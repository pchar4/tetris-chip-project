magic
tech scmos
timestamp 1712622712
<< metal1 >>
rect 14 3307 3490 3327
rect 38 3283 3466 3303
rect 14 3267 3490 3273
rect 530 3233 556 3236
rect 898 3233 916 3236
rect 1418 3233 1436 3236
rect 1610 3233 1660 3236
rect 1930 3233 1948 3236
rect 1962 3233 1996 3236
rect 2850 3233 2892 3236
rect 412 3223 437 3226
rect 530 3216 533 3233
rect 596 3223 637 3226
rect 924 3223 933 3226
rect 1050 3216 1053 3225
rect 1170 3223 1204 3226
rect 1444 3223 1453 3226
rect 1548 3223 1557 3226
rect 1604 3223 1653 3226
rect 1754 3223 1764 3226
rect 2004 3223 2013 3226
rect 74 3213 92 3216
rect 172 3213 197 3216
rect 284 3213 309 3216
rect 340 3213 373 3216
rect 380 3213 396 3216
rect 426 3213 444 3216
rect 476 3213 485 3216
rect 524 3213 533 3216
rect 594 3213 644 3216
rect 746 3213 764 3216
rect 788 3213 797 3216
rect 804 3213 813 3216
rect 818 3213 828 3216
rect 858 3213 892 3216
rect 962 3213 1004 3216
rect 1018 3213 1036 3216
rect 1050 3213 1061 3216
rect 1074 3213 1116 3216
rect 1156 3213 1197 3216
rect 1234 3213 1252 3216
rect 1298 3213 1324 3216
rect 1364 3213 1381 3216
rect 370 3205 373 3213
rect 746 3206 749 3213
rect 468 3203 493 3206
rect 642 3203 652 3206
rect 668 3203 685 3206
rect 708 3203 749 3206
rect 780 3203 789 3206
rect 794 3205 797 3213
rect 1450 3206 1453 3223
rect 2202 3216 2205 3225
rect 2338 3223 2356 3226
rect 2580 3223 2605 3226
rect 2900 3223 2917 3226
rect 3356 3223 3365 3226
rect 3394 3216 3397 3225
rect 1474 3213 1492 3216
rect 1506 3213 1532 3216
rect 1546 3213 1589 3216
rect 1690 3213 1700 3216
rect 1818 3206 1821 3214
rect 1826 3213 1852 3216
rect 1884 3213 1909 3216
rect 2084 3213 2093 3216
rect 2122 3213 2156 3216
rect 2202 3213 2220 3216
rect 2284 3213 2293 3216
rect 2332 3213 2349 3216
rect 866 3203 884 3206
rect 1052 3203 1060 3206
rect 1074 3203 1108 3206
rect 1140 3203 1148 3206
rect 1258 3203 1284 3206
rect 1290 3203 1316 3206
rect 1450 3203 1484 3206
rect 1514 3203 1524 3206
rect 1548 3203 1557 3206
rect 1578 3203 1588 3206
rect 1740 3203 1757 3206
rect 1794 3203 1812 3206
rect 1818 3203 1844 3206
rect 1916 3203 1925 3206
rect 2044 3203 2060 3206
rect 2116 3203 2148 3206
rect 2362 3203 2365 3214
rect 2386 3213 2404 3216
rect 2410 3213 2436 3216
rect 2466 3213 2476 3216
rect 2516 3213 2541 3216
rect 2410 3203 2428 3206
rect 2538 3205 2541 3213
rect 2578 3213 2613 3216
rect 2716 3213 2741 3216
rect 2820 3213 2829 3216
rect 2914 3213 2932 3216
rect 2986 3213 2997 3216
rect 3026 3213 3060 3216
rect 3236 3213 3261 3216
rect 3298 3213 3316 3216
rect 3330 3213 3340 3216
rect 3362 3213 3380 3216
rect 3394 3213 3412 3216
rect 2578 3205 2581 3213
rect 2594 3203 2612 3206
rect 2660 3203 2677 3206
rect 2778 3203 2804 3206
rect 2818 3203 2836 3206
rect 2906 3203 2924 3206
rect 2948 3203 2957 3206
rect 2994 3205 2997 3213
rect 3322 3203 3332 3206
rect 1706 3193 1732 3196
rect 1794 3193 1804 3196
rect 1890 3193 1908 3196
rect 2482 3193 2500 3196
rect 38 3167 3466 3173
rect 778 3143 796 3146
rect 1674 3136 1677 3145
rect 1804 3143 1813 3146
rect 202 3126 205 3134
rect 250 3126 253 3134
rect 418 3126 421 3134
rect 474 3133 485 3136
rect 508 3133 541 3136
rect 570 3133 580 3136
rect 626 3133 652 3136
rect 714 3133 748 3136
rect 764 3133 773 3136
rect 794 3133 804 3136
rect 810 3133 820 3136
rect 858 3133 876 3136
rect 946 3133 956 3136
rect 1010 3133 1020 3136
rect 1066 3133 1092 3136
rect 1122 3133 1132 3136
rect 1154 3133 1196 3136
rect 1226 3133 1236 3136
rect 1266 3133 1308 3136
rect 1338 3133 1348 3136
rect 1466 3133 1516 3136
rect 1586 3133 1644 3136
rect 1666 3133 1677 3136
rect 1754 3133 1788 3136
rect 116 3123 141 3126
rect 172 3123 205 3126
rect 242 3123 253 3126
rect 340 3123 365 3126
rect 396 3123 421 3126
rect 428 3123 444 3126
rect 474 3116 477 3133
rect 276 3113 293 3116
rect 460 3113 477 3116
rect 522 3123 540 3126
rect 610 3123 644 3126
rect 722 3123 740 3126
rect 772 3123 781 3126
rect 810 3125 813 3133
rect 858 3126 861 3133
rect 1834 3126 1837 3134
rect 1938 3133 1948 3136
rect 1972 3133 1981 3136
rect 2050 3133 2076 3136
rect 2082 3133 2108 3136
rect 2138 3126 2141 3134
rect 2170 3133 2212 3136
rect 2274 3133 2316 3136
rect 2378 3133 2413 3136
rect 844 3123 861 3126
rect 954 3123 964 3126
rect 978 3123 1004 3126
rect 1156 3123 1197 3126
rect 1218 3123 1228 3126
rect 1260 3123 1309 3126
rect 1372 3123 1389 3126
rect 1402 3123 1428 3126
rect 1482 3123 1524 3126
rect 1626 3123 1636 3126
rect 1668 3123 1677 3126
rect 1692 3123 1732 3126
rect 1770 3123 1780 3126
rect 1804 3123 1837 3126
rect 522 3093 525 3123
rect 604 3113 637 3116
rect 972 3113 989 3116
rect 1444 3113 1453 3116
rect 1468 3113 1477 3116
rect 1540 3113 1549 3116
rect 1874 3106 1877 3125
rect 1938 3123 1956 3126
rect 1970 3123 2004 3126
rect 2018 3123 2044 3126
rect 2084 3123 2101 3126
rect 2132 3123 2141 3126
rect 2298 3123 2308 3126
rect 2378 3125 2381 3133
rect 2386 3123 2428 3126
rect 2434 3123 2444 3126
rect 2458 3123 2461 3134
rect 2466 3133 2492 3136
rect 2522 3133 2540 3136
rect 2594 3133 2628 3136
rect 2772 3133 2781 3136
rect 2786 3133 2796 3136
rect 2876 3133 2884 3136
rect 2964 3133 2973 3136
rect 2994 3133 3020 3136
rect 3034 3133 3052 3136
rect 3066 3133 3100 3136
rect 3124 3133 3133 3136
rect 2778 3126 2781 3133
rect 3138 3126 3141 3134
rect 3252 3133 3260 3136
rect 3394 3133 3412 3136
rect 2474 3123 2500 3126
rect 2514 3123 2532 3126
rect 2572 3123 2613 3126
rect 2650 3123 2660 3126
rect 2698 3123 2748 3126
rect 2778 3123 2804 3126
rect 2810 3123 2852 3126
rect 2906 3123 2948 3126
rect 2962 3123 2988 3126
rect 3028 3123 3053 3126
rect 3060 3123 3101 3126
rect 3122 3123 3141 3126
rect 3148 3123 3181 3126
rect 3194 3123 3212 3126
rect 3268 3123 3285 3126
rect 3332 3123 3357 3126
rect 3420 3123 3437 3126
rect 1938 3116 1941 3123
rect 1916 3113 1941 3116
rect 1972 3113 1981 3116
rect 2020 3113 2029 3116
rect 2164 3113 2197 3116
rect 2460 3113 2485 3116
rect 2676 3113 2693 3116
rect 3068 3113 3093 3116
rect 1850 3103 1877 3106
rect 14 3067 3490 3073
rect 810 3033 844 3036
rect 236 3023 261 3026
rect 428 3023 445 3026
rect 604 3023 629 3026
rect 116 3013 141 3016
rect 172 3013 197 3016
rect 204 3013 220 3016
rect 300 3013 325 3016
rect 356 3013 389 3016
rect 396 3013 412 3016
rect 434 3013 452 3016
rect 194 3005 197 3013
rect 386 3005 389 3013
rect 482 3006 485 3014
rect 490 3013 516 3016
rect 562 3013 572 3016
rect 666 3013 676 3016
rect 698 3013 708 3016
rect 810 3006 813 3033
rect 818 3023 828 3026
rect 852 3023 861 3026
rect 916 3023 941 3026
rect 1260 3023 1277 3026
rect 1308 3023 1333 3026
rect 1428 3023 1445 3026
rect 2068 3023 2077 3026
rect 858 3013 884 3016
rect 922 3013 948 3016
rect 978 3006 981 3014
rect 1082 3013 1092 3016
rect 1098 3013 1124 3016
rect 1218 3013 1244 3016
rect 1266 3013 1292 3016
rect 1322 3013 1340 3016
rect 1386 3013 1412 3016
rect 1442 3013 1452 3016
rect 1548 3013 1565 3016
rect 1604 3013 1621 3016
rect 1626 3013 1644 3016
rect 1722 3013 1748 3016
rect 1802 3013 1812 3016
rect 1954 3013 1972 3016
rect 1986 3013 1996 3016
rect 2042 3013 2052 3016
rect 2066 3013 2108 3016
rect 450 3003 460 3006
rect 482 3003 517 3006
rect 546 3003 564 3006
rect 610 3003 636 3006
rect 754 3003 764 3006
rect 796 3003 813 3006
rect 866 3003 876 3006
rect 930 3003 956 3006
rect 978 3003 989 3006
rect 1002 3003 1012 3006
rect 1260 3003 1269 3006
rect 1274 3003 1284 3006
rect 1364 3003 1381 3006
rect 1394 3003 1404 3006
rect 1434 3003 1460 3006
rect 1506 3003 1524 3006
rect 1546 3003 1580 3006
rect 1668 3003 1685 3006
rect 1730 3003 1756 3006
rect 1786 3003 1820 3006
rect 1850 3003 1876 3006
rect 1898 3003 1924 3006
rect 2034 3003 2044 3006
rect 2074 3003 2100 3006
rect 2114 3003 2117 3014
rect 2178 3013 2188 3016
rect 2228 3013 2237 3016
rect 2274 3013 2308 3016
rect 2354 3013 2404 3016
rect 2410 3013 2436 3016
rect 2274 3006 2277 3013
rect 2514 3006 2517 3036
rect 2858 3016 2861 3026
rect 2586 3013 2636 3016
rect 2660 3013 2669 3016
rect 2706 3013 2756 3016
rect 2786 3013 2820 3016
rect 2826 3013 2861 3016
rect 2866 3013 2884 3016
rect 2940 3013 2949 3016
rect 3028 3013 3045 3016
rect 3218 3013 3252 3016
rect 2170 3003 2180 3006
rect 2194 3003 2204 3006
rect 2266 3003 2277 3006
rect 2362 3003 2396 3006
rect 2418 3003 2428 3006
rect 2458 3003 2476 3006
rect 2482 3003 2532 3006
rect 2554 3003 2572 3006
rect 2578 3003 2644 3006
rect 2658 3003 2668 3006
rect 2714 3003 2748 3006
rect 2826 3003 2836 3006
rect 2850 3003 2876 3006
rect 2900 3003 2925 3006
rect 2970 3003 3020 3006
rect 3034 3003 3044 3006
rect 3068 3003 3101 3006
rect 3202 3003 3244 3006
rect 778 2993 788 2996
rect 2242 2993 2252 2996
rect 2826 2983 2829 3003
rect 38 2967 3466 2973
rect 74 2943 92 2946
rect 100 2933 117 2936
rect 132 2933 149 2936
rect 156 2933 197 2936
rect 330 2926 333 2935
rect 346 2926 349 2945
rect 714 2936 717 2946
rect 546 2926 549 2935
rect 626 2933 636 2936
rect 658 2933 677 2936
rect 714 2933 741 2936
rect 804 2933 844 2936
rect 860 2933 869 2936
rect 890 2933 900 2936
rect 924 2933 964 2936
rect 1186 2933 1212 2936
rect 1268 2933 1301 2936
rect 1570 2933 1588 2936
rect 1722 2933 1748 2936
rect 1820 2933 1837 2936
rect 1858 2933 1884 2936
rect 108 2923 125 2926
rect 236 2923 261 2926
rect 292 2923 333 2926
rect 340 2923 349 2926
rect 370 2923 380 2926
rect 460 2923 485 2926
rect 516 2923 549 2926
rect 556 2923 572 2926
rect 618 2923 628 2926
rect 658 2925 661 2933
rect 666 2923 676 2926
rect 738 2925 741 2933
rect 1834 2926 1837 2933
rect 2010 2926 2013 2935
rect 2202 2926 2205 2935
rect 2340 2933 2349 2936
rect 2394 2933 2404 2936
rect 2460 2933 2509 2936
rect 2514 2926 2517 2935
rect 994 2923 1004 2926
rect 1010 2923 1028 2926
rect 1092 2923 1117 2926
rect 1154 2923 1164 2926
rect 1202 2923 1220 2926
rect 1282 2923 1308 2926
rect 1340 2923 1349 2926
rect 1388 2923 1413 2926
rect 1508 2923 1533 2926
rect 1570 2923 1596 2926
rect 1666 2923 1692 2926
rect 1724 2923 1733 2926
rect 1778 2923 1796 2926
rect 1834 2923 1852 2926
rect 2010 2923 2021 2926
rect 2154 2923 2188 2926
rect 2202 2923 2213 2926
rect 2250 2923 2276 2926
rect 2338 2923 2380 2926
rect 2386 2923 2412 2926
rect 2490 2923 2517 2926
rect 2706 2923 2724 2926
rect 3068 2923 3077 2926
rect 3268 2923 3293 2926
rect 3324 2923 3333 2926
rect 396 2913 421 2916
rect 588 2913 621 2916
rect 1908 2913 1917 2916
rect 2826 2913 2844 2916
rect 3076 2913 3085 2916
rect 2834 2903 2860 2906
rect 3090 2903 3140 2906
rect 14 2867 3490 2873
rect 3178 2833 3236 2836
rect 564 2823 581 2826
rect 1172 2823 1189 2826
rect 1660 2823 1677 2826
rect 2116 2823 2125 2826
rect 3172 2823 3220 2826
rect 340 2813 365 2816
rect 634 2813 652 2816
rect 706 2813 724 2816
rect 754 2813 772 2816
rect 1052 2813 1077 2816
rect 1108 2813 1133 2816
rect 1140 2813 1156 2816
rect 1338 2813 1356 2816
rect 1508 2813 1517 2816
rect 1556 2813 1581 2816
rect 1716 2813 1741 2816
rect 1778 2813 1796 2816
rect 1868 2813 1893 2816
rect 2012 2813 2037 2816
rect 2068 2813 2077 2816
rect 2084 2813 2100 2816
rect 2180 2813 2205 2816
rect 2276 2813 2301 2816
rect 2332 2813 2341 2816
rect 2548 2813 2557 2816
rect 2628 2813 2653 2816
rect 2684 2813 2693 2816
rect 2956 2813 2965 2816
rect 3146 2813 3164 2816
rect 3284 2813 3301 2816
rect 3428 2813 3437 2816
rect 410 2803 436 2806
rect 450 2803 460 2806
rect 466 2803 484 2806
rect 522 2803 540 2806
rect 564 2803 573 2806
rect 612 2803 645 2806
rect 676 2803 701 2806
rect 746 2803 764 2806
rect 836 2803 853 2806
rect 922 2803 940 2806
rect 980 2803 989 2806
rect 1130 2805 1133 2813
rect 1298 2803 1316 2806
rect 1618 2803 1636 2806
rect 2074 2805 2077 2813
rect 2338 2805 2341 2813
rect 2514 2803 2540 2806
rect 2564 2803 2589 2806
rect 2962 2805 2965 2813
rect 3250 2803 3276 2806
rect 402 2793 428 2796
rect 794 2793 828 2796
rect 2546 2793 2556 2796
rect 3298 2795 3301 2813
rect 3308 2803 3333 2806
rect 38 2767 3466 2773
rect 586 2726 589 2735
rect 602 2726 605 2745
rect 674 2743 692 2746
rect 674 2733 700 2736
rect 706 2733 716 2736
rect 882 2726 885 2735
rect 898 2726 901 2745
rect 1106 2743 1116 2746
rect 1642 2745 1652 2746
rect 1090 2726 1093 2735
rect 1106 2726 1109 2743
rect 1124 2733 1141 2736
rect 1242 2726 1245 2745
rect 1642 2743 1653 2745
rect 1332 2733 1349 2736
rect 1356 2733 1413 2736
rect 1572 2733 1605 2736
rect 1650 2726 1653 2743
rect 1660 2733 1669 2736
rect 1714 2726 1717 2756
rect 1818 2743 1828 2746
rect 1754 2733 1764 2736
rect 1788 2733 1805 2736
rect 1994 2733 2028 2736
rect 2066 2733 2076 2736
rect 2108 2733 2125 2736
rect 2172 2733 2189 2736
rect 2306 2733 2324 2736
rect 2122 2726 2125 2733
rect 2706 2726 2709 2745
rect 2722 2743 2756 2746
rect 2770 2743 2804 2746
rect 2730 2733 2764 2736
rect 2802 2733 2812 2736
rect 3188 2733 3197 2736
rect 3218 2733 3252 2736
rect 3282 2733 3292 2736
rect 148 2723 157 2726
rect 268 2723 293 2726
rect 324 2723 333 2726
rect 388 2723 413 2726
rect 500 2723 525 2726
rect 556 2723 589 2726
rect 596 2723 605 2726
rect 642 2723 660 2726
rect 724 2723 741 2726
rect 804 2723 821 2726
rect 860 2723 885 2726
rect 892 2723 901 2726
rect 1044 2723 1093 2726
rect 1100 2723 1109 2726
rect 1202 2723 1245 2726
rect 1260 2723 1325 2726
rect 1508 2723 1533 2726
rect 1620 2723 1653 2726
rect 1684 2723 1717 2726
rect 1732 2723 1765 2726
rect 1772 2723 1781 2726
rect 1796 2723 1821 2726
rect 1932 2723 1957 2726
rect 1988 2723 2005 2726
rect 2122 2723 2140 2726
rect 2244 2723 2269 2726
rect 2300 2723 2309 2726
rect 2380 2723 2389 2726
rect 2492 2723 2517 2726
rect 2700 2723 2709 2726
rect 2772 2723 2797 2726
rect 2826 2723 2836 2726
rect 2916 2723 2933 2726
rect 3028 2723 3053 2726
rect 3138 2706 3141 2725
rect 3162 2723 3172 2726
rect 3234 2723 3260 2726
rect 3276 2723 3293 2726
rect 3364 2723 3389 2726
rect 3122 2703 3141 2706
rect 14 2667 3490 2673
rect 3156 2623 3189 2626
rect 3434 2616 3437 2656
rect 82 2613 92 2616
rect 124 2613 149 2616
rect 188 2613 205 2616
rect 268 2613 285 2616
rect 290 2613 300 2616
rect 404 2613 429 2616
rect 460 2613 493 2616
rect 498 2613 508 2616
rect 524 2613 533 2616
rect 604 2613 613 2616
rect 820 2613 845 2616
rect 876 2613 885 2616
rect 980 2613 989 2616
rect 1028 2613 1053 2616
rect 1244 2613 1253 2616
rect 1300 2613 1309 2616
rect 1412 2613 1437 2616
rect 1482 2613 1500 2616
rect 1828 2613 1837 2616
rect 2060 2613 2069 2616
rect 2180 2613 2189 2616
rect 2236 2613 2269 2616
rect 2420 2613 2445 2616
rect 2556 2613 2581 2616
rect 2676 2613 2701 2616
rect 2732 2613 2741 2616
rect 2788 2613 2805 2616
rect 2916 2613 2925 2616
rect 2980 2613 2989 2616
rect 3084 2613 3093 2616
rect 3170 2613 3220 2616
rect 3330 2606 3333 2614
rect 3420 2613 3437 2616
rect 130 2603 164 2606
rect 186 2603 244 2606
rect 324 2603 357 2606
rect 466 2603 500 2606
rect 1474 2603 1508 2606
rect 2340 2603 2357 2606
rect 2468 2603 2476 2606
rect 2850 2603 2892 2606
rect 3050 2603 3076 2606
rect 3162 2603 3212 2606
rect 3292 2603 3333 2606
rect 3370 2603 3412 2606
rect 3250 2593 3284 2596
rect 3370 2593 3373 2603
rect 3378 2593 3404 2596
rect 38 2567 3466 2573
rect 306 2533 340 2536
rect 370 2533 420 2536
rect 538 2533 572 2536
rect 746 2533 812 2536
rect 828 2533 869 2536
rect 914 2533 964 2536
rect 1122 2533 1156 2536
rect 1178 2533 1197 2536
rect 1228 2533 1253 2536
rect 1562 2533 1596 2536
rect 1618 2533 1661 2536
rect 1740 2533 1757 2536
rect 1994 2533 2044 2536
rect 2060 2533 2093 2536
rect 2170 2533 2228 2536
rect 2290 2533 2324 2536
rect 2474 2533 2516 2536
rect 2538 2533 2597 2536
rect 2626 2533 2676 2536
rect 2698 2533 2741 2536
rect 2778 2533 2829 2536
rect 124 2523 149 2526
rect 236 2523 245 2526
rect 292 2523 332 2526
rect 562 2523 580 2526
rect 610 2523 620 2526
rect 748 2523 757 2526
rect 762 2523 804 2526
rect 836 2523 861 2526
rect 866 2523 876 2526
rect 988 2523 1021 2526
rect 1060 2523 1085 2526
rect 1116 2523 1141 2526
rect 1178 2525 1181 2533
rect 1186 2523 1204 2526
rect 1236 2523 1245 2526
rect 1292 2523 1309 2526
rect 1348 2523 1357 2526
rect 1396 2523 1421 2526
rect 1452 2523 1461 2526
rect 1556 2523 1588 2526
rect 1618 2525 1621 2533
rect 1626 2523 1660 2526
rect 1692 2523 1717 2526
rect 1746 2523 1756 2526
rect 1788 2523 1829 2526
rect 1868 2523 1885 2526
rect 1996 2523 2005 2526
rect 2068 2523 2109 2526
rect 2172 2523 2205 2526
rect 2252 2523 2261 2526
rect 2444 2523 2452 2526
rect 2538 2525 2541 2533
rect 2628 2523 2637 2526
rect 2698 2525 2701 2533
rect 2738 2523 2748 2526
rect 2778 2525 2781 2533
rect 3170 2526 3173 2535
rect 2860 2523 2877 2526
rect 2988 2523 3021 2526
rect 3084 2523 3093 2526
rect 3098 2523 3148 2526
rect 3162 2523 3173 2526
rect 3268 2523 3293 2526
rect 3324 2523 3333 2526
rect 3428 2523 3501 2526
rect 3018 2506 3021 2523
rect 3028 2513 3037 2516
rect 3196 2513 3213 2516
rect 3018 2503 3044 2506
rect 14 2467 3490 2473
rect 3498 2456 3501 2523
rect 3426 2453 3501 2456
rect 3322 2433 3341 2436
rect 3394 2433 3412 2436
rect 1316 2423 1333 2426
rect 1364 2423 1405 2426
rect 1436 2423 1453 2426
rect 3322 2423 3332 2426
rect 172 2413 181 2416
rect 228 2413 245 2416
rect 284 2413 293 2416
rect 340 2413 365 2416
rect 396 2413 413 2416
rect 452 2413 477 2416
rect 564 2413 573 2416
rect 620 2413 629 2416
rect 668 2413 685 2416
rect 892 2413 917 2416
rect 1188 2413 1213 2416
rect 1266 2413 1300 2416
rect 1314 2413 1348 2416
rect 1410 2413 1420 2416
rect 1556 2413 1581 2416
rect 1612 2413 1621 2416
rect 1668 2413 1693 2416
rect 1724 2413 1733 2416
rect 1804 2413 1829 2416
rect 1908 2413 1933 2416
rect 2004 2413 2029 2416
rect 2108 2413 2133 2416
rect 2204 2413 2229 2416
rect 2300 2413 2325 2416
rect 2500 2413 2509 2416
rect 2596 2413 2621 2416
rect 2700 2413 2725 2416
rect 2796 2413 2821 2416
rect 2892 2413 2917 2416
rect 2996 2413 3013 2416
rect 3148 2413 3157 2416
rect 3252 2413 3285 2416
rect 1066 2403 1100 2406
rect 1370 2403 1412 2406
rect 1442 2403 1460 2406
rect 1484 2403 1501 2406
rect 3282 2405 3285 2413
rect 3322 2406 3325 2423
rect 3338 2415 3341 2433
rect 3362 2423 3396 2426
rect 3420 2423 3429 2426
rect 3308 2403 3325 2406
rect 38 2367 3466 2373
rect 258 2333 268 2336
rect 306 2333 316 2336
rect 354 2333 396 2336
rect 426 2333 460 2336
rect 506 2333 524 2336
rect 548 2333 573 2336
rect 626 2333 660 2336
rect 690 2333 724 2336
rect 748 2333 781 2336
rect 812 2333 837 2336
rect 882 2333 900 2336
rect 930 2333 964 2336
rect 1034 2333 1068 2336
rect 1114 2333 1140 2336
rect 1170 2333 1212 2336
rect 1234 2326 1237 2335
rect 1284 2333 1293 2336
rect 1306 2333 1332 2336
rect 1356 2333 1365 2336
rect 1418 2333 1452 2336
rect 1474 2326 1477 2335
rect 1524 2333 1533 2336
rect 1770 2333 1788 2336
rect 1826 2333 1852 2336
rect 1882 2333 1916 2336
rect 1962 2333 1980 2336
rect 2004 2333 2037 2336
rect 2082 2333 2108 2336
rect 2204 2333 2229 2336
rect 2266 2333 2300 2336
rect 2330 2333 2364 2336
rect 2388 2333 2397 2336
rect 2402 2333 2428 2336
rect 2452 2333 2477 2336
rect 2482 2326 2485 2335
rect 2514 2333 2548 2336
rect 2572 2333 2597 2336
rect 2682 2333 2700 2336
rect 2794 2326 2797 2356
rect 3138 2343 3148 2346
rect 3322 2336 3325 2346
rect 2802 2333 2828 2336
rect 2852 2333 2861 2336
rect 2866 2333 2900 2336
rect 2954 2333 2988 2336
rect 3034 2333 3052 2336
rect 3156 2333 3172 2336
rect 3218 2333 3244 2336
rect 3258 2333 3276 2336
rect 3300 2333 3308 2336
rect 3322 2333 3364 2336
rect 3388 2333 3396 2336
rect 164 2323 189 2326
rect 220 2323 237 2326
rect 386 2323 404 2326
rect 618 2323 668 2326
rect 746 2323 796 2326
rect 874 2323 908 2326
rect 962 2323 972 2326
rect 1076 2323 1085 2326
rect 1162 2323 1220 2326
rect 1234 2323 1268 2326
rect 1354 2323 1396 2326
rect 1410 2323 1460 2326
rect 1474 2323 1508 2326
rect 1522 2323 1580 2326
rect 1850 2323 1860 2326
rect 1978 2323 1988 2326
rect 2090 2323 2116 2326
rect 2178 2323 2188 2326
rect 2258 2323 2308 2326
rect 2362 2323 2372 2326
rect 2450 2323 2485 2326
rect 2642 2323 2660 2326
rect 2794 2323 2836 2326
rect 2930 2323 2948 2326
rect 3082 2323 3092 2326
rect 3180 2323 3189 2326
rect 420 2313 437 2316
rect 484 2313 517 2316
rect 684 2313 717 2316
rect 748 2313 781 2316
rect 924 2313 957 2316
rect 1108 2313 1117 2316
rect 1164 2313 1197 2316
rect 1356 2313 1381 2316
rect 1412 2313 1445 2316
rect 1476 2313 1493 2316
rect 1596 2313 1613 2316
rect 1684 2313 1701 2316
rect 1876 2313 1901 2316
rect 2068 2313 2077 2316
rect 2260 2313 2269 2316
rect 2724 2313 2757 2316
rect 2852 2313 2877 2316
rect 3012 2313 3045 2316
rect 3188 2313 3205 2316
rect 3258 2315 3261 2333
rect 3298 2323 3333 2326
rect 3362 2323 3372 2326
rect 3394 2323 3429 2326
rect 3330 2313 3333 2323
rect 3426 2313 3429 2323
rect 1114 2303 1117 2313
rect 1610 2303 1613 2313
rect 14 2267 3490 2273
rect 116 2223 133 2226
rect 172 2223 181 2226
rect 244 2223 269 2226
rect 308 2223 325 2226
rect 364 2223 381 2226
rect 604 2223 629 2226
rect 1290 2223 1309 2226
rect 1820 2223 1837 2226
rect 1868 2223 1901 2226
rect 2300 2223 2309 2226
rect 2428 2223 2453 2226
rect 3004 2223 3021 2226
rect 3052 2223 3061 2226
rect 82 2213 100 2216
rect 122 2213 156 2216
rect 306 2213 349 2216
rect 356 2213 381 2216
rect 394 2213 404 2216
rect 426 2213 468 2216
rect 490 2213 524 2216
rect 548 2213 581 2216
rect 586 2213 596 2216
rect 602 2213 652 2216
rect 682 2213 724 2216
rect 796 2213 813 2216
rect 818 2213 852 2216
rect 866 2213 876 2216
rect 898 2213 932 2216
rect 964 2213 973 2216
rect 1020 2213 1045 2216
rect 1108 2213 1141 2216
rect 1170 2213 1204 2216
rect 82 2203 92 2206
rect 138 2203 148 2206
rect 186 2203 220 2206
rect 258 2203 284 2206
rect 308 2203 341 2206
rect 346 2205 349 2213
rect 378 2206 381 2213
rect 1290 2206 1293 2223
rect 1298 2213 1324 2216
rect 1402 2213 1412 2216
rect 1450 2213 1468 2216
rect 1570 2213 1596 2216
rect 1634 2213 1644 2216
rect 1708 2213 1717 2216
rect 1756 2213 1765 2216
rect 1770 2213 1812 2216
rect 1818 2213 1852 2216
rect 1866 2213 1916 2216
rect 2108 2213 2125 2216
rect 2194 2213 2228 2216
rect 2260 2213 2269 2216
rect 2274 2213 2292 2216
rect 2314 2213 2340 2216
rect 2394 2213 2420 2216
rect 2442 2213 2468 2216
rect 2474 2213 2492 2216
rect 2562 2213 2580 2216
rect 2634 2213 2652 2216
rect 2666 2213 2684 2216
rect 2690 2213 2724 2216
rect 2754 2213 2772 2216
rect 3002 2213 3036 2216
rect 3074 2213 3108 2216
rect 3170 2213 3196 2216
rect 3276 2213 3285 2216
rect 3412 2213 3429 2216
rect 2266 2206 2269 2213
rect 2394 2206 2397 2213
rect 2754 2206 2757 2213
rect 378 2203 396 2206
rect 420 2203 437 2206
rect 442 2203 460 2206
rect 530 2203 540 2206
rect 722 2203 732 2206
rect 802 2203 844 2206
rect 892 2203 925 2206
rect 1026 2203 1044 2206
rect 1068 2203 1085 2206
rect 1114 2203 1140 2206
rect 1170 2203 1212 2206
rect 1276 2203 1293 2206
rect 1298 2203 1316 2206
rect 1364 2203 1381 2206
rect 1450 2203 1460 2206
rect 1474 2203 1524 2206
rect 1548 2203 1581 2206
rect 1586 2203 1604 2206
rect 1626 2203 1636 2206
rect 1650 2203 1700 2206
rect 1762 2203 1804 2206
rect 1868 2203 1909 2206
rect 2010 2203 2044 2206
rect 2252 2203 2261 2206
rect 2266 2203 2277 2206
rect 2314 2203 2348 2206
rect 2364 2203 2397 2206
rect 2740 2203 2757 2206
rect 2890 2203 2908 2206
rect 2946 2203 2980 2206
rect 3052 2203 3069 2206
rect 3082 2203 3100 2206
rect 3298 2203 3348 2206
rect 3378 2203 3404 2206
rect 1298 2196 1301 2203
rect 1242 2193 1268 2196
rect 1282 2193 1301 2196
rect 1346 2193 1356 2196
rect 1506 2193 1516 2196
rect 3210 2193 3220 2196
rect 38 2167 3466 2173
rect 3010 2153 3029 2156
rect 882 2143 924 2146
rect 938 2143 948 2146
rect 122 2133 172 2136
rect 226 2133 276 2136
rect 292 2133 317 2136
rect 404 2133 429 2136
rect 602 2133 613 2136
rect 642 2133 660 2136
rect 682 2133 716 2136
rect 314 2126 317 2133
rect 124 2123 173 2126
rect 180 2123 189 2126
rect 234 2123 268 2126
rect 314 2123 332 2126
rect 354 2123 380 2126
rect 434 2123 452 2126
rect 610 2116 613 2133
rect 626 2123 652 2126
rect 754 2123 812 2126
rect 844 2123 853 2126
rect 938 2125 941 2143
rect 970 2126 973 2146
rect 1298 2143 1333 2146
rect 1330 2136 1333 2143
rect 3346 2136 3349 2146
rect 1018 2133 1028 2136
rect 1042 2133 1060 2136
rect 1076 2133 1109 2136
rect 1148 2133 1157 2136
rect 1162 2133 1188 2136
rect 1204 2133 1229 2136
rect 1234 2133 1252 2136
rect 1306 2133 1325 2136
rect 1330 2133 1340 2136
rect 1364 2133 1373 2136
rect 1380 2133 1389 2136
rect 1394 2133 1413 2136
rect 1452 2133 1477 2136
rect 1524 2133 1556 2136
rect 1618 2133 1636 2136
rect 1106 2126 1109 2133
rect 1410 2126 1413 2133
rect 1666 2126 1669 2135
rect 1692 2133 1709 2136
rect 1746 2133 1756 2136
rect 970 2123 988 2126
rect 1018 2123 1036 2126
rect 1106 2123 1124 2126
rect 1170 2123 1180 2126
rect 1212 2123 1221 2126
rect 1284 2123 1341 2126
rect 1388 2123 1405 2126
rect 1410 2123 1428 2126
rect 1466 2123 1500 2126
rect 1530 2123 1564 2126
rect 1652 2123 1669 2126
rect 1676 2123 1685 2126
rect 1778 2125 1781 2136
rect 1802 2133 1868 2136
rect 1898 2133 1908 2136
rect 1938 2126 1941 2136
rect 1946 2133 1964 2136
rect 2036 2133 2077 2136
rect 2108 2133 2117 2136
rect 2204 2133 2237 2136
rect 2242 2133 2252 2136
rect 2269 2133 2324 2136
rect 2394 2133 2403 2136
rect 2434 2133 2460 2136
rect 2476 2133 2517 2136
rect 2740 2133 2757 2136
rect 3010 2133 3036 2136
rect 3066 2133 3084 2136
rect 3116 2133 3141 2136
rect 3226 2133 3252 2136
rect 3266 2133 3292 2136
rect 3306 2133 3316 2136
rect 3346 2133 3356 2136
rect 1796 2123 1821 2126
rect 1892 2123 1909 2126
rect 1938 2123 1972 2126
rect 2140 2123 2165 2126
rect 2226 2123 2244 2126
rect 2306 2123 2316 2126
rect 2362 2123 2372 2126
rect 2378 2123 2411 2126
rect 2506 2123 2532 2126
rect 2652 2123 2669 2126
rect 2770 2123 2780 2126
rect 2826 2123 2836 2126
rect 2852 2123 2877 2126
rect 2914 2123 2940 2126
rect 3082 2123 3092 2126
rect 3220 2123 3245 2126
rect 3250 2123 3260 2126
rect 3338 2123 3364 2126
rect 3402 2123 3412 2126
rect 188 2113 197 2116
rect 340 2113 373 2116
rect 610 2113 645 2116
rect 732 2113 741 2116
rect 506 2103 532 2106
rect 850 2103 853 2123
rect 1218 2103 1221 2123
rect 1292 2113 1333 2116
rect 1402 2113 1405 2123
rect 1924 2113 1957 2116
rect 2428 2113 2445 2116
rect 2860 2113 2869 2116
rect 14 2067 3490 2073
rect 378 2033 420 2036
rect 188 2023 205 2026
rect 372 2023 381 2026
rect 404 2023 413 2026
rect 474 2016 477 2046
rect 506 2033 516 2036
rect 82 2013 109 2016
rect 140 2013 149 2016
rect 180 2013 189 2016
rect 330 2013 364 2016
rect 442 2013 477 2016
rect 482 2023 500 2026
rect 564 2023 573 2026
rect 714 2023 733 2026
rect 66 2003 92 2006
rect 186 2003 189 2013
rect 482 2006 485 2023
rect 714 2016 717 2023
rect 818 2016 821 2036
rect 962 2033 980 2036
rect 954 2023 964 2026
rect 1122 2016 1125 2046
rect 1850 2043 1869 2046
rect 1850 2016 1853 2043
rect 1970 2033 2028 2036
rect 1964 2023 1989 2026
rect 2036 2023 2045 2026
rect 2140 2023 2149 2026
rect 2188 2023 2197 2026
rect 546 2013 556 2016
rect 586 2013 603 2016
rect 636 2013 645 2016
rect 700 2013 717 2016
rect 722 2013 748 2016
rect 796 2013 812 2016
rect 818 2013 860 2016
rect 1012 2013 1021 2016
rect 1066 2013 1076 2016
rect 1090 2013 1100 2016
rect 1122 2013 1164 2016
rect 1178 2013 1197 2016
rect 1306 2013 1324 2016
rect 1346 2013 1356 2016
rect 1410 2013 1436 2016
rect 1474 2013 1484 2016
rect 1666 2013 1685 2016
rect 1788 2013 1805 2016
rect 1844 2013 1853 2016
rect 1858 2013 1884 2016
rect 2042 2013 2068 2016
rect 2170 2013 2180 2016
rect 2300 2013 2309 2016
rect 722 2006 725 2013
rect 282 2003 300 2006
rect 316 2003 341 2006
rect 466 2003 485 2006
rect 538 2003 548 2006
rect 570 2003 596 2006
rect 650 2003 676 2006
rect 692 2003 725 2006
rect 730 2003 740 2006
rect 770 2003 788 2006
rect 850 2003 868 2006
rect 884 2003 893 2006
rect 898 2003 908 2006
rect 1034 2003 1068 2006
rect 1082 2003 1092 2006
rect 1122 2003 1156 2006
rect 1178 2005 1181 2013
rect 1186 2003 1212 2006
rect 1242 2003 1252 2006
rect 1306 2003 1316 2006
rect 1340 2003 1348 2006
rect 1396 2003 1437 2006
rect 1466 2003 1476 2006
rect 1490 2003 1548 2006
rect 1588 2003 1613 2006
rect 1618 2003 1644 2006
rect 1666 2005 1669 2013
rect 1724 2003 1733 2006
rect 1836 2003 1869 2006
rect 1906 2003 1916 2006
rect 2042 2003 2060 2006
rect 2074 2003 2084 2006
rect 2194 2003 2244 2006
rect 2314 2003 2340 2006
rect 2354 2003 2357 2025
rect 2642 2023 2653 2026
rect 2642 2016 2645 2023
rect 2412 2013 2429 2016
rect 2442 2013 2476 2016
rect 2490 2013 2500 2016
rect 2588 2013 2597 2016
rect 2636 2013 2645 2016
rect 2650 2013 2676 2016
rect 2738 2013 2772 2016
rect 2962 2013 2972 2016
rect 3018 2013 3036 2016
rect 3050 2013 3100 2016
rect 3130 2013 3180 2016
rect 3252 2013 3261 2016
rect 3282 2013 3340 2016
rect 3356 2013 3365 2016
rect 2434 2003 2468 2006
rect 2580 2003 2597 2006
rect 2740 2003 2780 2006
rect 2796 2003 2837 2006
rect 2916 2003 2925 2006
rect 2954 2003 2964 2006
rect 3018 2003 3028 2006
rect 3052 2003 3061 2006
rect 3066 2003 3092 2006
rect 3130 2003 3172 2006
rect 3196 2003 3205 2006
rect 3210 2003 3244 2006
rect 3250 2003 3260 2006
rect 3290 2003 3332 2006
rect 730 1996 733 2003
rect 714 1993 733 1996
rect 938 1993 957 1996
rect 1268 1993 1285 1996
rect 1362 1993 1388 1996
rect 2194 1983 2197 2003
rect 2594 1983 2597 2003
rect 3226 1993 3236 1996
rect 38 1967 3466 1973
rect 162 1936 165 1945
rect 594 1943 612 1946
rect 114 1926 117 1934
rect 140 1933 165 1936
rect 172 1933 197 1936
rect 202 1933 220 1936
rect 236 1933 269 1936
rect 362 1933 380 1936
rect 426 1933 444 1936
rect 474 1933 508 1936
rect 538 1933 556 1936
rect 650 1933 668 1936
rect 690 1933 701 1936
rect 714 1933 724 1936
rect 748 1933 757 1936
rect 92 1923 117 1926
rect 154 1923 165 1926
rect 180 1923 189 1926
rect 194 1923 212 1926
rect 244 1923 253 1926
rect 154 1916 157 1923
rect 194 1916 197 1923
rect 140 1913 157 1916
rect 186 1913 197 1916
rect 250 1903 253 1923
rect 362 1916 365 1933
rect 698 1926 701 1933
rect 762 1926 765 1956
rect 884 1943 893 1946
rect 1482 1943 1500 1946
rect 1482 1936 1485 1943
rect 778 1933 788 1936
rect 842 1933 868 1936
rect 924 1933 933 1936
rect 994 1933 1011 1936
rect 1042 1926 1045 1936
rect 1066 1933 1092 1936
rect 1108 1933 1117 1936
rect 1122 1933 1140 1936
rect 1154 1933 1204 1936
rect 1210 1933 1236 1936
rect 1252 1933 1261 1936
rect 1332 1933 1341 1936
rect 1346 1933 1356 1936
rect 1378 1933 1412 1936
rect 1452 1933 1485 1936
rect 1490 1933 1508 1936
rect 1490 1926 1493 1933
rect 404 1923 413 1926
rect 474 1923 500 1926
rect 554 1923 564 1926
rect 580 1923 605 1926
rect 628 1923 645 1926
rect 698 1923 732 1926
rect 762 1923 780 1926
rect 826 1923 860 1926
rect 884 1923 901 1926
rect 1042 1923 1084 1926
rect 1116 1923 1141 1926
rect 1148 1923 1189 1926
rect 1212 1923 1221 1926
rect 1266 1923 1308 1926
rect 1370 1923 1420 1926
rect 1466 1923 1493 1926
rect 1514 1925 1517 1946
rect 1858 1936 1861 1956
rect 1882 1953 1901 1956
rect 3002 1943 3021 1946
rect 3114 1943 3148 1946
rect 3018 1936 3021 1943
rect 3250 1936 3253 1946
rect 3306 1936 3309 1946
rect 1554 1933 1588 1936
rect 1762 1933 1804 1936
rect 1850 1933 1861 1936
rect 1986 1933 2028 1936
rect 2052 1933 2061 1936
rect 2066 1933 2076 1936
rect 2090 1933 2101 1936
rect 2162 1933 2180 1936
rect 2196 1933 2237 1936
rect 2482 1933 2492 1936
rect 2604 1933 2613 1936
rect 2674 1933 2684 1936
rect 2714 1933 2748 1936
rect 2762 1933 2772 1936
rect 2996 1933 3013 1936
rect 3018 1933 3028 1936
rect 3052 1933 3061 1936
rect 3066 1933 3084 1936
rect 3108 1933 3133 1936
rect 3138 1933 3156 1936
rect 3162 1933 3188 1936
rect 3226 1933 3268 1936
rect 3292 1933 3309 1936
rect 3428 1933 3437 1936
rect 1850 1926 1853 1933
rect 1612 1923 1621 1926
rect 1658 1923 1692 1926
rect 1724 1923 1733 1926
rect 1786 1923 1796 1926
rect 1828 1923 1837 1926
rect 1844 1923 1853 1926
rect 1874 1923 1916 1926
rect 1954 1923 1972 1926
rect 2026 1923 2036 1926
rect 2090 1925 2093 1933
rect 2162 1926 2165 1933
rect 2762 1926 2765 1933
rect 2098 1923 2165 1926
rect 2274 1923 2291 1926
rect 2306 1923 2332 1926
rect 2698 1923 2765 1926
rect 2826 1923 2844 1926
rect 2850 1923 2900 1926
rect 2940 1923 2965 1926
rect 3082 1923 3092 1926
rect 3164 1923 3181 1926
rect 3186 1923 3196 1926
rect 3276 1923 3285 1926
rect 3348 1923 3357 1926
rect 1618 1916 1621 1923
rect 306 1913 324 1916
rect 348 1913 365 1916
rect 938 1913 964 1916
rect 1156 1913 1173 1916
rect 1372 1913 1405 1916
rect 1548 1913 1573 1916
rect 1618 1913 1628 1916
rect 1748 1913 1789 1916
rect 266 1903 292 1906
rect 2098 1883 2101 1923
rect 2269 1913 2277 1916
rect 2388 1913 2397 1916
rect 2434 1913 2453 1916
rect 2548 1913 2557 1916
rect 3052 1913 3061 1916
rect 3108 1913 3117 1916
rect 3220 1913 3237 1916
rect 2218 1903 2260 1906
rect 2298 1883 2301 1906
rect 2378 1903 2403 1906
rect 2530 1903 2564 1906
rect 14 1867 3490 1873
rect 666 1853 693 1856
rect 2682 1853 2701 1856
rect 626 1833 652 1836
rect 698 1833 714 1836
rect 1098 1833 1125 1836
rect 164 1823 181 1826
rect 268 1823 293 1826
rect 348 1823 357 1826
rect 146 1813 156 1816
rect 82 1803 108 1806
rect 124 1803 133 1806
rect 178 1786 181 1823
rect 602 1816 605 1826
rect 626 1823 636 1826
rect 660 1823 669 1826
rect 690 1823 700 1826
rect 884 1823 909 1826
rect 228 1813 245 1816
rect 266 1813 340 1816
rect 364 1813 397 1816
rect 444 1813 477 1816
rect 524 1813 557 1816
rect 596 1813 605 1816
rect 186 1803 220 1806
rect 242 1805 245 1813
rect 394 1806 397 1813
rect 268 1803 277 1806
rect 394 1803 420 1806
rect 436 1803 453 1806
rect 458 1803 500 1806
rect 522 1803 572 1806
rect 690 1793 693 1823
rect 698 1813 706 1816
rect 756 1813 781 1816
rect 796 1813 821 1816
rect 828 1813 837 1816
rect 858 1813 868 1816
rect 954 1813 988 1816
rect 1020 1813 1037 1816
rect 1042 1813 1052 1816
rect 1122 1815 1125 1833
rect 1370 1816 1373 1836
rect 1842 1833 1852 1836
rect 1906 1833 1916 1836
rect 2010 1833 2036 1836
rect 2378 1826 2381 1836
rect 2450 1833 2469 1836
rect 2538 1833 2557 1836
rect 2450 1826 2453 1833
rect 1754 1823 1804 1826
rect 1900 1823 1909 1826
rect 1924 1823 1933 1826
rect 1948 1823 1957 1826
rect 2002 1823 2020 1826
rect 2340 1823 2381 1826
rect 2420 1823 2453 1826
rect 2484 1823 2493 1826
rect 2490 1816 2493 1823
rect 1194 1813 1204 1816
rect 1226 1813 1252 1816
rect 1300 1813 1309 1816
rect 1340 1813 1373 1816
rect 1388 1813 1396 1816
rect 1428 1813 1437 1816
rect 1500 1813 1517 1816
rect 1666 1813 1701 1816
rect 1940 1813 1957 1816
rect 1962 1813 1996 1816
rect 2236 1813 2253 1816
rect 698 1812 701 1813
rect 730 1803 748 1806
rect 788 1803 797 1806
rect 810 1803 820 1806
rect 884 1803 901 1806
rect 940 1803 957 1806
rect 986 1803 996 1806
rect 1012 1803 1021 1806
rect 1050 1803 1060 1806
rect 1180 1803 1189 1806
rect 1226 1803 1229 1813
rect 1306 1806 1309 1813
rect 1514 1806 1517 1813
rect 1268 1803 1285 1806
rect 1306 1803 1317 1806
rect 1346 1803 1380 1806
rect 1420 1803 1469 1806
rect 1492 1803 1509 1806
rect 1514 1803 1532 1806
rect 1548 1803 1581 1806
rect 1586 1803 1596 1806
rect 1634 1803 1644 1806
rect 1698 1805 1701 1813
rect 1714 1803 1717 1813
rect 1746 1806 1749 1813
rect 1746 1803 1757 1806
rect 1810 1803 1813 1813
rect 1906 1803 1909 1813
rect 1970 1803 1988 1806
rect 2164 1803 2173 1806
rect 2178 1803 2212 1806
rect 2228 1803 2237 1806
rect 2250 1803 2253 1813
rect 2314 1813 2332 1816
rect 2338 1813 2388 1816
rect 2394 1813 2411 1816
rect 2490 1813 2501 1816
rect 2508 1813 2533 1816
rect 2554 1815 2557 1833
rect 2572 1823 2581 1826
rect 2612 1823 2621 1826
rect 2610 1813 2621 1816
rect 2706 1813 2716 1816
rect 2890 1813 2908 1816
rect 2938 1813 2956 1816
rect 2988 1813 3005 1816
rect 3074 1813 3092 1816
rect 3122 1813 3148 1816
rect 2314 1806 2317 1813
rect 2258 1803 2284 1806
rect 2300 1803 2317 1806
rect 2578 1803 2588 1806
rect 770 1793 780 1796
rect 178 1783 189 1786
rect 274 1783 325 1786
rect 954 1783 957 1803
rect 1162 1793 1172 1796
rect 1314 1795 1317 1803
rect 2578 1793 2581 1803
rect 2618 1793 2621 1813
rect 2676 1803 2685 1806
rect 2698 1803 2708 1806
rect 2740 1803 2781 1806
rect 2804 1803 2813 1806
rect 2834 1803 2860 1806
rect 2890 1803 2893 1813
rect 3234 1806 3237 1815
rect 3300 1813 3333 1816
rect 3348 1813 3357 1816
rect 3364 1813 3397 1816
rect 2930 1803 2964 1806
rect 2980 1803 3013 1806
rect 3074 1803 3084 1806
rect 3130 1803 3140 1806
rect 3234 1803 3292 1806
rect 3298 1803 3340 1806
rect 3354 1805 3357 1813
rect 3210 1793 3220 1796
rect 3258 1793 3284 1796
rect 38 1767 3466 1773
rect 378 1743 388 1746
rect 650 1736 653 1756
rect 2162 1753 2181 1756
rect 850 1743 875 1746
rect 898 1736 901 1746
rect 1148 1743 1173 1746
rect 1170 1736 1173 1743
rect 130 1726 133 1736
rect 194 1733 220 1736
rect 250 1726 253 1736
rect 554 1733 564 1736
rect 594 1733 628 1736
rect 650 1733 669 1736
rect 682 1733 724 1736
rect 124 1723 157 1726
rect 180 1723 205 1726
rect 250 1723 300 1726
rect 450 1723 500 1726
rect 524 1723 541 1726
rect 412 1713 421 1716
rect 410 1703 428 1706
rect 554 1703 557 1733
rect 770 1726 773 1736
rect 858 1733 884 1736
rect 898 1733 940 1736
rect 1026 1733 1060 1736
rect 1170 1733 1180 1736
rect 1226 1726 1229 1746
rect 2522 1743 2541 1746
rect 3226 1743 3252 1746
rect 1234 1733 1276 1736
rect 1450 1733 1476 1736
rect 1636 1733 1653 1736
rect 1722 1733 1732 1736
rect 1762 1733 1773 1736
rect 1858 1733 1877 1736
rect 1900 1733 1909 1736
rect 1948 1733 1965 1736
rect 2026 1733 2036 1736
rect 2090 1733 2108 1736
rect 2154 1733 2188 1736
rect 2290 1733 2300 1736
rect 2372 1733 2389 1736
rect 2402 1733 2428 1736
rect 2458 1733 2492 1736
rect 2516 1733 2533 1736
rect 1770 1726 1773 1733
rect 636 1723 653 1726
rect 698 1723 714 1726
rect 770 1723 796 1726
rect 802 1723 837 1726
rect 852 1723 877 1726
rect 978 1723 1004 1726
rect 1210 1723 1220 1726
rect 1226 1723 1284 1726
rect 1500 1723 1509 1726
rect 1610 1723 1620 1726
rect 1634 1723 1676 1726
rect 1756 1723 1765 1726
rect 1770 1723 1788 1726
rect 1826 1723 1829 1733
rect 1836 1723 1869 1726
rect 1874 1725 1877 1733
rect 1908 1723 1925 1726
rect 644 1713 653 1716
rect 698 1683 701 1723
rect 1372 1713 1389 1716
rect 1412 1713 1421 1716
rect 1436 1713 1453 1716
rect 1506 1713 1516 1716
rect 1796 1713 1805 1716
rect 1844 1713 1861 1716
rect 1506 1693 1509 1713
rect 1522 1703 1532 1706
rect 1954 1703 1957 1726
rect 1962 1703 1965 1733
rect 2018 1723 2028 1726
rect 2060 1723 2101 1726
rect 2106 1723 2116 1726
rect 2122 1723 2140 1726
rect 2196 1723 2228 1726
rect 2260 1723 2306 1726
rect 2330 1723 2348 1726
rect 2386 1723 2420 1726
rect 2452 1723 2477 1726
rect 2500 1723 2509 1726
rect 1980 1713 1989 1716
rect 2004 1713 2013 1716
rect 2124 1713 2133 1716
rect 2148 1713 2189 1716
rect 2204 1713 2221 1716
rect 2316 1713 2341 1716
rect 1978 1703 1996 1706
rect 2010 1703 2013 1713
rect 2538 1706 2541 1743
rect 2554 1733 2564 1736
rect 2642 1733 2652 1736
rect 2706 1733 2724 1736
rect 2770 1733 2796 1736
rect 2852 1733 2861 1736
rect 2924 1733 2933 1736
rect 2994 1733 3036 1736
rect 3052 1733 3069 1736
rect 3082 1733 3108 1736
rect 3154 1733 3164 1736
rect 3220 1733 3229 1736
rect 2562 1723 2572 1726
rect 2698 1723 2732 1726
rect 2818 1723 2829 1726
rect 2882 1723 2900 1726
rect 2946 1723 2964 1726
rect 2996 1723 3005 1726
rect 3010 1723 3028 1726
rect 3060 1723 3085 1726
rect 3138 1723 3172 1726
rect 2578 1713 2588 1716
rect 2818 1715 2821 1723
rect 2852 1713 2893 1716
rect 2538 1703 2549 1706
rect 2578 1703 2604 1706
rect 2578 1693 2581 1703
rect 14 1667 3490 1673
rect 354 1633 380 1636
rect 348 1623 357 1626
rect 388 1623 397 1626
rect 530 1623 549 1626
rect 652 1623 661 1626
rect 692 1623 717 1626
rect 116 1613 125 1616
rect 164 1614 173 1616
rect 122 1606 125 1613
rect 162 1613 173 1614
rect 236 1613 261 1616
rect 306 1613 340 1616
rect 162 1606 165 1613
rect 394 1606 397 1623
rect 538 1616 541 1623
rect 658 1616 661 1623
rect 714 1616 717 1623
rect 778 1616 781 1625
rect 882 1616 885 1625
rect 1132 1623 1141 1626
rect 1298 1623 1308 1626
rect 1332 1623 1349 1626
rect 1434 1616 1437 1646
rect 2066 1636 2069 1656
rect 1506 1633 1539 1636
rect 1626 1633 1660 1636
rect 2066 1633 2085 1636
rect 2170 1633 2197 1636
rect 2258 1633 2285 1636
rect 2418 1633 2468 1636
rect 2618 1633 2653 1636
rect 2834 1633 2860 1636
rect 2970 1633 2980 1636
rect 1524 1623 1533 1626
rect 1548 1623 1581 1626
rect 1626 1623 1644 1626
rect 1674 1623 1701 1626
rect 1860 1623 1901 1626
rect 452 1613 461 1616
rect 474 1613 492 1616
rect 524 1613 533 1616
rect 538 1613 555 1616
rect 588 1613 605 1616
rect 658 1613 669 1616
rect 714 1613 725 1616
rect 732 1613 749 1616
rect 778 1613 789 1616
rect 882 1613 893 1616
rect 978 1613 1020 1616
rect 1114 1613 1124 1616
rect 1434 1613 1468 1616
rect 1562 1613 1581 1616
rect 1620 1613 1637 1616
rect 82 1603 100 1606
rect 122 1603 133 1606
rect 162 1603 212 1606
rect 250 1603 276 1606
rect 306 1603 332 1606
rect 394 1603 428 1606
rect 554 1603 564 1606
rect 580 1603 589 1606
rect 692 1603 709 1606
rect 722 1605 725 1613
rect 786 1606 789 1613
rect 738 1603 756 1606
rect 786 1603 796 1606
rect 818 1603 860 1606
rect 916 1603 925 1606
rect 946 1603 956 1606
rect 980 1603 997 1606
rect 1002 1603 1011 1606
rect 1074 1603 1100 1606
rect 1194 1603 1204 1606
rect 1228 1603 1245 1606
rect 1266 1603 1284 1606
rect 1338 1603 1364 1606
rect 1428 1603 1469 1606
rect 1562 1603 1596 1606
rect 1612 1603 1621 1606
rect 116 1593 125 1596
rect 1170 1593 1180 1596
rect 1194 1593 1197 1603
rect 1674 1596 1677 1623
rect 1724 1613 1733 1616
rect 1778 1613 1804 1616
rect 1852 1613 1885 1616
rect 2002 1613 2012 1616
rect 2044 1613 2053 1616
rect 2138 1613 2156 1616
rect 2194 1615 2197 1633
rect 2218 1613 2252 1616
rect 2282 1615 2285 1633
rect 2618 1626 2621 1633
rect 2300 1623 2309 1626
rect 2364 1623 2373 1626
rect 2412 1623 2429 1626
rect 2434 1623 2451 1626
rect 2330 1613 2348 1616
rect 1682 1603 1716 1606
rect 1722 1603 1732 1606
rect 1802 1603 1812 1606
rect 1834 1603 1844 1606
rect 1906 1603 1916 1606
rect 1956 1603 2013 1606
rect 2066 1603 2124 1606
rect 2314 1603 2340 1606
rect 2482 1603 2485 1626
rect 2596 1623 2621 1626
rect 2626 1623 2644 1626
rect 2762 1623 2788 1626
rect 2812 1623 2844 1626
rect 2626 1616 2629 1623
rect 2556 1613 2580 1616
rect 2610 1613 2629 1616
rect 2708 1613 2725 1616
rect 2898 1613 2956 1616
rect 3026 1613 3036 1616
rect 3060 1613 3069 1616
rect 3148 1613 3173 1616
rect 3204 1613 3237 1616
rect 3372 1613 3397 1616
rect 2522 1603 2548 1606
rect 2562 1603 2572 1606
rect 2674 1603 2700 1606
rect 2706 1603 2773 1606
rect 2874 1603 2884 1606
rect 2906 1603 2948 1606
rect 3042 1603 3052 1606
rect 3218 1603 3244 1606
rect 3316 1603 3325 1606
rect 1674 1593 1685 1596
rect 2106 1593 2116 1596
rect 2418 1593 2437 1596
rect 2674 1593 2692 1596
rect 2722 1593 2740 1596
rect 122 1583 125 1593
rect 38 1567 3466 1573
rect 378 1553 397 1556
rect 450 1543 468 1546
rect 130 1533 140 1536
rect 330 1533 348 1536
rect 386 1533 413 1536
rect 548 1533 565 1536
rect 74 1513 100 1516
rect 74 1496 77 1513
rect 106 1506 109 1525
rect 138 1523 148 1526
rect 252 1523 285 1526
rect 356 1523 381 1526
rect 386 1516 389 1533
rect 444 1523 461 1526
rect 506 1523 524 1526
rect 124 1513 133 1516
rect 156 1513 173 1516
rect 378 1513 389 1516
rect 82 1503 109 1506
rect 266 1503 316 1506
rect 562 1496 565 1533
rect 602 1526 605 1556
rect 1802 1553 1813 1556
rect 922 1543 972 1546
rect 1266 1543 1308 1546
rect 732 1533 749 1536
rect 898 1533 916 1536
rect 1068 1533 1093 1536
rect 1130 1533 1140 1536
rect 1260 1533 1277 1536
rect 1316 1533 1333 1536
rect 1370 1533 1396 1536
rect 682 1523 716 1526
rect 802 1523 828 1526
rect 924 1523 933 1526
rect 1012 1523 1029 1526
rect 1130 1523 1148 1526
rect 1210 1523 1220 1526
rect 1268 1523 1293 1526
rect 1394 1523 1404 1526
rect 1490 1516 1493 1536
rect 1516 1533 1525 1536
rect 1634 1533 1644 1536
rect 1626 1523 1652 1526
rect 1802 1516 1805 1553
rect 2058 1543 2068 1546
rect 2746 1543 2756 1546
rect 1860 1533 1885 1536
rect 1930 1533 1964 1536
rect 1980 1533 1989 1536
rect 2058 1533 2076 1536
rect 2082 1533 2116 1536
rect 2178 1533 2188 1536
rect 2218 1533 2244 1536
rect 2260 1533 2293 1536
rect 2306 1533 2316 1536
rect 2218 1526 2221 1533
rect 2402 1526 2405 1534
rect 1810 1523 1853 1526
rect 2084 1523 2101 1526
rect 2154 1523 2196 1526
rect 2210 1523 2221 1526
rect 2268 1523 2277 1526
rect 2306 1523 2324 1526
rect 2338 1523 2405 1526
rect 668 1513 701 1516
rect 738 1513 764 1516
rect 788 1513 821 1516
rect 836 1513 868 1516
rect 1068 1513 1077 1516
rect 1420 1513 1437 1516
rect 1444 1513 1453 1516
rect 1468 1513 1493 1516
rect 1562 1513 1596 1516
rect 1668 1513 1685 1516
rect 1708 1513 1717 1516
rect 1732 1513 1749 1516
rect 1780 1513 1789 1516
rect 1802 1513 1813 1516
rect 2020 1513 2029 1516
rect 2044 1513 2053 1516
rect 2154 1513 2157 1523
rect 2490 1516 2493 1534
rect 2506 1533 2516 1536
rect 2578 1533 2604 1536
rect 2676 1533 2701 1536
rect 2706 1526 2709 1534
rect 2732 1533 2741 1536
rect 2770 1533 2804 1536
rect 2828 1533 2837 1536
rect 2850 1533 2860 1536
rect 2866 1533 2900 1536
rect 2930 1533 2956 1536
rect 2514 1523 2524 1526
rect 2572 1523 2597 1526
rect 2602 1523 2612 1526
rect 2674 1523 2709 1526
rect 2866 1525 2869 1533
rect 2978 1526 2981 1534
rect 3098 1533 3108 1536
rect 3250 1533 3284 1536
rect 3314 1526 3317 1534
rect 3362 1533 3372 1536
rect 3402 1526 3405 1534
rect 2978 1523 2989 1526
rect 3116 1523 3141 1526
rect 3244 1523 3269 1526
rect 3308 1523 3317 1526
rect 3396 1523 3405 1526
rect 3412 1523 3421 1526
rect 2602 1516 2605 1523
rect 2340 1513 2349 1516
rect 2364 1513 2373 1516
rect 2482 1513 2493 1516
rect 2508 1513 2517 1516
rect 2586 1513 2605 1516
rect 2620 1513 2637 1516
rect 2828 1513 2837 1516
rect 2986 1506 2989 1523
rect 3004 1513 3013 1516
rect 3034 1513 3068 1516
rect 570 1503 612 1506
rect 1762 1503 1772 1506
rect 2018 1503 2036 1506
rect 2986 1503 3020 1506
rect 74 1493 85 1496
rect 562 1493 573 1496
rect 14 1467 3490 1473
rect 314 1433 340 1436
rect 522 1433 549 1436
rect 714 1433 733 1436
rect 1290 1433 1325 1436
rect 2002 1433 2021 1436
rect 2146 1433 2164 1436
rect 2242 1433 2268 1436
rect 2322 1433 2356 1436
rect 2978 1433 3037 1436
rect 714 1426 717 1433
rect 146 1416 149 1426
rect 164 1423 205 1426
rect 228 1423 237 1426
rect 348 1423 365 1426
rect 381 1423 413 1426
rect 474 1416 477 1426
rect 522 1423 541 1426
rect 594 1423 612 1426
rect 636 1423 645 1426
rect 708 1423 717 1426
rect 538 1416 541 1423
rect 138 1413 156 1416
rect 210 1413 220 1416
rect 138 1406 141 1413
rect 82 1403 108 1406
rect 124 1403 141 1406
rect 274 1406 277 1414
rect 354 1413 372 1416
rect 378 1413 413 1416
rect 452 1413 477 1416
rect 516 1413 533 1416
rect 538 1413 555 1416
rect 274 1403 301 1406
rect 354 1403 364 1406
rect 514 1403 564 1406
rect 298 1393 301 1403
rect 386 1393 405 1396
rect 618 1393 621 1414
rect 770 1413 804 1416
rect 666 1403 684 1406
rect 826 1405 829 1426
rect 844 1423 869 1426
rect 1124 1423 1141 1426
rect 1290 1416 1293 1433
rect 1380 1423 1389 1426
rect 1628 1423 1661 1426
rect 1794 1423 1821 1426
rect 1860 1423 1917 1426
rect 1996 1423 2005 1426
rect 922 1413 940 1416
rect 978 1413 988 1416
rect 1066 1413 1108 1416
rect 1164 1413 1173 1416
rect 1212 1413 1237 1416
rect 1258 1413 1269 1416
rect 1276 1413 1293 1416
rect 1330 1413 1340 1416
rect 1354 1413 1365 1416
rect 1372 1413 1381 1416
rect 1018 1403 1036 1406
rect 1074 1403 1100 1406
rect 1130 1403 1156 1406
rect 1162 1403 1204 1406
rect 1210 1403 1236 1406
rect 1258 1405 1261 1413
rect 1282 1403 1332 1406
rect 1362 1405 1365 1413
rect 916 1393 925 1396
rect 1186 1393 1196 1396
rect 522 1383 549 1386
rect 1386 1383 1389 1423
rect 1394 1413 1436 1416
rect 1556 1413 1565 1416
rect 1572 1413 1612 1416
rect 1754 1413 1772 1416
rect 1794 1406 1797 1423
rect 1802 1413 1828 1416
rect 1418 1403 1428 1406
rect 1538 1403 1548 1406
rect 1554 1403 1564 1406
rect 1578 1403 1604 1406
rect 1634 1403 1676 1406
rect 1724 1403 1764 1406
rect 1788 1403 1797 1406
rect 2018 1406 2021 1433
rect 2052 1423 2069 1426
rect 2130 1423 2148 1426
rect 2220 1423 2237 1426
rect 2242 1416 2245 1433
rect 2276 1423 2285 1426
rect 2108 1413 2125 1416
rect 2186 1413 2204 1416
rect 2234 1413 2245 1416
rect 2018 1403 2028 1406
rect 2082 1403 2092 1406
rect 2186 1403 2196 1406
rect 1650 1393 1668 1396
rect 1698 1393 1716 1396
rect 2108 1393 2125 1396
rect 2282 1383 2285 1423
rect 2322 1416 2325 1433
rect 2330 1423 2340 1426
rect 2746 1423 2765 1426
rect 2994 1423 3028 1426
rect 2746 1416 2749 1423
rect 2316 1413 2325 1416
rect 2370 1413 2396 1416
rect 2410 1413 2428 1416
rect 2452 1413 2461 1416
rect 2466 1413 2500 1416
rect 2506 1406 2509 1416
rect 2524 1413 2565 1416
rect 2652 1413 2669 1416
rect 2674 1413 2700 1416
rect 2732 1413 2749 1416
rect 2754 1413 2780 1416
rect 2820 1413 2837 1416
rect 2842 1413 2860 1416
rect 2908 1413 2956 1416
rect 3034 1415 3037 1433
rect 3058 1426 3061 1436
rect 3052 1423 3061 1426
rect 3348 1423 3365 1426
rect 3100 1413 3133 1416
rect 3180 1413 3189 1416
rect 3276 1413 3332 1416
rect 2754 1406 2757 1413
rect 2290 1403 2308 1406
rect 2370 1403 2388 1406
rect 2402 1403 2436 1406
rect 2466 1403 2492 1406
rect 2506 1403 2516 1406
rect 2538 1403 2580 1406
rect 2618 1403 2636 1406
rect 2650 1403 2708 1406
rect 2724 1403 2757 1406
rect 2762 1403 2772 1406
rect 2794 1403 2852 1406
rect 2866 1403 2892 1406
rect 2922 1403 2948 1406
rect 2972 1403 2989 1406
rect 3058 1403 3092 1406
rect 3172 1403 3189 1406
rect 3250 1403 3268 1406
rect 3354 1403 3372 1406
rect 2452 1393 2461 1396
rect 2762 1393 2765 1403
rect 3058 1393 3084 1396
rect 3106 1383 3157 1386
rect 38 1367 3466 1373
rect 338 1353 365 1356
rect 682 1353 693 1356
rect 2602 1353 2629 1356
rect 386 1336 389 1346
rect 82 1333 92 1336
rect 164 1333 213 1336
rect 386 1333 397 1336
rect 514 1333 564 1336
rect 580 1333 597 1336
rect 66 1323 100 1326
rect 172 1323 197 1326
rect 282 1323 300 1326
rect 381 1323 389 1326
rect 394 1325 397 1333
rect 420 1323 429 1326
rect 546 1323 555 1326
rect 252 1313 269 1316
rect 594 1313 597 1333
rect 618 1323 636 1326
rect 682 1316 685 1353
rect 1242 1343 1260 1346
rect 1378 1343 1404 1346
rect 1242 1336 1245 1343
rect 834 1333 844 1336
rect 882 1333 900 1336
rect 922 1333 932 1336
rect 978 1333 1020 1336
rect 1052 1333 1069 1336
rect 1098 1333 1132 1336
rect 1212 1333 1245 1336
rect 1458 1336 1461 1346
rect 1676 1343 1709 1346
rect 1458 1333 1476 1336
rect 1508 1333 1525 1336
rect 1610 1333 1660 1336
rect 1748 1333 1757 1336
rect 882 1326 885 1333
rect 730 1323 740 1326
rect 852 1323 885 1326
rect 930 1323 940 1326
rect 970 1323 1028 1326
rect 1084 1323 1093 1326
rect 1140 1323 1149 1326
rect 1162 1323 1181 1326
rect 1282 1323 1292 1326
rect 1322 1323 1356 1326
rect 1362 1323 1372 1326
rect 1450 1323 1484 1326
rect 1554 1323 1572 1326
rect 1634 1323 1652 1326
rect 1722 1323 1732 1326
rect 1802 1325 1805 1346
rect 1906 1343 1948 1346
rect 1986 1343 2020 1346
rect 2154 1336 2157 1346
rect 2442 1343 2468 1346
rect 1834 1333 1868 1336
rect 1930 1333 1956 1336
rect 2018 1333 2028 1336
rect 2034 1333 2044 1336
rect 2106 1333 2116 1336
rect 2154 1333 2204 1336
rect 2306 1333 2324 1336
rect 2348 1333 2365 1336
rect 2386 1333 2396 1336
rect 2434 1333 2476 1336
rect 2482 1333 2501 1336
rect 2522 1333 2532 1336
rect 2570 1333 2588 1336
rect 1866 1323 1876 1326
rect 2036 1323 2093 1326
rect 2186 1323 2196 1326
rect 2234 1323 2268 1326
rect 2346 1323 2404 1326
rect 652 1313 685 1316
rect 690 1313 700 1316
rect 794 1313 804 1316
rect 1796 1313 1805 1316
rect 202 1303 244 1306
rect 706 1303 716 1306
rect 2186 1293 2189 1323
rect 2284 1313 2309 1316
rect 2498 1313 2501 1333
rect 2578 1323 2596 1326
rect 2602 1316 2605 1353
rect 2738 1346 2741 1356
rect 2682 1343 2716 1346
rect 2738 1343 2764 1346
rect 2858 1343 2877 1346
rect 2858 1336 2861 1343
rect 2610 1333 2636 1336
rect 2724 1333 2749 1336
rect 2762 1333 2812 1336
rect 2844 1333 2861 1336
rect 2866 1333 2892 1336
rect 2930 1333 2972 1336
rect 2986 1333 3020 1336
rect 3050 1326 3053 1335
rect 3306 1333 3340 1336
rect 3370 1333 3388 1336
rect 2626 1323 2644 1326
rect 2676 1323 2693 1326
rect 2732 1323 2741 1326
rect 2780 1323 2789 1326
rect 2866 1323 2900 1326
rect 2930 1323 2964 1326
rect 2988 1323 3028 1326
rect 3042 1323 3053 1326
rect 3060 1323 3077 1326
rect 3132 1323 3149 1326
rect 3210 1323 3220 1326
rect 3330 1323 3341 1326
rect 3378 1323 3396 1326
rect 3330 1316 3333 1323
rect 3378 1316 3381 1323
rect 2602 1313 2621 1316
rect 3308 1313 3333 1316
rect 3364 1313 3381 1316
rect 1306 1283 1341 1286
rect 14 1267 3490 1273
rect 266 1243 277 1246
rect 218 1233 244 1236
rect 266 1226 269 1243
rect 274 1233 308 1236
rect 618 1233 637 1236
rect 858 1233 876 1236
rect 116 1223 141 1226
rect 172 1223 189 1226
rect 202 1223 228 1226
rect 252 1223 269 1226
rect 316 1223 333 1226
rect 410 1223 437 1226
rect 90 1203 100 1206
rect 138 1203 148 1206
rect 186 1203 189 1223
rect 410 1216 413 1223
rect 466 1216 469 1224
rect 354 1213 372 1216
rect 404 1213 413 1216
rect 418 1213 460 1216
rect 466 1213 477 1216
rect 484 1213 501 1216
rect 506 1213 548 1216
rect 634 1215 637 1233
rect 722 1216 725 1225
rect 788 1223 797 1226
rect 834 1223 860 1226
rect 1396 1223 1421 1226
rect 658 1213 716 1216
rect 722 1213 740 1216
rect 930 1213 940 1216
rect 1076 1213 1085 1216
rect 1162 1213 1172 1216
rect 1324 1213 1373 1216
rect 338 1203 380 1206
rect 396 1203 445 1206
rect 514 1203 555 1206
rect 572 1203 589 1206
rect 666 1203 708 1206
rect 722 1203 732 1206
rect 914 1203 932 1206
rect 1036 1203 1045 1206
rect 1098 1203 1140 1206
rect 1268 1203 1293 1206
rect 1298 1203 1316 1206
rect 1370 1205 1373 1213
rect 1402 1213 1436 1216
rect 1290 1196 1293 1203
rect 1402 1196 1405 1213
rect 1410 1203 1444 1206
rect 1490 1196 1493 1216
rect 1516 1213 1525 1216
rect 1540 1213 1557 1216
rect 1562 1213 1596 1216
rect 1634 1206 1637 1236
rect 1770 1233 1813 1236
rect 3146 1233 3180 1236
rect 3250 1233 3276 1236
rect 3354 1233 3381 1236
rect 1498 1203 1508 1206
rect 1532 1203 1557 1206
rect 1578 1203 1597 1206
rect 1620 1203 1637 1206
rect 1642 1223 1661 1226
rect 1692 1223 1717 1226
rect 1722 1223 1732 1226
rect 1786 1223 1804 1226
rect 1018 1193 1028 1196
rect 1106 1193 1132 1196
rect 1290 1193 1308 1196
rect 1402 1193 1421 1196
rect 1460 1193 1493 1196
rect 1642 1196 1645 1223
rect 1722 1216 1725 1223
rect 1658 1213 1676 1216
rect 1714 1213 1725 1216
rect 1810 1215 1813 1233
rect 1948 1223 1981 1226
rect 2012 1223 2021 1226
rect 2060 1223 2069 1226
rect 2196 1223 2221 1226
rect 2332 1223 2341 1226
rect 3218 1223 3260 1226
rect 3284 1223 3293 1226
rect 2338 1216 2341 1223
rect 3354 1216 3357 1233
rect 3362 1223 3372 1226
rect 1850 1213 1876 1216
rect 1898 1213 1932 1216
rect 1978 1213 1996 1216
rect 2010 1213 2093 1216
rect 2132 1213 2165 1216
rect 2188 1213 2221 1216
rect 2090 1206 2093 1213
rect 2226 1206 2229 1215
rect 2260 1213 2269 1216
rect 2306 1213 2316 1216
rect 2338 1213 2349 1216
rect 2356 1213 2365 1216
rect 2490 1213 2508 1216
rect 2546 1213 2596 1216
rect 2652 1213 2669 1216
rect 2756 1213 2765 1216
rect 2868 1213 2901 1216
rect 2932 1213 2949 1216
rect 3108 1213 3117 1216
rect 3324 1213 3357 1216
rect 3378 1215 3381 1233
rect 2546 1206 2549 1213
rect 1650 1203 1668 1206
rect 1692 1203 1701 1206
rect 1892 1203 1901 1206
rect 1948 1203 1973 1206
rect 2012 1203 2037 1206
rect 2090 1203 2101 1206
rect 2130 1203 2180 1206
rect 2194 1203 2229 1206
rect 2258 1203 2308 1206
rect 2332 1203 2341 1206
rect 2412 1203 2429 1206
rect 2444 1203 2461 1206
rect 2466 1203 2493 1206
rect 2522 1203 2532 1206
rect 2538 1203 2549 1206
rect 2676 1203 2701 1206
rect 2772 1203 2821 1206
rect 2836 1203 2853 1206
rect 2860 1203 2869 1206
rect 2930 1203 2956 1206
rect 2988 1203 2997 1206
rect 3002 1203 3036 1206
rect 3060 1203 3069 1206
rect 3074 1203 3092 1206
rect 3298 1203 3316 1206
rect 1642 1193 1653 1196
rect 1698 1193 1701 1203
rect 2362 1193 2404 1196
rect 2690 1193 2740 1196
rect 2810 1193 2828 1196
rect 2842 1193 2852 1196
rect 2874 1193 2916 1196
rect 3108 1193 3117 1196
rect 38 1167 3466 1173
rect 506 1153 525 1156
rect 850 1146 853 1156
rect 130 1143 141 1146
rect 290 1143 301 1146
rect 556 1143 565 1146
rect 844 1143 853 1146
rect 954 1143 980 1146
rect 1146 1143 1164 1146
rect 1514 1143 1533 1146
rect 1810 1143 1852 1146
rect 130 1126 133 1143
rect 138 1133 156 1136
rect 170 1133 196 1136
rect 210 1133 252 1136
rect 268 1133 293 1136
rect 66 1123 92 1126
rect 130 1123 164 1126
rect 170 1123 204 1126
rect 276 1123 293 1126
rect 172 1113 189 1116
rect 290 1113 293 1123
rect 298 1116 301 1143
rect 404 1133 413 1136
rect 450 1133 460 1136
rect 476 1133 501 1136
rect 570 1133 580 1136
rect 658 1133 676 1136
rect 714 1133 724 1136
rect 754 1133 772 1136
rect 802 1133 828 1136
rect 858 1133 884 1136
rect 898 1133 948 1136
rect 954 1133 988 1136
rect 1002 1133 1036 1136
rect 1146 1133 1172 1136
rect 1242 1133 1260 1136
rect 1362 1133 1372 1136
rect 1410 1133 1444 1136
rect 754 1126 757 1133
rect 802 1126 805 1133
rect 362 1123 380 1126
rect 418 1123 452 1126
rect 484 1123 493 1126
rect 514 1123 532 1126
rect 556 1123 581 1126
rect 588 1123 613 1126
rect 362 1116 365 1123
rect 298 1113 308 1116
rect 332 1113 365 1116
rect 418 1113 421 1123
rect 610 1106 613 1123
rect 634 1106 637 1125
rect 658 1123 684 1126
rect 690 1123 732 1126
rect 746 1123 757 1126
rect 770 1123 805 1126
rect 810 1123 820 1126
rect 844 1123 853 1126
rect 956 1123 973 1126
rect 1018 1123 1044 1126
rect 1180 1123 1221 1126
rect 1226 1123 1236 1126
rect 1396 1123 1405 1126
rect 1434 1123 1452 1126
rect 1226 1116 1229 1123
rect 1514 1116 1517 1143
rect 1530 1136 1533 1143
rect 1522 1126 1525 1136
rect 1530 1133 1540 1136
rect 1602 1133 1611 1136
rect 1636 1133 1676 1136
rect 1690 1133 1708 1136
rect 1738 1133 1772 1136
rect 1788 1133 1853 1136
rect 1860 1133 1885 1136
rect 1900 1133 1909 1136
rect 1914 1126 1917 1146
rect 1986 1143 1996 1146
rect 2898 1143 2932 1146
rect 2962 1143 2972 1146
rect 2004 1133 2021 1136
rect 2098 1133 2108 1136
rect 2234 1126 2237 1136
rect 2258 1133 2284 1136
rect 2306 1133 2316 1136
rect 2338 1133 2380 1136
rect 2404 1133 2421 1136
rect 2434 1133 2452 1136
rect 2474 1133 2540 1136
rect 2554 1133 2564 1136
rect 2626 1133 2636 1136
rect 2690 1133 2748 1136
rect 2754 1133 2828 1136
rect 2940 1133 2973 1136
rect 3026 1133 3036 1136
rect 3058 1133 3068 1136
rect 3092 1133 3140 1136
rect 2338 1126 2341 1133
rect 1522 1123 1548 1126
rect 1578 1123 1620 1126
rect 1658 1123 1684 1126
rect 1698 1123 1716 1126
rect 1746 1123 1764 1126
rect 1908 1123 1917 1126
rect 1938 1123 1964 1126
rect 2012 1123 2061 1126
rect 652 1113 669 1116
rect 748 1113 757 1116
rect 1194 1113 1229 1116
rect 1306 1113 1316 1116
rect 1340 1113 1349 1116
rect 1484 1113 1493 1116
rect 1514 1113 1525 1116
rect 2034 1113 2068 1116
rect 2074 1106 2077 1125
rect 2116 1123 2141 1126
rect 2234 1123 2301 1126
rect 2324 1123 2341 1126
rect 2514 1123 2548 1126
rect 2666 1123 2741 1126
rect 2754 1125 2757 1133
rect 2788 1123 2805 1126
rect 2810 1123 2845 1126
rect 2092 1113 2101 1116
rect 2556 1113 2565 1116
rect 2580 1113 2597 1116
rect 2850 1113 2868 1116
rect 2874 1106 2877 1125
rect 3018 1123 3044 1126
rect 3162 1123 3180 1126
rect 3242 1123 3260 1126
rect 3290 1123 3333 1126
rect 3330 1116 3333 1123
rect 3092 1113 3125 1116
rect 3330 1113 3348 1116
rect 298 1103 324 1106
rect 594 1103 637 1106
rect 1322 1103 1332 1106
rect 2066 1103 2077 1106
rect 2122 1103 2188 1106
rect 2842 1103 2877 1106
rect 3378 1103 3396 1106
rect 14 1067 3490 1073
rect 2154 1053 2173 1056
rect 154 1023 173 1026
rect 268 1023 309 1026
rect 170 1016 173 1023
rect 562 1016 565 1046
rect 690 1033 701 1036
rect 1066 1033 1108 1036
rect 2098 1033 2133 1036
rect 2186 1033 2204 1036
rect 2346 1033 2365 1036
rect 2666 1033 2677 1036
rect 2682 1033 2716 1036
rect 2794 1033 2805 1036
rect 2842 1033 2860 1036
rect 2882 1033 2917 1036
rect 2978 1033 2996 1036
rect 652 1023 685 1026
rect 108 1013 117 1016
rect 132 1013 165 1016
rect 170 1013 188 1016
rect 234 1013 260 1016
rect 282 1013 324 1016
rect 418 1013 436 1016
rect 442 1013 460 1016
rect 532 1013 565 1016
rect 618 1013 636 1016
rect 698 1015 701 1033
rect 2098 1026 2101 1033
rect 780 1023 789 1026
rect 988 1023 1021 1026
rect 1116 1023 1141 1026
rect 2012 1023 2021 1026
rect 2084 1023 2101 1026
rect 2106 1023 2124 1026
rect 2148 1023 2181 1026
rect 2188 1023 2197 1026
rect 2212 1023 2237 1026
rect 2332 1023 2357 1026
rect 730 1013 764 1016
rect 810 1013 820 1016
rect 844 1013 853 1016
rect 898 1013 924 1016
rect 986 1013 1028 1016
rect 1282 1013 1317 1016
rect 1450 1013 1492 1016
rect 1516 1013 1525 1016
rect 1554 1013 1572 1016
rect 1780 1013 1789 1016
rect 1834 1013 1876 1016
rect 1898 1013 1924 1016
rect 1930 1013 1972 1016
rect 1978 1013 1996 1016
rect 2034 1013 2068 1016
rect 2082 1013 2101 1016
rect 2330 1013 2365 1016
rect 234 1006 237 1013
rect 114 1003 124 1006
rect 146 1003 165 1006
rect 170 1003 196 1006
rect 212 1003 237 1006
rect 266 1003 316 1006
rect 340 1003 357 1006
rect 364 1003 381 1006
rect 402 1003 428 1006
rect 594 1003 628 1006
rect 738 1003 756 1006
rect 780 1003 805 1006
rect 810 1003 828 1006
rect 858 1003 884 1006
rect 898 1003 916 1006
rect 938 1003 964 1006
rect 1178 1003 1212 1006
rect 1234 1003 1268 1006
rect 1274 1003 1292 1006
rect 474 993 492 996
rect 844 993 869 996
rect 898 993 901 1003
rect 1314 996 1317 1013
rect 2402 1006 2405 1014
rect 2490 1013 2516 1016
rect 1330 1003 1348 1006
rect 1388 1003 1413 1006
rect 1474 1003 1484 1006
rect 1508 1003 1517 1006
rect 1522 1003 1564 1006
rect 1610 1003 1652 1006
rect 1666 1003 1692 1006
rect 1738 1003 1764 1006
rect 1820 1003 1868 1006
rect 1978 1003 1988 1006
rect 2012 1003 2053 1006
rect 2218 1003 2244 1006
rect 2282 1003 2308 1006
rect 2332 1003 2341 1006
rect 2370 1003 2380 1006
rect 2402 1003 2452 1006
rect 2474 1003 2508 1006
rect 2522 1003 2525 1025
rect 2666 1016 2669 1033
rect 2674 1023 2700 1026
rect 2666 1013 2685 1016
rect 2802 1015 2805 1033
rect 2834 1023 2844 1026
rect 2874 1023 2908 1026
rect 2914 1015 2917 1033
rect 2980 1023 2989 1026
rect 3220 1023 3229 1026
rect 2946 1013 2972 1016
rect 3084 1013 3101 1016
rect 3194 1013 3204 1016
rect 3250 1013 3276 1016
rect 3306 1013 3332 1016
rect 2538 1003 2572 1006
rect 2594 1003 2636 1006
rect 2938 1003 2964 1006
rect 3220 1003 3268 1006
rect 3300 1003 3309 1006
rect 3314 1003 3340 1006
rect 3378 1003 3412 1006
rect 1514 996 1517 1003
rect 3306 996 3309 1003
rect 1052 993 1061 996
rect 1186 993 1204 996
rect 1314 993 1340 996
rect 1354 993 1380 996
rect 1514 993 1541 996
rect 1602 993 1644 996
rect 1780 993 1797 996
rect 1802 993 1812 996
rect 1826 993 1853 996
rect 3306 993 3325 996
rect 3394 993 3404 996
rect 1626 983 1629 993
rect 38 967 3466 973
rect 2234 946 2237 956
rect 194 943 220 946
rect 386 943 404 946
rect 898 943 916 946
rect 1258 943 1276 946
rect 1314 943 1372 946
rect 1626 943 1644 946
rect 1666 943 1708 946
rect 1906 943 1916 946
rect 2234 943 2261 946
rect 3210 943 3220 946
rect 82 933 108 936
rect 114 933 125 936
rect 164 933 181 936
rect 228 933 245 936
rect 290 933 300 936
rect 378 933 412 936
rect 498 933 524 936
rect 540 933 581 936
rect 778 933 796 936
rect 820 933 845 936
rect 890 933 924 936
rect 1034 933 1068 936
rect 1084 933 1093 936
rect 122 926 125 933
rect 242 926 245 933
rect 122 923 148 926
rect 242 923 253 926
rect 274 923 308 926
rect 428 923 437 926
rect 498 916 501 933
rect 548 923 565 926
rect 586 923 604 926
rect 730 923 740 926
rect 316 913 325 916
rect 338 913 348 916
rect 452 913 461 916
rect 476 913 501 916
rect 620 913 629 916
rect 666 913 700 916
rect 820 913 837 916
rect 626 906 629 913
rect 842 906 845 933
rect 932 923 941 926
rect 1002 923 1028 926
rect 1042 923 1060 926
rect 1092 923 1149 926
rect 1170 923 1173 935
rect 1258 933 1284 936
rect 1298 933 1308 936
rect 1322 933 1380 936
rect 1386 933 1396 936
rect 1498 933 1508 936
rect 1532 933 1573 936
rect 1578 933 1588 936
rect 1612 933 1621 936
rect 1634 933 1652 936
rect 1722 933 1732 936
rect 1770 933 1796 936
rect 1820 933 1853 936
rect 1962 933 1972 936
rect 1996 933 2013 936
rect 2042 933 2077 936
rect 2100 933 2109 936
rect 2138 933 2156 936
rect 2170 933 2189 936
rect 2212 933 2269 936
rect 2322 933 2388 936
rect 2404 933 2429 936
rect 2434 933 2444 936
rect 2466 933 2508 936
rect 2530 933 2557 936
rect 2594 933 2644 936
rect 2690 933 2700 936
rect 1570 926 1573 933
rect 1178 923 1204 926
rect 1394 923 1437 926
rect 1490 923 1516 926
rect 1570 923 1596 926
rect 1660 923 1685 926
rect 1778 923 1804 926
rect 1818 923 1829 926
rect 2036 923 2061 926
rect 2074 925 2077 933
rect 2108 923 2149 926
rect 2164 923 2181 926
rect 2186 925 2189 933
rect 2316 923 2325 926
rect 2370 923 2380 926
rect 2412 923 2421 926
rect 2452 923 2493 926
rect 2530 925 2533 933
rect 2730 926 2733 935
rect 3210 933 3228 936
rect 3258 933 3276 936
rect 2538 923 2564 926
rect 2596 923 2605 926
rect 2610 923 2636 926
rect 2722 923 2733 926
rect 1434 916 1437 923
rect 1826 916 1829 923
rect 2602 916 2605 923
rect 876 913 893 916
rect 980 913 989 916
rect 1172 913 1181 916
rect 1220 913 1245 916
rect 1434 913 1452 916
rect 1476 913 1501 916
rect 1532 913 1541 916
rect 1826 913 1860 916
rect 2044 913 2069 916
rect 2172 913 2181 916
rect 2242 913 2276 916
rect 2324 913 2333 916
rect 2602 913 2621 916
rect 2796 913 2805 916
rect 2898 913 2908 916
rect 2914 906 2917 925
rect 2938 923 2972 926
rect 2978 923 2996 926
rect 3002 923 3020 926
rect 3084 923 3109 926
rect 3250 923 3301 926
rect 3356 923 3389 926
rect 3298 916 3301 923
rect 3298 913 3316 916
rect 3386 906 3389 923
rect 3402 906 3405 925
rect 354 903 364 906
rect 442 903 468 906
rect 626 903 645 906
rect 842 903 853 906
rect 1442 903 1468 906
rect 1834 903 1876 906
rect 2234 903 2292 906
rect 2826 903 2868 906
rect 2882 903 2917 906
rect 3322 903 3332 906
rect 3386 903 3405 906
rect 14 867 3490 873
rect 738 853 757 856
rect 1130 853 1173 856
rect 226 833 284 836
rect 618 833 660 836
rect 826 833 836 836
rect 2242 833 2292 836
rect 268 823 277 826
rect 292 823 333 826
rect 644 823 653 826
rect 732 823 749 826
rect 786 823 820 826
rect 972 823 981 826
rect 1028 823 1061 826
rect 1260 823 1285 826
rect 1684 823 1725 826
rect 1932 823 1957 826
rect 2138 823 2156 826
rect 2180 823 2221 826
rect 2236 823 2253 826
rect 2258 823 2276 826
rect 2300 823 2333 826
rect 108 813 133 816
rect 140 813 181 816
rect 220 813 261 816
rect 372 813 405 816
rect 444 813 461 816
rect 466 813 492 816
rect 530 813 564 816
rect 690 813 716 816
rect 402 806 405 813
rect 746 806 749 823
rect 2258 816 2261 823
rect 2570 816 2573 826
rect 2892 823 2901 826
rect 2932 823 2965 826
rect 780 813 805 816
rect 850 813 884 816
rect 1034 813 1076 816
rect 1138 813 1188 816
rect 1242 813 1252 816
rect 1338 813 1388 816
rect 1482 813 1524 816
rect 1594 813 1612 816
rect 1626 813 1661 816
rect 1756 813 1773 816
rect 1796 813 1805 816
rect 1860 813 1901 816
rect 1946 813 1972 816
rect 2002 813 2036 816
rect 2090 813 2149 816
rect 2228 813 2237 816
rect 2242 813 2261 816
rect 2306 813 2340 816
rect 2362 813 2388 816
rect 2538 813 2548 816
rect 2570 813 2596 816
rect 2626 813 2684 816
rect 2708 813 2741 816
rect 2780 813 2805 816
rect 3004 813 3029 816
rect 3220 813 3245 816
rect 3292 813 3301 816
rect 3308 813 3317 816
rect 3332 813 3341 816
rect 3410 813 3420 816
rect 114 803 132 806
rect 170 803 196 806
rect 212 803 229 806
rect 330 803 348 806
rect 364 803 397 806
rect 402 803 420 806
rect 436 803 461 806
rect 516 803 572 806
rect 588 803 637 806
rect 732 803 741 806
rect 746 803 772 806
rect 866 803 876 806
rect 914 803 948 806
rect 1028 803 1037 806
rect 1042 803 1068 806
rect 1124 803 1149 806
rect 1258 803 1292 806
rect 1330 803 1380 806
rect 1418 803 1452 806
rect 1490 803 1516 806
rect 1548 803 1557 806
rect 1570 803 1604 806
rect 1626 805 1629 813
rect 1634 803 1660 806
rect 1684 803 1709 806
rect 1714 803 1748 806
rect 1754 803 1788 806
rect 1810 803 1844 806
rect 1938 803 1964 806
rect 1988 803 2013 806
rect 2018 803 2028 806
rect 2082 803 2108 806
rect 2186 803 2220 806
rect 2386 803 2396 806
rect 2410 803 2420 806
rect 2450 803 2492 806
rect 2690 803 2700 806
rect 2842 803 2868 806
rect 3066 803 3084 806
rect 3154 803 3196 806
rect 3202 803 3212 806
rect 3258 803 3284 806
rect 394 796 397 803
rect 394 793 405 796
rect 754 793 764 796
rect 682 783 701 786
rect 1146 783 1149 803
rect 1706 796 1709 803
rect 2018 796 2021 803
rect 1706 793 1725 796
rect 1730 793 1740 796
rect 1860 793 1869 796
rect 2002 793 2021 796
rect 3162 793 3188 796
rect 3258 793 3276 796
rect 3314 795 3317 813
rect 3338 803 3388 806
rect 1730 786 1733 793
rect 1690 783 1733 786
rect 38 767 3466 773
rect 1306 746 1309 756
rect 730 743 748 746
rect 1066 743 1132 746
rect 1300 743 1309 746
rect 1490 743 1516 746
rect 3148 743 3157 746
rect 82 733 92 736
rect 132 733 173 736
rect 210 733 220 736
rect 322 733 332 736
rect 450 733 492 736
rect 594 733 612 736
rect 682 733 692 736
rect 756 733 765 736
rect 786 733 796 736
rect 842 733 860 736
rect 916 733 933 736
rect 170 726 173 733
rect 930 726 933 733
rect 1050 733 1060 736
rect 1050 726 1053 733
rect 1338 726 1341 734
rect 1364 733 1389 736
rect 1426 733 1460 736
rect 1490 733 1524 736
rect 1570 726 1573 734
rect 1642 733 1660 736
rect 1850 733 1860 736
rect 2154 733 2172 736
rect 2194 733 2244 736
rect 2260 733 2309 736
rect 2386 733 2396 736
rect 2418 733 2468 736
rect 2484 733 2525 736
rect 2546 733 2572 736
rect 2594 733 2604 736
rect 2618 733 2660 736
rect 2940 733 2949 736
rect 2962 733 2980 736
rect 3010 733 3036 736
rect 3084 733 3101 736
rect 3114 733 3132 736
rect 3162 733 3180 736
rect 3250 733 3292 736
rect 3306 733 3316 736
rect 3332 733 3349 736
rect 3354 733 3412 736
rect 3346 726 3349 733
rect 66 723 100 726
rect 140 723 149 726
rect 170 723 221 726
rect 314 723 340 726
rect 444 723 477 726
rect 522 723 556 726
rect 586 723 604 726
rect 642 723 676 726
rect 700 723 733 726
rect 764 723 773 726
rect 794 723 804 726
rect 834 723 901 726
rect 930 723 941 726
rect 962 723 1028 726
rect 1042 723 1053 726
rect 1068 723 1133 726
rect 1300 723 1341 726
rect 1532 723 1573 726
rect 1612 723 1621 726
rect 1626 723 1652 726
rect 1676 723 1693 726
rect 1746 723 1780 726
rect 1850 723 1868 726
rect 2042 723 2052 726
rect 2196 723 2236 726
rect 2298 723 2308 726
rect 2346 723 2388 726
rect 2434 723 2460 726
rect 2498 723 2540 726
rect 2586 723 2612 726
rect 2722 723 2732 726
rect 2812 723 2829 726
rect 2916 723 2941 726
rect 3148 723 3173 726
rect 3178 723 3188 726
rect 3300 723 3308 726
rect 3346 723 3405 726
rect 348 713 381 716
rect 388 713 397 716
rect 412 713 421 716
rect 1042 715 1045 723
rect 1252 713 1269 716
rect 1364 713 1389 716
rect 1682 713 1716 716
rect 1922 713 1948 716
rect 1972 713 2005 716
rect 2060 713 2093 716
rect 1386 706 1389 713
rect 2098 706 2101 715
rect 2124 713 2157 716
rect 2620 713 2661 716
rect 3244 713 3285 716
rect 250 703 300 706
rect 370 703 404 706
rect 1162 703 1172 706
rect 1386 703 1405 706
rect 1706 703 1732 706
rect 1818 703 1828 706
rect 2066 703 2101 706
rect 378 693 381 703
rect 14 667 3490 673
rect 3226 653 3269 656
rect 682 633 732 636
rect 954 633 996 636
rect 1010 633 1052 636
rect 116 623 141 626
rect 156 623 197 626
rect 274 616 277 626
rect 308 623 325 626
rect 620 623 645 626
rect 740 623 757 626
rect 828 623 837 626
rect 892 623 917 626
rect 980 623 989 626
rect 1036 623 1045 626
rect 1228 623 1237 626
rect 1282 616 1285 636
rect 1362 633 1373 636
rect 1348 623 1357 626
rect 148 613 189 616
rect 236 613 277 616
rect 306 613 332 616
rect 364 613 373 616
rect 540 613 549 616
rect 556 613 573 616
rect 626 613 660 616
rect 772 613 805 616
rect 890 613 932 616
rect 1138 613 1164 616
rect 1202 613 1212 616
rect 1226 613 1245 616
rect 1250 613 1260 616
rect 1282 613 1332 616
rect 1370 615 1373 633
rect 1506 633 1532 636
rect 1450 616 1453 625
rect 1506 616 1509 633
rect 1626 626 1629 636
rect 1770 633 1788 636
rect 2346 633 2381 636
rect 2386 633 2396 636
rect 2418 633 2452 636
rect 1626 623 1636 626
rect 1660 623 1669 626
rect 1724 623 1741 626
rect 1772 623 1781 626
rect 1892 623 1901 626
rect 2068 623 2093 626
rect 2116 623 2125 626
rect 2324 623 2373 626
rect 2378 625 2381 633
rect 2418 623 2436 626
rect 2460 623 2493 626
rect 2508 623 2533 626
rect 3180 623 3205 626
rect 3300 623 3317 626
rect 1450 613 1461 616
rect 1468 613 1509 616
rect 1612 613 1629 616
rect 1674 613 1708 616
rect 1722 613 1757 616
rect 114 603 140 606
rect 228 603 285 606
rect 356 603 397 606
rect 402 603 428 606
rect 442 603 452 606
rect 490 603 532 606
rect 676 603 709 606
rect 746 603 764 606
rect 786 603 804 606
rect 842 603 868 606
rect 892 603 909 606
rect 1114 603 1124 606
rect 1194 603 1204 606
rect 1226 605 1229 613
rect 1276 603 1285 606
rect 1290 603 1324 606
rect 1402 603 1428 606
rect 1690 603 1700 606
rect 1754 605 1757 613
rect 1778 593 1781 615
rect 1802 613 1860 616
rect 1866 613 1884 616
rect 1948 613 1957 616
rect 1962 613 1988 616
rect 2108 613 2149 616
rect 2156 613 2189 616
rect 2266 613 2284 616
rect 2298 613 2316 616
rect 2466 613 2493 616
rect 2178 606 2181 613
rect 1906 603 1940 606
rect 1970 603 1980 606
rect 2004 603 2021 606
rect 2082 603 2100 606
rect 2114 603 2148 606
rect 2178 603 2204 606
rect 2490 605 2493 613
rect 2530 606 2533 623
rect 3202 616 3205 623
rect 2572 613 2581 616
rect 2764 613 2813 616
rect 2852 613 2916 616
rect 3004 613 3037 616
rect 3044 613 3061 616
rect 3106 606 3109 615
rect 3114 613 3164 616
rect 3202 613 3212 616
rect 3242 613 3284 616
rect 3340 613 3349 616
rect 3362 613 3380 616
rect 2530 603 2541 606
rect 2564 603 2628 606
rect 2644 603 2653 606
rect 2690 603 2708 606
rect 2746 603 2756 606
rect 2770 603 2780 606
rect 2876 603 2917 606
rect 2946 603 2996 606
rect 3026 603 3036 606
rect 3050 603 3084 606
rect 3106 603 3149 606
rect 3180 603 3189 606
rect 3194 603 3204 606
rect 3226 603 3276 606
rect 3346 603 3388 606
rect 2666 593 2700 596
rect 2738 593 2748 596
rect 2962 593 2988 596
rect 38 567 3466 573
rect 554 543 596 546
rect 124 533 133 536
rect 170 533 204 536
rect 220 533 229 536
rect 170 526 173 533
rect 66 523 100 526
rect 148 523 173 526
rect 178 523 196 526
rect 242 523 245 534
rect 268 533 301 536
rect 418 533 428 536
rect 442 533 452 536
rect 538 533 548 536
rect 282 523 324 526
rect 466 523 508 526
rect 514 523 532 526
rect 554 525 557 543
rect 628 533 669 536
rect 770 533 788 536
rect 804 533 837 536
rect 914 526 917 534
rect 962 533 972 536
rect 994 533 1036 536
rect 1052 533 1061 536
rect 1074 526 1077 556
rect 1082 536 1085 556
rect 1082 533 1092 536
rect 1106 533 1140 536
rect 1156 533 1173 536
rect 1186 533 1204 536
rect 1218 533 1228 536
rect 1266 533 1284 536
rect 1330 533 1348 536
rect 1362 533 1404 536
rect 1458 533 1468 536
rect 1484 533 1493 536
rect 1578 533 1620 536
rect 1682 533 1708 536
rect 1786 533 1804 536
rect 700 523 725 526
rect 762 523 780 526
rect 812 523 837 526
rect 906 523 917 526
rect 938 523 964 526
rect 1002 523 1028 526
rect 1074 523 1100 526
rect 1106 523 1132 526
rect 1202 523 1212 526
rect 1218 523 1221 533
rect 1842 526 1845 546
rect 3218 543 3229 546
rect 1226 523 1236 526
rect 1274 523 1292 526
rect 1306 523 1316 526
rect 1428 523 1445 526
rect 1450 523 1460 526
rect 1634 523 1652 526
rect 1724 523 1733 526
rect 1770 523 1796 526
rect 1828 523 1845 526
rect 1882 533 1924 536
rect 1940 533 1988 536
rect 2092 533 2148 536
rect 2178 533 2204 536
rect 2220 533 2245 536
rect 2282 533 2292 536
rect 2306 533 2348 536
rect 2364 533 2389 536
rect 2466 533 2492 536
rect 178 516 181 523
rect 162 513 181 516
rect 346 503 372 506
rect 714 503 748 506
rect 906 503 909 523
rect 1882 516 1885 533
rect 2514 526 2517 535
rect 2530 533 2580 536
rect 2682 533 2716 536
rect 2730 526 2733 535
rect 2826 533 2836 536
rect 2922 533 2948 536
rect 2972 533 2981 536
rect 3042 533 3068 536
rect 3106 533 3116 536
rect 3148 533 3157 536
rect 3170 533 3188 536
rect 3212 533 3221 536
rect 3226 526 3229 543
rect 3274 533 3300 536
rect 3324 533 3333 536
rect 3364 533 3389 536
rect 3394 526 3397 535
rect 3420 533 3437 536
rect 1962 523 1980 526
rect 2050 523 2076 526
rect 2100 523 2109 526
rect 2178 523 2196 526
rect 2228 523 2261 526
rect 2330 523 2340 526
rect 2372 523 2397 526
rect 2402 523 2412 526
rect 2426 523 2452 526
rect 2458 523 2517 526
rect 2524 523 2557 526
rect 2570 523 2588 526
rect 2724 523 2733 526
rect 2818 523 2876 526
rect 2916 523 2956 526
rect 2970 523 3004 526
rect 3058 523 3076 526
rect 3162 523 3196 526
rect 3226 523 3244 526
rect 3298 523 3308 526
rect 3378 523 3397 526
rect 1108 513 1117 516
rect 1364 513 1381 516
rect 1668 513 1677 516
rect 1764 513 1789 516
rect 1834 513 1852 516
rect 1876 513 1885 516
rect 2172 513 2189 516
rect 2420 513 2445 516
rect 2460 513 2493 516
rect 2612 513 2645 516
rect 2652 513 2661 516
rect 2892 513 2901 516
rect 2972 513 2989 516
rect 3092 513 3101 516
rect 3212 513 3229 516
rect 3260 513 3269 516
rect 3364 513 3381 516
rect 1498 503 1548 506
rect 1730 503 1756 506
rect 1850 503 1868 506
rect 14 467 3490 473
rect 146 423 165 426
rect 180 423 197 426
rect 324 423 349 426
rect 404 423 413 426
rect 428 423 461 426
rect 884 423 901 426
rect 932 423 941 426
rect 1052 423 1061 426
rect 1076 423 1125 426
rect 146 416 149 423
rect 132 413 149 416
rect 154 413 172 416
rect 186 413 228 416
rect 266 413 316 416
rect 356 413 389 416
rect 442 413 468 416
rect 578 413 596 416
rect 602 413 661 416
rect 692 413 740 416
rect 772 413 797 416
rect 818 413 828 416
rect 850 413 869 416
rect 876 413 885 416
rect 890 413 924 416
rect 1002 413 1044 416
rect 1068 413 1085 416
rect 1154 413 1172 416
rect 124 403 141 406
rect 146 403 164 406
rect 226 403 236 406
rect 252 403 277 406
rect 322 403 348 406
rect 514 403 565 406
rect 506 393 548 396
rect 658 395 661 413
rect 668 403 684 406
rect 764 403 773 406
rect 802 403 820 406
rect 844 403 861 406
rect 866 405 869 413
rect 906 403 916 406
rect 954 403 972 406
rect 994 403 1036 406
rect 1050 403 1060 406
rect 1122 403 1132 406
rect 1178 403 1181 425
rect 1516 423 1557 426
rect 1674 416 1677 425
rect 1778 416 1781 426
rect 1820 423 1853 426
rect 1956 423 1965 426
rect 2004 423 2029 426
rect 2324 423 2373 426
rect 2604 423 2613 426
rect 2026 416 2029 423
rect 1194 413 1236 416
rect 1276 413 1285 416
rect 1300 413 1309 416
rect 1364 413 1373 416
rect 1420 413 1429 416
rect 1476 413 1500 416
rect 1634 413 1668 416
rect 1674 413 1692 416
rect 1770 413 1781 416
rect 1794 413 1804 416
rect 1914 413 1940 416
rect 2026 413 2044 416
rect 2050 413 2060 416
rect 2140 413 2189 416
rect 2338 413 2380 416
rect 2420 413 2429 416
rect 2490 413 2508 416
rect 2514 413 2524 416
rect 2538 413 2572 416
rect 2650 413 2668 416
rect 2828 413 2845 416
rect 2980 413 3005 416
rect 3092 413 3101 416
rect 3140 413 3165 416
rect 3364 413 3389 416
rect 1194 403 1228 406
rect 1242 403 1260 406
rect 1356 403 1365 406
rect 1370 405 1373 413
rect 1538 403 1556 406
rect 1586 403 1596 406
rect 1620 403 1653 406
rect 1770 405 1773 413
rect 2842 406 2845 413
rect 1820 403 1837 406
rect 1884 403 1925 406
rect 1970 403 1988 406
rect 2026 403 2036 406
rect 2154 403 2204 406
rect 2220 403 2245 406
rect 2250 403 2276 406
rect 2362 403 2372 406
rect 2842 403 2860 406
rect 1298 393 1348 396
rect 38 367 3466 373
rect 2106 346 2109 356
rect 834 343 860 346
rect 1266 336 1269 346
rect 2106 343 2125 346
rect 82 333 100 336
rect 124 333 133 336
rect 178 333 204 336
rect 338 333 372 336
rect 426 333 444 336
rect 474 333 524 336
rect 540 333 573 336
rect 658 333 668 336
rect 698 333 756 336
rect 826 333 868 336
rect 954 333 988 336
rect 1002 333 1044 336
rect 1146 333 1172 336
rect 1210 333 1220 336
rect 1266 333 1276 336
rect 1290 333 1300 336
rect 1322 333 1396 336
rect 1482 333 1493 336
rect 1642 333 1652 336
rect 1698 333 1724 336
rect 1746 333 1772 336
rect 1818 333 1828 336
rect 1842 333 1876 336
rect 1900 333 1909 336
rect 1978 333 2028 336
rect 2058 333 2076 336
rect 426 326 429 333
rect 570 326 573 333
rect 226 323 252 326
rect 396 323 429 326
rect 468 323 501 326
rect 570 323 588 326
rect 652 323 676 326
rect 730 323 764 326
rect 770 323 780 326
rect 786 323 820 326
rect 876 323 885 326
rect 890 323 924 326
rect 1052 323 1069 326
rect 1146 316 1149 333
rect 1482 326 1485 333
rect 1698 326 1701 333
rect 2098 326 2101 335
rect 2106 333 2148 336
rect 2258 333 2268 336
rect 2404 333 2453 336
rect 2474 333 2484 336
rect 1196 323 1221 326
rect 1228 323 1261 326
rect 1324 323 1333 326
rect 1404 323 1413 326
rect 1428 323 1485 326
rect 1524 323 1533 326
rect 1554 323 1596 326
rect 1660 323 1701 326
rect 1754 323 1780 326
rect 1786 323 1836 326
rect 1842 323 1884 326
rect 1980 323 2005 326
rect 2036 323 2084 326
rect 2098 323 2125 326
rect 2130 323 2140 326
rect 2172 323 2221 326
rect 2250 323 2276 326
rect 2282 323 2332 326
rect 2346 323 2380 326
rect 2458 323 2485 326
rect 2492 323 2509 326
rect 2530 323 2556 326
rect 260 313 301 316
rect 308 313 317 316
rect 332 313 357 316
rect 596 313 629 316
rect 828 313 837 316
rect 1004 313 1045 316
rect 1116 313 1149 316
rect 1436 313 1477 316
rect 274 303 324 306
rect 1074 303 1108 306
rect 1474 303 1477 313
rect 1554 303 1557 323
rect 2530 316 2533 323
rect 1668 313 1685 316
rect 1844 313 1869 316
rect 1900 313 1941 316
rect 2044 313 2069 316
rect 2100 313 2133 316
rect 2284 313 2325 316
rect 2340 313 2373 316
rect 2476 313 2485 316
rect 2500 313 2533 316
rect 2610 313 2644 316
rect 2674 313 2716 316
rect 1866 303 1869 313
rect 1938 303 1941 313
rect 2722 306 2725 325
rect 2836 323 2861 326
rect 2956 323 2981 326
rect 3012 323 3037 326
rect 3076 323 3085 326
rect 3220 323 3245 326
rect 3364 323 3389 326
rect 2586 303 2596 306
rect 2626 303 2660 306
rect 2690 303 2725 306
rect 14 267 3490 273
rect 194 233 204 236
rect 362 233 404 236
rect 906 233 916 236
rect 938 233 988 236
rect 1130 233 1156 236
rect 1378 233 1420 236
rect 2442 233 2468 236
rect 2610 233 2645 236
rect 212 223 245 226
rect 370 223 388 226
rect 460 223 501 226
rect 554 223 573 226
rect 636 223 669 226
rect 764 223 773 226
rect 884 223 893 226
rect 924 223 933 226
rect 1338 223 1348 226
rect 1386 223 1404 226
rect 2188 223 2221 226
rect 2396 223 2405 226
rect 2426 223 2452 226
rect 2578 223 2636 226
rect 66 213 108 216
rect 140 213 165 216
rect 242 206 245 223
rect 570 216 573 223
rect 426 213 452 216
rect 458 213 525 216
rect 532 213 565 216
rect 570 213 580 216
rect 610 213 620 216
rect 132 203 173 206
rect 242 203 253 206
rect 276 203 293 206
rect 418 203 444 206
rect 522 205 525 213
rect 666 206 669 223
rect 756 213 789 216
rect 828 213 869 216
rect 1010 213 1028 216
rect 1108 213 1125 216
rect 1194 213 1204 216
rect 1236 213 1245 216
rect 1258 213 1276 216
rect 1308 213 1333 216
rect 1450 213 1460 216
rect 1498 213 1548 216
rect 786 206 789 213
rect 1586 206 1589 215
rect 1594 213 1652 216
rect 1658 213 1701 216
rect 1724 213 1765 216
rect 1786 213 1804 216
rect 1890 213 1924 216
rect 1956 213 2012 216
rect 2050 213 2092 216
rect 1698 206 1701 213
rect 2154 206 2157 216
rect 2162 213 2180 216
rect 2186 213 2228 216
rect 2260 213 2301 216
rect 2306 213 2316 216
rect 2348 213 2357 216
rect 2626 213 2629 223
rect 2642 215 2645 233
rect 3170 233 3189 236
rect 3170 216 3173 233
rect 2676 213 2701 216
rect 2770 213 2796 216
rect 2844 213 2893 216
rect 2930 213 2948 216
rect 3012 213 3053 216
rect 3132 213 3173 216
rect 3186 215 3189 233
rect 3220 213 3261 216
rect 3300 213 3325 216
rect 3412 213 3437 216
rect 2306 206 2309 213
rect 594 203 612 206
rect 666 203 677 206
rect 706 203 748 206
rect 786 203 804 206
rect 826 203 868 206
rect 1002 203 1036 206
rect 1058 203 1100 206
rect 1242 203 1284 206
rect 1442 203 1468 206
rect 1586 203 1629 206
rect 1698 203 1716 206
rect 1746 203 1772 206
rect 1954 203 2004 206
rect 2026 203 2077 206
rect 2090 203 2100 206
rect 2154 203 2172 206
rect 2202 203 2236 206
rect 2282 203 2309 206
rect 2340 203 2349 206
rect 2764 203 2781 206
rect 2866 203 2900 206
rect 2930 203 2940 206
rect 1738 193 1764 196
rect 2018 193 2028 196
rect 3050 195 3053 213
rect 3060 203 3093 206
rect 3226 203 3268 206
rect 3346 203 3380 206
rect 38 167 3466 173
rect 810 136 813 146
rect 1330 143 1356 146
rect 122 133 180 136
rect 234 133 244 136
rect 348 133 357 136
rect 426 133 436 136
rect 532 133 557 136
rect 562 133 572 136
rect 610 133 636 136
rect 610 126 613 133
rect 658 126 661 135
rect 684 133 717 136
rect 764 133 797 136
rect 810 133 820 136
rect 892 133 949 136
rect 986 133 1020 136
rect 1042 126 1045 135
rect 1050 133 1092 136
rect 1108 133 1157 136
rect 1162 126 1165 135
rect 1252 133 1285 136
rect 1316 133 1349 136
rect 1354 133 1364 136
rect 1436 133 1461 136
rect 1540 133 1549 136
rect 1562 133 1572 136
rect 1698 133 1748 136
rect 1820 133 1829 136
rect 1834 133 1844 136
rect 1858 133 1876 136
rect 1954 133 1972 136
rect 2010 133 2044 136
rect 1354 126 1357 133
rect 2058 126 2061 135
rect 2074 133 2124 136
rect 2258 133 2292 136
rect 2338 133 2357 136
rect 2402 133 2452 136
rect 2650 133 2676 136
rect 2698 133 2708 136
rect 2836 133 2861 136
rect 2338 126 2341 133
rect 2954 126 2957 134
rect 3010 126 3013 134
rect 3074 126 3077 134
rect 3090 133 3100 136
rect 3146 133 3180 136
rect 3204 133 3221 136
rect 3250 133 3260 136
rect 3314 126 3317 136
rect 3370 133 3412 136
rect 178 123 188 126
rect 226 123 236 126
rect 268 123 317 126
rect 420 123 437 126
rect 444 123 501 126
rect 546 123 613 126
rect 644 123 661 126
rect 802 123 828 126
rect 834 123 868 126
rect 906 123 948 126
rect 980 123 1013 126
rect 1018 123 1028 126
rect 1042 123 1077 126
rect 1122 123 1165 126
rect 1172 123 1181 126
rect 1194 123 1236 126
rect 1250 123 1300 126
rect 1314 123 1357 126
rect 1378 123 1420 126
rect 1450 123 1500 126
rect 1548 123 1557 126
rect 1580 123 1613 126
rect 1706 123 1740 126
rect 1828 123 1845 126
rect 1852 123 1877 126
rect 1890 123 1924 126
rect 1946 123 1980 126
rect 2052 123 2061 126
rect 2068 123 2117 126
rect 2132 123 2149 126
rect 196 113 229 116
rect 684 113 733 116
rect 836 113 861 116
rect 1252 113 1261 116
rect 1316 113 1325 116
rect 1508 113 1517 116
rect 1586 113 1620 116
rect 1644 113 1661 116
rect 1692 113 1733 116
rect 1940 113 1965 116
rect 1996 113 2037 116
rect 2140 113 2149 116
rect 2146 106 2149 113
rect 2162 106 2165 125
rect 2316 123 2341 126
rect 2346 123 2364 126
rect 2426 123 2444 126
rect 2186 113 2228 116
rect 2252 113 2277 116
rect 2556 113 2565 116
rect 2618 106 2621 125
rect 2642 123 2684 126
rect 2690 123 2716 126
rect 2930 123 2957 126
rect 2986 123 3013 126
rect 3020 123 3077 126
rect 3084 123 3101 126
rect 3226 123 3244 126
rect 3250 123 3317 126
rect 3346 123 3364 126
rect 3378 123 3429 126
rect 3226 116 3229 123
rect 3204 113 3229 116
rect 3346 115 3349 123
rect 1650 103 1684 106
rect 2146 103 2165 106
rect 2186 103 2244 106
rect 2530 103 2572 106
rect 2586 103 2621 106
rect 14 67 3490 73
rect 38 37 3466 57
rect 14 13 3490 33
<< metal2 >>
rect 14 13 34 3327
rect 506 3306 509 3326
rect 38 37 58 3303
rect 434 3223 461 3226
rect 74 3036 77 3216
rect 82 3193 85 3206
rect 146 3166 149 3206
rect 194 3176 197 3216
rect 226 3193 229 3216
rect 194 3173 245 3176
rect 258 3173 261 3206
rect 306 3193 309 3216
rect 70 3033 77 3036
rect 90 3163 149 3166
rect 70 2966 73 3033
rect 90 2983 93 3163
rect 138 3123 141 3136
rect 210 3106 213 3126
rect 202 3103 213 3106
rect 218 3106 221 3136
rect 242 3133 245 3173
rect 266 3133 277 3136
rect 314 3133 317 3176
rect 226 3113 229 3126
rect 234 3123 245 3126
rect 234 3106 237 3123
rect 218 3103 237 3106
rect 242 3103 245 3116
rect 202 3056 205 3103
rect 202 3053 213 3056
rect 138 2993 141 3016
rect 154 2976 157 3036
rect 210 3033 213 3053
rect 218 3026 221 3103
rect 258 3033 261 3126
rect 362 3123 365 3136
rect 290 3093 293 3116
rect 386 3046 389 3206
rect 394 3176 397 3216
rect 410 3193 413 3206
rect 394 3173 405 3176
rect 402 3066 405 3173
rect 418 3126 421 3146
rect 370 3043 389 3046
rect 394 3063 405 3066
rect 414 3123 421 3126
rect 210 3023 221 3026
rect 146 2973 157 2976
rect 70 2963 77 2966
rect 74 2943 77 2963
rect 82 2836 85 2966
rect 122 2943 125 2956
rect 146 2943 149 2973
rect 202 2953 205 3016
rect 210 3003 213 3023
rect 258 3013 261 3026
rect 322 3013 325 3026
rect 234 2993 237 3006
rect 74 2833 85 2836
rect 74 2756 77 2833
rect 114 2813 117 2936
rect 146 2933 157 2936
rect 122 2923 141 2926
rect 138 2913 141 2923
rect 154 2856 157 2933
rect 162 2913 165 2926
rect 194 2876 197 2936
rect 210 2933 213 2986
rect 274 2983 277 3006
rect 258 2923 261 2946
rect 194 2873 229 2876
rect 154 2853 161 2856
rect 90 2776 93 2806
rect 158 2776 161 2853
rect 90 2773 125 2776
rect 74 2753 85 2756
rect 82 2646 85 2753
rect 122 2733 125 2773
rect 154 2773 161 2776
rect 154 2723 157 2773
rect 170 2756 173 2816
rect 226 2813 229 2873
rect 266 2846 269 2866
rect 266 2843 273 2846
rect 202 2773 205 2806
rect 270 2776 273 2843
rect 290 2826 293 2926
rect 338 2846 341 2956
rect 346 2916 349 2926
rect 354 2923 357 2936
rect 362 2923 365 2936
rect 370 2933 373 3043
rect 394 3026 397 3063
rect 386 3023 397 3026
rect 386 2956 389 3023
rect 402 2993 405 3046
rect 414 3036 417 3123
rect 426 3076 429 3216
rect 458 3213 461 3223
rect 450 3193 453 3206
rect 482 3163 485 3216
rect 490 3203 493 3226
rect 498 3203 501 3306
rect 506 3303 513 3306
rect 510 3236 513 3303
rect 506 3233 513 3236
rect 506 3156 509 3233
rect 522 3176 525 3306
rect 562 3266 565 3340
rect 578 3323 581 3340
rect 522 3173 529 3176
rect 434 3133 437 3156
rect 474 3153 509 3156
rect 450 3133 461 3136
rect 442 3106 445 3126
rect 474 3116 477 3153
rect 482 3143 501 3146
rect 482 3133 485 3143
rect 466 3113 477 3116
rect 442 3103 453 3106
rect 426 3073 437 3076
rect 414 3033 421 3036
rect 386 2953 405 2956
rect 394 2933 397 2946
rect 370 2916 373 2926
rect 402 2916 405 2953
rect 346 2913 373 2916
rect 394 2913 405 2916
rect 338 2843 349 2846
rect 290 2823 297 2826
rect 166 2753 173 2756
rect 166 2686 169 2753
rect 242 2733 245 2776
rect 266 2773 273 2776
rect 166 2683 173 2686
rect 74 2643 85 2646
rect 74 2626 77 2643
rect 170 2626 173 2683
rect 74 2623 109 2626
rect 74 2606 77 2623
rect 70 2603 77 2606
rect 70 2506 73 2603
rect 82 2513 85 2616
rect 106 2613 109 2623
rect 146 2623 173 2626
rect 98 2593 101 2606
rect 114 2603 117 2616
rect 146 2613 149 2623
rect 122 2546 125 2606
rect 130 2593 133 2606
rect 154 2596 157 2616
rect 170 2603 173 2616
rect 178 2603 181 2616
rect 202 2613 205 2726
rect 266 2686 269 2773
rect 250 2683 269 2686
rect 154 2593 181 2596
rect 186 2593 189 2606
rect 122 2543 133 2546
rect 70 2503 77 2506
rect 74 2376 77 2503
rect 98 2466 101 2536
rect 130 2496 133 2543
rect 90 2463 101 2466
rect 122 2493 133 2496
rect 74 2373 85 2376
rect 90 2373 93 2463
rect 122 2426 125 2493
rect 146 2456 149 2526
rect 178 2523 181 2593
rect 146 2453 165 2456
rect 122 2423 129 2426
rect 74 2266 77 2366
rect 82 2356 85 2373
rect 114 2366 117 2416
rect 126 2366 129 2423
rect 106 2363 117 2366
rect 122 2363 129 2366
rect 82 2353 93 2356
rect 70 2263 77 2266
rect 70 2026 73 2263
rect 90 2256 93 2353
rect 82 2253 93 2256
rect 82 2216 85 2253
rect 106 2216 109 2363
rect 82 2213 93 2216
rect 106 2213 117 2216
rect 82 2193 85 2206
rect 90 2183 93 2213
rect 114 2203 117 2213
rect 122 2156 125 2363
rect 138 2333 141 2376
rect 162 2346 165 2453
rect 178 2413 181 2516
rect 210 2456 213 2536
rect 234 2486 237 2616
rect 250 2536 253 2683
rect 258 2603 261 2616
rect 282 2613 285 2816
rect 294 2776 297 2823
rect 290 2773 297 2776
rect 314 2773 317 2806
rect 346 2796 349 2843
rect 394 2836 397 2913
rect 394 2833 405 2836
rect 362 2813 365 2826
rect 338 2793 349 2796
rect 290 2723 293 2773
rect 330 2706 333 2726
rect 322 2703 333 2706
rect 322 2636 325 2703
rect 322 2633 333 2636
rect 250 2533 257 2536
rect 202 2453 213 2456
rect 230 2483 237 2486
rect 202 2373 205 2453
rect 230 2406 233 2483
rect 242 2433 245 2526
rect 254 2466 257 2533
rect 250 2463 257 2466
rect 230 2403 237 2406
rect 162 2343 173 2346
rect 170 2296 173 2343
rect 162 2293 173 2296
rect 82 2153 125 2156
rect 82 2026 85 2153
rect 106 2143 125 2146
rect 90 2083 93 2126
rect 98 2113 101 2136
rect 106 2123 109 2143
rect 106 2026 109 2046
rect 70 2023 77 2026
rect 82 2023 93 2026
rect 66 1983 69 2006
rect 66 1473 69 1836
rect 66 1323 69 1406
rect 74 1306 77 2023
rect 82 1933 85 2016
rect 90 1916 93 2023
rect 98 2023 109 2026
rect 98 1923 101 2023
rect 114 2016 117 2136
rect 122 2133 125 2143
rect 106 2013 117 2016
rect 122 2013 125 2036
rect 114 2003 125 2006
rect 106 1916 109 1996
rect 86 1913 93 1916
rect 98 1913 109 1916
rect 86 1846 89 1913
rect 86 1843 93 1846
rect 82 1603 85 1826
rect 90 1673 93 1843
rect 90 1613 93 1626
rect 82 1503 85 1596
rect 82 1483 85 1496
rect 82 1393 85 1436
rect 90 1403 93 1606
rect 82 1333 85 1346
rect 70 1303 77 1306
rect 70 1146 73 1303
rect 70 1143 77 1146
rect 66 743 69 1126
rect 66 723 69 736
rect 66 316 69 626
rect 74 383 77 1143
rect 82 1096 85 1296
rect 90 1203 93 1386
rect 98 1166 101 1913
rect 122 1856 125 1926
rect 106 1853 125 1856
rect 130 1853 133 2226
rect 162 2216 165 2293
rect 186 2226 189 2326
rect 234 2323 237 2403
rect 242 2343 245 2416
rect 250 2306 253 2463
rect 290 2413 293 2616
rect 306 2533 309 2606
rect 314 2596 317 2616
rect 322 2603 325 2616
rect 330 2613 333 2633
rect 338 2603 341 2793
rect 362 2696 365 2776
rect 354 2693 365 2696
rect 354 2613 357 2693
rect 394 2686 397 2816
rect 402 2793 405 2833
rect 410 2816 413 3016
rect 418 2963 421 3033
rect 426 3003 429 3026
rect 434 3013 437 3073
rect 450 3036 453 3103
rect 466 3056 469 3113
rect 466 3053 477 3056
rect 450 3033 461 3036
rect 442 3023 453 3026
rect 418 2913 421 2936
rect 410 2813 421 2816
rect 410 2723 413 2806
rect 418 2773 421 2813
rect 426 2746 429 2786
rect 434 2766 437 2986
rect 450 2973 453 3006
rect 458 2956 461 3033
rect 466 3013 469 3026
rect 474 2966 477 3053
rect 482 3026 485 3126
rect 490 3113 493 3136
rect 498 3123 501 3143
rect 506 3106 509 3136
rect 502 3103 509 3106
rect 482 3023 493 3026
rect 490 3013 493 3023
rect 502 2986 505 3103
rect 502 2983 509 2986
rect 474 2963 501 2966
rect 458 2953 477 2956
rect 442 2833 461 2836
rect 442 2813 445 2833
rect 450 2803 453 2826
rect 458 2816 461 2833
rect 466 2816 469 2826
rect 458 2813 469 2816
rect 450 2773 453 2796
rect 466 2783 469 2806
rect 474 2793 477 2953
rect 482 2923 485 2946
rect 434 2763 477 2766
rect 426 2743 433 2746
rect 430 2686 433 2743
rect 474 2733 477 2763
rect 490 2743 493 2826
rect 498 2806 501 2963
rect 506 2903 509 2983
rect 514 2823 517 3166
rect 526 3106 529 3173
rect 538 3133 541 3266
rect 546 3263 565 3266
rect 602 3263 605 3340
rect 618 3303 621 3340
rect 634 3296 637 3340
rect 630 3293 637 3296
rect 546 3213 549 3263
rect 630 3236 633 3293
rect 562 3223 565 3236
rect 618 3233 633 3236
rect 642 3283 661 3286
rect 570 3136 573 3206
rect 578 3143 581 3216
rect 594 3213 597 3226
rect 594 3193 597 3206
rect 546 3123 549 3136
rect 554 3106 557 3126
rect 526 3103 541 3106
rect 546 3103 557 3106
rect 522 3073 525 3096
rect 522 2993 525 3006
rect 522 2916 525 2986
rect 530 2933 533 3016
rect 538 2916 541 3103
rect 546 3013 549 3026
rect 546 2963 549 3006
rect 554 2996 557 3076
rect 562 3003 565 3136
rect 570 3133 581 3136
rect 570 3023 573 3126
rect 578 3026 581 3133
rect 602 3126 605 3136
rect 586 3053 589 3126
rect 594 3123 605 3126
rect 594 3113 597 3123
rect 610 3073 613 3126
rect 578 3023 613 3026
rect 578 3003 581 3023
rect 554 2993 573 2996
rect 562 2933 565 2986
rect 570 2976 573 2993
rect 570 2973 577 2976
rect 522 2913 529 2916
rect 526 2836 529 2913
rect 522 2833 529 2836
rect 538 2913 549 2916
rect 498 2803 509 2806
rect 442 2696 445 2726
rect 506 2696 509 2803
rect 522 2783 525 2833
rect 538 2816 541 2913
rect 554 2843 557 2926
rect 574 2916 577 2973
rect 586 2953 589 3016
rect 602 2973 605 3006
rect 610 3003 613 3023
rect 618 2946 621 3233
rect 642 3226 645 3283
rect 634 3223 645 3226
rect 642 3213 653 3216
rect 658 3213 661 3283
rect 674 3213 677 3256
rect 682 3213 685 3266
rect 698 3223 701 3340
rect 626 3043 629 3136
rect 634 3113 637 3206
rect 642 3183 645 3206
rect 650 3106 653 3213
rect 682 3193 685 3206
rect 642 3103 653 3106
rect 658 3103 661 3126
rect 642 3036 645 3103
rect 626 3023 629 3036
rect 634 3033 645 3036
rect 634 3016 637 3033
rect 658 3023 661 3096
rect 630 3013 637 3016
rect 630 2956 633 3013
rect 642 2983 645 3016
rect 666 3013 669 3136
rect 674 3083 677 3126
rect 682 3123 685 3156
rect 690 3133 693 3206
rect 698 3203 701 3216
rect 714 3213 717 3296
rect 706 3133 709 3206
rect 714 3133 717 3186
rect 674 3006 677 3056
rect 698 3033 701 3126
rect 714 3113 717 3126
rect 722 3123 725 3306
rect 730 3246 733 3266
rect 730 3243 737 3246
rect 734 3126 737 3243
rect 730 3123 737 3126
rect 730 3106 733 3123
rect 722 3103 733 3106
rect 706 3026 709 3056
rect 722 3046 725 3103
rect 586 2933 589 2946
rect 610 2943 621 2946
rect 626 2953 633 2956
rect 610 2916 613 2943
rect 618 2923 621 2936
rect 626 2916 629 2953
rect 650 2933 653 3006
rect 658 2993 661 3006
rect 666 3003 677 3006
rect 698 3023 709 3026
rect 714 3043 725 3046
rect 666 2986 669 3003
rect 658 2983 669 2986
rect 574 2913 581 2916
rect 530 2813 541 2816
rect 530 2796 533 2813
rect 530 2793 541 2796
rect 538 2756 541 2793
rect 546 2776 549 2816
rect 546 2773 557 2776
rect 522 2723 525 2756
rect 538 2753 549 2756
rect 442 2693 453 2696
rect 362 2683 397 2686
rect 426 2683 433 2686
rect 314 2593 325 2596
rect 314 2576 317 2593
rect 314 2573 325 2576
rect 322 2526 325 2573
rect 314 2523 325 2526
rect 314 2436 317 2523
rect 298 2433 317 2436
rect 298 2356 301 2433
rect 314 2393 317 2406
rect 274 2353 301 2356
rect 242 2303 253 2306
rect 242 2246 245 2303
rect 242 2243 253 2246
rect 162 2213 173 2216
rect 138 2193 141 2206
rect 170 2203 173 2213
rect 138 2116 141 2136
rect 138 2113 145 2116
rect 142 2036 145 2113
rect 138 2033 145 2036
rect 106 1283 109 1853
rect 114 1793 117 1816
rect 114 1603 117 1736
rect 122 1596 125 1846
rect 130 1813 133 1836
rect 130 1733 133 1806
rect 130 1713 133 1726
rect 138 1713 141 2033
rect 146 1843 149 2016
rect 154 1993 157 2086
rect 170 2026 173 2126
rect 178 2106 181 2226
rect 186 2223 237 2226
rect 234 2216 237 2223
rect 186 2193 189 2206
rect 226 2196 229 2216
rect 234 2213 245 2216
rect 242 2203 245 2213
rect 250 2196 253 2243
rect 258 2213 261 2336
rect 274 2303 277 2353
rect 290 2333 293 2346
rect 306 2323 309 2336
rect 322 2323 325 2346
rect 338 2333 341 2436
rect 346 2426 349 2576
rect 354 2533 357 2606
rect 362 2523 365 2683
rect 378 2603 381 2616
rect 370 2533 373 2556
rect 418 2546 421 2626
rect 426 2613 429 2683
rect 450 2546 453 2693
rect 498 2693 509 2696
rect 466 2573 469 2606
rect 490 2596 493 2616
rect 498 2613 501 2693
rect 546 2686 549 2753
rect 538 2683 549 2686
rect 514 2603 517 2626
rect 530 2613 533 2626
rect 538 2613 541 2683
rect 562 2636 565 2906
rect 578 2846 581 2913
rect 570 2843 581 2846
rect 602 2913 613 2916
rect 602 2846 605 2913
rect 602 2843 613 2846
rect 570 2816 573 2843
rect 578 2823 605 2826
rect 570 2813 589 2816
rect 570 2753 573 2806
rect 586 2793 589 2813
rect 594 2803 597 2816
rect 602 2813 605 2823
rect 610 2803 613 2843
rect 618 2833 621 2916
rect 626 2913 633 2916
rect 630 2836 633 2913
rect 642 2903 645 2926
rect 658 2863 661 2983
rect 698 2976 701 3023
rect 714 3003 717 3043
rect 666 2973 717 2976
rect 666 2923 669 2973
rect 674 2963 709 2966
rect 674 2933 677 2963
rect 682 2923 685 2936
rect 698 2933 701 2956
rect 706 2936 709 2963
rect 714 2943 717 2973
rect 722 2943 725 3016
rect 730 3003 733 3026
rect 738 2946 741 3016
rect 746 3003 749 3340
rect 778 3216 781 3340
rect 882 3246 885 3340
rect 914 3323 917 3340
rect 954 3326 957 3340
rect 1034 3326 1037 3340
rect 946 3323 957 3326
rect 962 3323 973 3326
rect 878 3243 885 3246
rect 762 3213 781 3216
rect 786 3213 789 3236
rect 754 3183 757 3206
rect 754 3093 757 3126
rect 762 3023 765 3213
rect 770 3166 773 3206
rect 770 3163 781 3166
rect 770 3133 773 3146
rect 778 3143 781 3163
rect 778 3073 781 3126
rect 754 2963 757 3006
rect 770 2953 773 3016
rect 778 2983 781 2996
rect 786 2946 789 3206
rect 794 3053 797 3166
rect 802 3106 805 3226
rect 810 3133 813 3216
rect 818 3213 821 3226
rect 850 3223 861 3226
rect 850 3206 853 3216
rect 858 3213 861 3223
rect 818 3126 821 3206
rect 834 3126 837 3206
rect 842 3203 853 3206
rect 842 3183 845 3203
rect 850 3173 853 3196
rect 818 3123 829 3126
rect 834 3123 845 3126
rect 866 3116 869 3206
rect 878 3186 881 3243
rect 890 3233 901 3236
rect 890 3213 893 3233
rect 898 3203 901 3226
rect 906 3213 909 3266
rect 946 3256 949 3323
rect 914 3253 949 3256
rect 858 3113 869 3116
rect 874 3183 881 3186
rect 802 3103 813 3106
rect 810 3046 813 3103
rect 738 2943 789 2946
rect 794 3043 813 3046
rect 738 2936 741 2943
rect 706 2933 741 2936
rect 690 2893 693 2926
rect 706 2923 709 2933
rect 746 2913 749 2936
rect 626 2833 633 2836
rect 618 2813 621 2826
rect 602 2743 605 2776
rect 610 2716 613 2736
rect 618 2723 621 2746
rect 602 2713 613 2716
rect 602 2666 605 2713
rect 602 2663 613 2666
rect 554 2633 565 2636
rect 530 2603 541 2606
rect 490 2593 533 2596
rect 538 2593 541 2603
rect 418 2543 429 2546
rect 410 2506 413 2526
rect 402 2503 413 2506
rect 346 2423 357 2426
rect 290 2246 293 2316
rect 274 2243 293 2246
rect 226 2193 253 2196
rect 186 2123 189 2166
rect 194 2133 197 2146
rect 178 2103 185 2106
rect 182 2026 185 2103
rect 162 2023 173 2026
rect 178 2023 185 2026
rect 146 1813 149 1826
rect 154 1806 157 1986
rect 162 1936 165 2023
rect 170 2003 173 2016
rect 162 1933 173 1936
rect 162 1866 165 1926
rect 170 1873 173 1933
rect 162 1863 173 1866
rect 146 1803 157 1806
rect 130 1613 133 1646
rect 138 1613 141 1686
rect 146 1613 149 1786
rect 114 1593 125 1596
rect 130 1593 133 1606
rect 114 1513 117 1593
rect 122 1583 133 1586
rect 122 1536 125 1576
rect 130 1543 133 1583
rect 138 1536 141 1606
rect 154 1603 157 1726
rect 122 1533 133 1536
rect 138 1533 149 1536
rect 130 1513 133 1526
rect 114 1436 117 1506
rect 114 1433 125 1436
rect 114 1413 117 1426
rect 90 1163 101 1166
rect 90 1123 93 1163
rect 106 1156 109 1226
rect 114 1163 117 1406
rect 98 1153 109 1156
rect 98 1133 101 1153
rect 106 1113 109 1126
rect 114 1096 117 1136
rect 122 1133 125 1433
rect 130 1126 133 1476
rect 138 1433 141 1526
rect 146 1423 149 1533
rect 138 1323 141 1396
rect 146 1383 149 1406
rect 154 1376 157 1536
rect 162 1396 165 1856
rect 170 1783 173 1863
rect 170 1633 173 1736
rect 170 1613 173 1626
rect 170 1423 173 1516
rect 162 1393 169 1396
rect 146 1373 157 1376
rect 146 1233 149 1373
rect 154 1323 157 1346
rect 166 1306 169 1393
rect 162 1303 169 1306
rect 162 1236 165 1303
rect 162 1233 173 1236
rect 138 1213 141 1226
rect 138 1143 141 1206
rect 154 1203 157 1216
rect 170 1203 173 1233
rect 122 1123 133 1126
rect 82 1093 93 1096
rect 90 1026 93 1093
rect 106 1093 117 1096
rect 106 1036 109 1093
rect 106 1033 117 1036
rect 86 1023 93 1026
rect 86 946 89 1023
rect 114 1013 117 1033
rect 98 1003 117 1006
rect 86 943 93 946
rect 98 943 101 956
rect 82 333 85 936
rect 90 926 93 943
rect 90 923 97 926
rect 94 826 97 923
rect 90 823 97 826
rect 90 586 93 823
rect 98 723 101 806
rect 106 783 109 1003
rect 114 953 117 996
rect 122 976 125 1106
rect 130 1096 133 1123
rect 138 1113 141 1136
rect 130 1093 137 1096
rect 134 996 137 1093
rect 146 1003 149 1166
rect 162 1133 173 1136
rect 134 993 149 996
rect 122 973 129 976
rect 114 933 117 946
rect 114 843 117 926
rect 126 846 129 973
rect 122 843 129 846
rect 114 823 117 836
rect 114 803 117 816
rect 122 806 125 843
rect 138 826 141 936
rect 130 823 141 826
rect 130 813 133 823
rect 146 806 149 993
rect 122 803 133 806
rect 98 603 101 636
rect 106 623 109 746
rect 114 733 117 756
rect 114 723 125 726
rect 130 716 133 803
rect 142 803 149 806
rect 142 746 145 803
rect 142 743 149 746
rect 122 713 133 716
rect 122 616 125 713
rect 146 636 149 743
rect 154 646 157 1026
rect 162 1013 165 1133
rect 170 1113 173 1126
rect 162 713 165 1006
rect 170 916 173 1016
rect 178 933 181 2023
rect 186 1923 189 2006
rect 194 1996 197 2116
rect 202 2113 205 2126
rect 210 2043 213 2116
rect 226 2096 229 2136
rect 218 2093 229 2096
rect 202 2023 213 2026
rect 202 2003 205 2023
rect 218 2013 221 2093
rect 234 2083 237 2156
rect 250 2123 253 2193
rect 258 2163 261 2206
rect 266 2146 269 2226
rect 262 2143 269 2146
rect 226 2003 229 2046
rect 234 2013 237 2036
rect 250 2013 253 2116
rect 262 2086 265 2143
rect 258 2083 265 2086
rect 194 1993 221 1996
rect 218 1986 221 1993
rect 242 1986 245 2006
rect 218 1983 229 1986
rect 186 1903 189 1916
rect 194 1886 197 1936
rect 186 1883 197 1886
rect 186 1843 189 1883
rect 202 1876 205 1936
rect 210 1923 213 1946
rect 194 1873 205 1876
rect 186 1793 189 1806
rect 186 1613 189 1786
rect 194 1733 197 1873
rect 202 1723 205 1756
rect 186 1216 189 1606
rect 194 1383 197 1716
rect 210 1703 213 1836
rect 218 1813 221 1966
rect 226 1923 229 1983
rect 238 1983 245 1986
rect 238 1926 241 1983
rect 234 1923 241 1926
rect 250 1923 253 2006
rect 234 1833 237 1923
rect 258 1916 261 2083
rect 266 1943 269 2076
rect 274 1963 277 2243
rect 290 2233 333 2236
rect 290 2213 293 2233
rect 306 2196 309 2216
rect 322 2213 325 2226
rect 282 2193 309 2196
rect 282 2123 285 2193
rect 290 2076 293 2136
rect 322 2133 325 2146
rect 298 2093 301 2126
rect 282 2073 293 2076
rect 282 2003 285 2073
rect 290 1993 293 2046
rect 298 2013 309 2016
rect 266 1933 277 1936
rect 242 1913 261 1916
rect 218 1683 221 1746
rect 226 1663 229 1826
rect 234 1793 237 1826
rect 234 1743 237 1756
rect 202 1613 205 1626
rect 210 1606 213 1656
rect 218 1613 221 1636
rect 226 1606 229 1646
rect 202 1603 213 1606
rect 218 1603 229 1606
rect 202 1443 205 1603
rect 194 1223 197 1326
rect 202 1303 205 1426
rect 210 1413 213 1536
rect 218 1533 221 1603
rect 234 1596 237 1726
rect 242 1716 245 1913
rect 250 1823 253 1906
rect 250 1733 253 1816
rect 258 1796 261 1906
rect 266 1903 269 1926
rect 274 1833 277 1916
rect 282 1863 285 1926
rect 266 1803 269 1816
rect 274 1803 277 1816
rect 258 1793 265 1796
rect 242 1713 253 1716
rect 250 1646 253 1713
rect 262 1676 265 1793
rect 274 1713 277 1786
rect 262 1673 269 1676
rect 226 1593 237 1596
rect 242 1643 253 1646
rect 218 1483 221 1526
rect 226 1466 229 1593
rect 242 1586 245 1643
rect 250 1603 253 1626
rect 234 1583 245 1586
rect 234 1533 237 1583
rect 258 1576 261 1616
rect 266 1613 269 1673
rect 254 1573 261 1576
rect 222 1463 229 1466
rect 234 1463 237 1516
rect 210 1393 213 1406
rect 222 1396 225 1463
rect 242 1453 245 1536
rect 254 1466 257 1573
rect 254 1463 261 1466
rect 258 1443 261 1463
rect 234 1423 261 1426
rect 234 1413 245 1416
rect 258 1413 261 1423
rect 266 1413 269 1606
rect 274 1413 277 1666
rect 282 1613 285 1796
rect 290 1743 293 1976
rect 298 1913 301 1936
rect 306 1903 309 1916
rect 298 1846 301 1866
rect 298 1843 305 1846
rect 302 1766 305 1843
rect 298 1763 305 1766
rect 290 1693 293 1736
rect 290 1616 293 1656
rect 298 1643 301 1763
rect 314 1746 317 2126
rect 322 1773 325 2016
rect 330 2013 333 2233
rect 338 2203 341 2316
rect 346 2186 349 2416
rect 354 2343 357 2423
rect 362 2403 365 2416
rect 378 2366 381 2476
rect 402 2456 405 2503
rect 402 2453 413 2456
rect 386 2416 389 2436
rect 386 2413 397 2416
rect 410 2413 413 2453
rect 426 2433 429 2543
rect 434 2533 437 2546
rect 442 2543 453 2546
rect 442 2523 445 2543
rect 506 2533 509 2556
rect 522 2533 525 2546
rect 498 2523 509 2526
rect 370 2363 381 2366
rect 354 2323 357 2336
rect 370 2316 373 2363
rect 394 2346 397 2413
rect 410 2386 413 2406
rect 426 2393 429 2406
rect 410 2383 421 2386
rect 342 2183 349 2186
rect 354 2313 373 2316
rect 386 2343 397 2346
rect 342 2116 345 2183
rect 354 2123 357 2313
rect 342 2113 349 2116
rect 338 2003 341 2046
rect 330 1803 333 1986
rect 306 1743 317 1746
rect 306 1726 309 1743
rect 314 1733 325 1736
rect 306 1723 317 1726
rect 306 1633 309 1716
rect 290 1613 301 1616
rect 306 1613 309 1626
rect 282 1503 285 1526
rect 218 1393 225 1396
rect 210 1226 213 1336
rect 218 1233 221 1393
rect 226 1293 229 1386
rect 242 1336 245 1413
rect 250 1393 253 1406
rect 242 1333 249 1336
rect 234 1253 237 1326
rect 186 1213 197 1216
rect 186 1163 189 1206
rect 186 1113 189 1126
rect 170 913 177 916
rect 174 836 177 913
rect 170 833 177 836
rect 170 803 173 833
rect 178 703 181 816
rect 186 803 189 1106
rect 194 933 197 1213
rect 202 1013 205 1226
rect 210 1223 217 1226
rect 214 1156 217 1223
rect 214 1153 221 1156
rect 210 1003 213 1136
rect 210 936 213 956
rect 206 933 213 936
rect 206 866 209 933
rect 206 863 213 866
rect 210 846 213 863
rect 218 853 221 1153
rect 226 936 229 1236
rect 234 953 237 1216
rect 246 1146 249 1333
rect 258 1166 261 1406
rect 266 1173 269 1406
rect 282 1396 285 1496
rect 278 1393 285 1396
rect 278 1336 281 1393
rect 274 1333 281 1336
rect 290 1333 293 1606
rect 306 1583 309 1606
rect 314 1593 317 1723
rect 322 1713 325 1726
rect 322 1586 325 1676
rect 314 1583 325 1586
rect 298 1513 301 1546
rect 306 1506 309 1576
rect 314 1513 317 1583
rect 330 1573 333 1796
rect 338 1783 341 1926
rect 322 1513 325 1566
rect 330 1533 333 1546
rect 306 1503 333 1506
rect 298 1403 301 1466
rect 274 1243 277 1333
rect 258 1163 269 1166
rect 242 1143 249 1146
rect 242 1103 245 1143
rect 250 1123 261 1126
rect 266 1096 269 1163
rect 274 1113 277 1236
rect 250 1093 269 1096
rect 250 1026 253 1093
rect 242 1023 253 1026
rect 226 933 237 936
rect 234 863 237 933
rect 210 843 237 846
rect 154 643 181 646
rect 146 633 169 636
rect 138 623 157 626
rect 90 583 97 586
rect 94 446 97 583
rect 90 443 97 446
rect 90 396 93 443
rect 98 413 101 426
rect 106 413 109 616
rect 122 613 129 616
rect 114 523 117 606
rect 126 566 129 613
rect 122 563 129 566
rect 122 506 125 563
rect 130 543 149 546
rect 130 533 133 543
rect 118 503 125 506
rect 118 436 121 503
rect 118 433 125 436
rect 90 393 97 396
rect 94 326 97 393
rect 106 336 109 406
rect 114 366 117 416
rect 122 396 125 433
rect 130 403 133 526
rect 138 456 141 536
rect 146 523 149 543
rect 154 493 157 623
rect 166 536 169 633
rect 166 533 173 536
rect 138 453 149 456
rect 138 403 141 416
rect 146 403 149 453
rect 162 423 165 516
rect 170 496 173 533
rect 178 513 181 643
rect 186 613 189 726
rect 194 633 197 826
rect 202 813 205 836
rect 226 826 229 836
rect 218 823 229 826
rect 194 596 197 626
rect 202 613 205 806
rect 218 793 221 823
rect 226 773 229 806
rect 210 723 213 736
rect 218 716 221 726
rect 226 723 229 746
rect 210 703 213 716
rect 218 713 225 716
rect 222 636 225 713
rect 222 633 229 636
rect 210 603 213 616
rect 218 596 221 616
rect 194 593 221 596
rect 170 493 177 496
rect 174 436 177 493
rect 170 433 177 436
rect 202 436 205 556
rect 226 533 229 633
rect 210 523 221 526
rect 226 513 229 526
rect 234 506 237 843
rect 242 733 245 1023
rect 282 1013 285 1326
rect 298 1316 301 1396
rect 306 1393 309 1446
rect 306 1333 309 1366
rect 314 1323 317 1436
rect 322 1383 325 1456
rect 330 1413 333 1503
rect 338 1463 341 1746
rect 338 1373 341 1446
rect 338 1326 341 1356
rect 334 1323 341 1326
rect 298 1313 325 1316
rect 290 1143 293 1286
rect 298 1196 301 1256
rect 298 1193 305 1196
rect 290 1123 293 1136
rect 302 1126 305 1193
rect 302 1123 309 1126
rect 290 1086 293 1116
rect 298 1103 301 1116
rect 290 1083 297 1086
rect 294 1016 297 1083
rect 306 1023 309 1123
rect 314 1086 317 1186
rect 322 1103 325 1313
rect 334 1246 337 1323
rect 334 1243 341 1246
rect 330 1213 333 1226
rect 338 1203 341 1243
rect 330 1113 333 1126
rect 314 1083 325 1086
rect 294 1013 309 1016
rect 250 993 253 1006
rect 250 933 253 956
rect 250 916 253 926
rect 258 923 261 936
rect 266 916 269 1006
rect 274 923 277 946
rect 250 913 269 916
rect 250 896 253 913
rect 282 906 285 966
rect 290 933 293 946
rect 298 916 301 956
rect 278 903 285 906
rect 294 913 301 916
rect 250 893 257 896
rect 254 836 257 893
rect 250 833 257 836
rect 250 723 253 833
rect 258 793 261 816
rect 242 553 245 716
rect 250 693 253 706
rect 250 543 253 616
rect 242 516 245 526
rect 250 523 253 536
rect 258 516 261 786
rect 266 563 269 856
rect 278 846 281 903
rect 274 843 281 846
rect 274 826 277 843
rect 294 826 297 913
rect 274 823 285 826
rect 294 823 301 826
rect 274 803 277 816
rect 282 806 285 823
rect 282 803 289 806
rect 274 623 277 796
rect 286 746 289 803
rect 282 743 289 746
rect 282 713 285 743
rect 290 713 293 726
rect 242 513 261 516
rect 266 513 269 526
rect 234 503 245 506
rect 202 433 213 436
rect 170 416 173 433
rect 122 393 141 396
rect 114 363 125 366
rect 106 333 117 336
rect 90 323 97 326
rect 66 313 77 316
rect 74 236 77 313
rect 66 233 77 236
rect 66 143 69 233
rect 90 203 93 323
rect 106 313 109 326
rect 114 306 117 333
rect 122 313 125 363
rect 130 343 133 366
rect 130 326 133 336
rect 138 333 141 393
rect 130 323 149 326
rect 154 306 157 416
rect 114 303 157 306
rect 162 413 173 416
rect 186 413 189 426
rect 114 203 117 303
rect 162 286 165 413
rect 154 283 165 286
rect 154 236 157 283
rect 154 233 165 236
rect 122 133 125 216
rect 162 196 165 233
rect 154 193 165 196
rect 170 193 173 206
rect 154 126 157 193
rect 154 123 165 126
rect 178 123 181 336
rect 194 233 197 426
rect 210 346 213 433
rect 242 413 245 503
rect 258 413 261 436
rect 226 396 229 406
rect 266 396 269 416
rect 274 403 277 616
rect 282 593 285 606
rect 290 603 293 626
rect 298 613 301 823
rect 306 793 309 1013
rect 322 936 325 1083
rect 338 1023 341 1116
rect 346 1006 349 2113
rect 362 2106 365 2306
rect 386 2236 389 2343
rect 418 2333 421 2383
rect 426 2323 429 2336
rect 370 2233 389 2236
rect 370 2123 373 2233
rect 378 2206 381 2226
rect 394 2213 397 2226
rect 378 2203 397 2206
rect 386 2123 389 2136
rect 394 2123 397 2203
rect 418 2166 421 2236
rect 426 2213 429 2226
rect 434 2203 437 2316
rect 466 2293 469 2516
rect 474 2376 477 2416
rect 506 2413 509 2523
rect 514 2516 517 2526
rect 530 2523 533 2593
rect 554 2586 557 2633
rect 578 2603 581 2616
rect 610 2613 613 2663
rect 626 2623 629 2833
rect 634 2793 637 2816
rect 666 2813 669 2836
rect 642 2723 645 2806
rect 658 2793 661 2806
rect 674 2743 677 2846
rect 682 2813 685 2826
rect 738 2823 741 2896
rect 650 2626 653 2736
rect 674 2656 677 2736
rect 690 2726 693 2746
rect 698 2733 701 2806
rect 706 2736 709 2816
rect 714 2786 717 2806
rect 738 2793 741 2806
rect 746 2786 749 2836
rect 754 2826 757 2926
rect 762 2923 765 2936
rect 770 2923 773 2943
rect 778 2833 781 2936
rect 786 2913 789 2926
rect 794 2896 797 3043
rect 810 3023 821 3026
rect 858 3023 861 3113
rect 874 3026 877 3183
rect 914 3176 917 3253
rect 922 3216 925 3246
rect 930 3223 933 3236
rect 946 3216 949 3226
rect 922 3213 933 3216
rect 882 3173 917 3176
rect 930 3173 933 3213
rect 882 3116 885 3173
rect 890 3143 893 3166
rect 898 3143 901 3156
rect 890 3126 893 3136
rect 890 3123 901 3126
rect 882 3113 893 3116
rect 874 3023 885 3026
rect 802 2963 805 3016
rect 834 3003 837 3016
rect 802 2903 805 2916
rect 794 2893 805 2896
rect 754 2823 789 2826
rect 714 2783 749 2786
rect 754 2796 757 2816
rect 786 2803 789 2816
rect 754 2793 797 2796
rect 706 2733 733 2736
rect 690 2723 709 2726
rect 674 2653 709 2656
rect 646 2623 653 2626
rect 554 2583 565 2586
rect 538 2516 541 2536
rect 562 2523 565 2583
rect 646 2576 649 2623
rect 634 2573 649 2576
rect 626 2533 629 2556
rect 514 2513 541 2516
rect 610 2433 613 2526
rect 634 2506 637 2573
rect 658 2556 661 2616
rect 682 2603 685 2616
rect 706 2613 709 2653
rect 650 2553 661 2556
rect 642 2533 645 2546
rect 650 2523 653 2553
rect 722 2533 725 2646
rect 618 2503 637 2506
rect 474 2373 485 2376
rect 538 2373 541 2406
rect 482 2333 485 2373
rect 506 2323 509 2336
rect 514 2313 517 2336
rect 530 2313 533 2326
rect 466 2223 477 2226
rect 402 2163 421 2166
rect 358 2103 365 2106
rect 358 2026 361 2103
rect 370 2086 373 2116
rect 370 2083 381 2086
rect 358 2023 365 2026
rect 354 1873 357 2006
rect 362 1903 365 2023
rect 370 1923 373 2066
rect 378 2033 381 2083
rect 402 2056 405 2163
rect 394 2053 405 2056
rect 378 2006 381 2026
rect 378 2003 389 2006
rect 378 1923 381 1936
rect 386 1923 389 2003
rect 394 1973 397 2053
rect 410 2046 413 2126
rect 402 2043 413 2046
rect 402 2003 405 2043
rect 410 2023 413 2036
rect 410 1983 413 2016
rect 354 1823 373 1826
rect 354 1803 357 1816
rect 354 1633 357 1726
rect 354 1536 357 1626
rect 362 1546 365 1736
rect 370 1623 373 1823
rect 394 1813 397 1936
rect 410 1906 413 1976
rect 406 1903 413 1906
rect 406 1836 409 1903
rect 402 1833 409 1836
rect 402 1753 405 1833
rect 410 1813 413 1826
rect 370 1583 373 1616
rect 378 1553 381 1746
rect 418 1743 421 2156
rect 442 2136 445 2206
rect 426 1933 429 2136
rect 442 2133 449 2136
rect 434 2063 437 2126
rect 446 2056 449 2133
rect 442 2053 449 2056
rect 442 2026 445 2053
rect 458 2036 461 2136
rect 466 2123 469 2223
rect 474 2043 477 2136
rect 434 2023 445 2026
rect 434 1933 437 2023
rect 434 1816 437 1926
rect 442 1906 445 2016
rect 450 2006 453 2036
rect 458 2033 477 2036
rect 466 2013 469 2026
rect 450 2003 469 2006
rect 466 1963 469 2003
rect 458 1933 461 1946
rect 474 1933 477 2033
rect 482 1973 485 2206
rect 490 2043 493 2216
rect 450 1913 453 1926
rect 442 1903 449 1906
rect 446 1836 449 1903
rect 466 1866 469 1926
rect 458 1863 469 1866
rect 446 1833 453 1836
rect 426 1746 429 1816
rect 434 1813 445 1816
rect 442 1756 445 1813
rect 450 1803 453 1833
rect 458 1803 461 1863
rect 474 1813 477 1926
rect 474 1786 477 1806
rect 470 1783 477 1786
rect 442 1753 453 1756
rect 426 1743 445 1746
rect 362 1543 373 1546
rect 354 1533 365 1536
rect 362 1513 365 1533
rect 354 1413 357 1486
rect 354 1393 357 1406
rect 354 1193 357 1376
rect 362 1353 365 1426
rect 370 1346 373 1543
rect 378 1523 381 1546
rect 378 1463 381 1516
rect 378 1413 381 1456
rect 386 1413 389 1736
rect 394 1713 397 1736
rect 410 1733 437 1736
rect 410 1726 413 1733
rect 402 1723 413 1726
rect 418 1723 429 1726
rect 410 1663 413 1706
rect 418 1703 421 1716
rect 394 1583 397 1646
rect 362 1343 373 1346
rect 354 1103 357 1176
rect 314 933 325 936
rect 338 1003 349 1006
rect 354 1003 357 1026
rect 338 936 341 1003
rect 354 953 357 996
rect 338 933 349 936
rect 314 803 317 933
rect 322 853 325 916
rect 338 893 341 916
rect 330 823 333 836
rect 306 703 309 776
rect 330 746 333 806
rect 338 793 341 816
rect 330 743 341 746
rect 322 733 333 736
rect 306 593 309 616
rect 314 613 317 726
rect 322 713 325 733
rect 282 523 285 536
rect 290 506 293 576
rect 322 573 325 626
rect 330 566 333 636
rect 338 603 341 743
rect 346 653 349 933
rect 354 923 357 936
rect 354 903 357 916
rect 354 813 357 896
rect 346 613 349 626
rect 354 603 357 786
rect 298 513 301 536
rect 306 506 309 546
rect 314 533 317 566
rect 322 563 333 566
rect 286 503 293 506
rect 298 503 309 506
rect 226 393 269 396
rect 202 343 213 346
rect 202 316 205 343
rect 226 333 229 386
rect 210 323 229 326
rect 202 313 229 316
rect 226 303 229 313
rect 234 246 237 393
rect 286 386 289 503
rect 298 396 301 503
rect 314 406 317 476
rect 306 403 317 406
rect 298 393 309 396
rect 266 383 289 386
rect 266 366 269 383
rect 258 363 269 366
rect 242 333 245 356
rect 258 286 261 363
rect 258 283 269 286
rect 274 283 277 336
rect 226 243 237 246
rect 186 213 189 226
rect 194 203 197 216
rect 226 186 229 243
rect 250 213 253 236
rect 250 196 253 206
rect 258 203 261 266
rect 266 213 269 283
rect 282 196 285 216
rect 290 203 293 326
rect 298 313 301 346
rect 306 296 309 393
rect 314 323 317 403
rect 322 316 325 563
rect 330 486 333 536
rect 338 503 341 526
rect 354 513 357 576
rect 346 493 349 506
rect 330 483 337 486
rect 334 356 337 483
rect 362 473 365 1343
rect 370 1253 373 1336
rect 370 1056 373 1246
rect 378 1173 381 1376
rect 386 1343 389 1396
rect 386 1323 389 1336
rect 386 1213 389 1256
rect 394 1166 397 1556
rect 402 1393 405 1606
rect 418 1546 421 1676
rect 410 1543 421 1546
rect 410 1533 413 1543
rect 410 1443 413 1526
rect 418 1473 421 1536
rect 426 1523 429 1723
rect 434 1713 437 1733
rect 442 1703 445 1743
rect 450 1723 453 1753
rect 458 1696 461 1756
rect 470 1706 473 1783
rect 470 1703 477 1706
rect 454 1693 461 1696
rect 454 1636 457 1693
rect 434 1613 437 1636
rect 454 1633 461 1636
rect 442 1566 445 1606
rect 434 1563 445 1566
rect 434 1533 437 1563
rect 450 1543 453 1586
rect 458 1536 461 1633
rect 442 1533 461 1536
rect 442 1526 445 1533
rect 434 1523 445 1526
rect 410 1423 421 1426
rect 426 1416 429 1466
rect 434 1453 437 1523
rect 410 1373 413 1416
rect 418 1413 429 1416
rect 434 1413 437 1426
rect 418 1356 421 1413
rect 410 1353 421 1356
rect 402 1316 405 1336
rect 410 1326 413 1353
rect 418 1333 421 1346
rect 426 1343 429 1406
rect 442 1403 445 1476
rect 450 1386 453 1466
rect 442 1383 453 1386
rect 410 1323 421 1326
rect 402 1313 413 1316
rect 410 1283 413 1313
rect 418 1276 421 1323
rect 378 1163 397 1166
rect 402 1273 421 1276
rect 378 1106 381 1163
rect 386 1133 389 1146
rect 394 1113 397 1126
rect 378 1103 397 1106
rect 370 1053 389 1056
rect 370 1013 373 1026
rect 378 1003 381 1046
rect 386 996 389 1053
rect 370 993 389 996
rect 370 913 373 993
rect 394 976 397 1103
rect 402 1096 405 1273
rect 410 1203 413 1216
rect 418 1203 421 1216
rect 410 1136 413 1196
rect 410 1133 421 1136
rect 410 1103 413 1126
rect 418 1123 421 1133
rect 426 1126 429 1326
rect 442 1316 445 1383
rect 442 1313 453 1316
rect 450 1293 453 1313
rect 458 1283 461 1526
rect 434 1143 437 1226
rect 442 1196 445 1206
rect 450 1203 461 1206
rect 466 1196 469 1686
rect 474 1613 477 1703
rect 482 1613 485 1966
rect 490 1893 493 2016
rect 498 1996 501 2246
rect 522 2223 533 2226
rect 514 2193 517 2206
rect 522 2186 525 2223
rect 538 2216 541 2306
rect 514 2183 525 2186
rect 530 2213 541 2216
rect 506 2033 509 2106
rect 514 2026 517 2183
rect 522 2123 525 2176
rect 506 2023 517 2026
rect 522 2023 525 2036
rect 506 2013 509 2023
rect 498 1993 505 1996
rect 502 1906 505 1993
rect 514 1976 517 2023
rect 530 1983 533 2213
rect 546 2153 549 2316
rect 538 2103 541 2116
rect 546 2013 549 2126
rect 554 2006 557 2346
rect 570 2333 573 2416
rect 562 2276 565 2296
rect 562 2273 569 2276
rect 566 2146 569 2273
rect 578 2213 581 2256
rect 586 2213 589 2336
rect 602 2333 613 2336
rect 594 2223 597 2326
rect 610 2233 613 2316
rect 618 2293 621 2503
rect 626 2413 629 2496
rect 714 2453 717 2526
rect 730 2506 733 2733
rect 738 2723 741 2736
rect 754 2723 757 2793
rect 778 2723 781 2766
rect 802 2733 805 2893
rect 818 2723 821 2796
rect 826 2616 829 2996
rect 834 2923 837 2936
rect 850 2913 853 2926
rect 858 2923 861 3016
rect 866 2993 869 3006
rect 882 2986 885 3023
rect 890 2993 893 3113
rect 898 3093 901 3123
rect 906 3106 909 3136
rect 914 3123 917 3146
rect 906 3103 913 3106
rect 910 3046 913 3103
rect 910 3043 917 3046
rect 898 2986 901 3016
rect 882 2983 901 2986
rect 882 2946 885 2983
rect 866 2943 885 2946
rect 866 2933 869 2943
rect 842 2803 845 2816
rect 850 2803 853 2846
rect 866 2823 869 2926
rect 858 2783 861 2806
rect 866 2753 869 2816
rect 738 2533 741 2546
rect 746 2533 749 2586
rect 762 2556 765 2616
rect 794 2603 797 2616
rect 818 2613 829 2616
rect 842 2613 845 2676
rect 874 2626 877 2936
rect 882 2923 885 2943
rect 882 2823 885 2916
rect 890 2833 893 2956
rect 906 2936 909 3036
rect 914 2953 917 3043
rect 922 3013 925 3066
rect 930 3003 933 3136
rect 938 3106 941 3216
rect 946 3213 957 3216
rect 962 3213 965 3236
rect 970 3156 973 3323
rect 1026 3323 1037 3326
rect 1026 3256 1029 3323
rect 1026 3253 1037 3256
rect 1034 3236 1037 3253
rect 1034 3233 1045 3236
rect 1018 3223 1037 3226
rect 946 3133 949 3146
rect 954 3123 957 3156
rect 966 3153 973 3156
rect 986 3213 1021 3216
rect 966 3106 969 3153
rect 978 3123 981 3146
rect 986 3113 989 3213
rect 994 3193 997 3206
rect 1010 3136 1013 3156
rect 1018 3146 1021 3206
rect 1026 3173 1029 3206
rect 1034 3183 1037 3223
rect 1042 3163 1045 3233
rect 1018 3143 1037 3146
rect 994 3133 1013 3136
rect 1034 3133 1037 3143
rect 938 3103 949 3106
rect 966 3103 973 3106
rect 946 3046 949 3103
rect 938 3043 949 3046
rect 970 3086 973 3103
rect 970 3083 989 3086
rect 938 3023 941 3043
rect 954 3013 965 3016
rect 970 2963 973 3083
rect 906 2933 917 2936
rect 906 2913 909 2926
rect 914 2843 917 2933
rect 922 2913 925 2946
rect 954 2923 965 2926
rect 882 2793 885 2806
rect 922 2756 925 2806
rect 930 2793 933 2846
rect 946 2803 949 2886
rect 970 2826 973 2926
rect 978 2886 981 2996
rect 986 2893 989 3006
rect 1002 3003 1005 3056
rect 1010 3023 1013 3126
rect 1026 3066 1029 3126
rect 1034 3123 1045 3126
rect 1026 3063 1037 3066
rect 1026 3016 1029 3046
rect 1034 3023 1037 3063
rect 1018 2996 1021 3016
rect 1026 3013 1037 3016
rect 1050 3013 1053 3340
rect 1066 3326 1069 3340
rect 1066 3323 1077 3326
rect 1074 3276 1077 3323
rect 1066 3273 1077 3276
rect 1066 3256 1069 3273
rect 1066 3253 1085 3256
rect 1058 3093 1061 3216
rect 1066 3053 1069 3216
rect 1074 3213 1077 3246
rect 1082 3216 1085 3253
rect 1082 3213 1093 3216
rect 1074 3193 1077 3206
rect 1034 3003 1037 3013
rect 1042 2996 1045 3006
rect 1018 2993 1045 2996
rect 994 2933 1005 2936
rect 994 2886 997 2926
rect 978 2883 997 2886
rect 1002 2883 1005 2933
rect 1010 2843 1013 2926
rect 1018 2913 1021 2936
rect 1042 2846 1045 2993
rect 1074 2983 1077 3166
rect 1090 3156 1093 3213
rect 1082 3153 1093 3156
rect 1082 3013 1085 3153
rect 1106 3136 1109 3340
rect 1162 3293 1173 3296
rect 1122 3203 1125 3216
rect 1130 3213 1133 3246
rect 1146 3203 1149 3226
rect 1162 3223 1165 3246
rect 1170 3223 1173 3293
rect 1186 3206 1189 3340
rect 1178 3203 1189 3206
rect 1090 3133 1109 3136
rect 1090 3113 1093 3133
rect 1114 3126 1117 3136
rect 1122 3133 1125 3156
rect 1146 3133 1149 3146
rect 1098 3076 1101 3126
rect 1106 3123 1117 3126
rect 1106 3103 1109 3123
rect 1098 3073 1109 3076
rect 1090 3063 1101 3066
rect 1098 3013 1101 3063
rect 1106 3006 1109 3073
rect 1114 3063 1117 3116
rect 1082 3003 1109 3006
rect 1122 3003 1125 3126
rect 1130 3003 1133 3106
rect 1138 3063 1141 3126
rect 1154 3053 1157 3136
rect 1178 3116 1181 3203
rect 1194 3193 1197 3216
rect 1202 3176 1205 3256
rect 1210 3213 1213 3236
rect 1218 3233 1253 3236
rect 1226 3203 1229 3226
rect 1250 3216 1253 3233
rect 1234 3183 1237 3216
rect 1250 3213 1261 3216
rect 1242 3176 1245 3206
rect 1258 3203 1261 3213
rect 1202 3173 1245 3176
rect 1194 3123 1197 3156
rect 1202 3123 1205 3173
rect 1210 3133 1221 3136
rect 1226 3133 1229 3166
rect 1250 3133 1253 3146
rect 1210 3123 1221 3126
rect 1178 3113 1189 3116
rect 1186 3073 1189 3113
rect 1210 3083 1213 3123
rect 1242 3116 1245 3126
rect 1218 3113 1245 3116
rect 1266 3053 1269 3216
rect 1290 3213 1293 3256
rect 1298 3213 1301 3246
rect 1306 3206 1309 3236
rect 1274 3203 1293 3206
rect 1298 3203 1309 3206
rect 1274 3193 1277 3203
rect 1298 3176 1301 3203
rect 1290 3173 1301 3176
rect 1290 3106 1293 3173
rect 1306 3113 1309 3126
rect 1314 3123 1317 3206
rect 1322 3203 1333 3206
rect 1338 3173 1341 3216
rect 1378 3213 1381 3236
rect 1354 3186 1357 3206
rect 1354 3183 1365 3186
rect 1330 3126 1333 3136
rect 1338 3133 1341 3166
rect 1362 3133 1365 3183
rect 1378 3166 1381 3186
rect 1374 3163 1381 3166
rect 1322 3123 1333 3126
rect 1290 3103 1301 3106
rect 1322 3103 1325 3123
rect 1146 3023 1173 3026
rect 1146 3016 1149 3023
rect 1138 3013 1149 3016
rect 1042 2843 1053 2846
rect 970 2823 981 2826
rect 954 2783 957 2806
rect 898 2743 901 2756
rect 922 2753 933 2756
rect 962 2753 965 2816
rect 906 2673 909 2736
rect 914 2723 917 2746
rect 930 2636 933 2753
rect 962 2723 965 2736
rect 986 2723 989 2806
rect 1026 2783 1029 2806
rect 1050 2766 1053 2843
rect 1042 2763 1053 2766
rect 1042 2716 1045 2763
rect 1066 2723 1069 2966
rect 1098 2856 1101 3003
rect 1146 2983 1149 3006
rect 1154 2973 1157 3016
rect 1114 2923 1117 2946
rect 1138 2933 1165 2936
rect 1138 2906 1141 2933
rect 1146 2913 1149 2926
rect 1138 2903 1149 2906
rect 1154 2903 1157 2926
rect 1162 2906 1165 2933
rect 1170 2926 1173 3023
rect 1178 3013 1181 3026
rect 1186 2993 1189 3006
rect 1178 2933 1181 2946
rect 1170 2923 1181 2926
rect 1178 2913 1181 2923
rect 1186 2906 1189 2936
rect 1162 2903 1189 2906
rect 1098 2853 1109 2856
rect 1074 2793 1077 2816
rect 1106 2776 1109 2853
rect 1098 2773 1109 2776
rect 1042 2713 1053 2716
rect 866 2623 877 2626
rect 922 2633 933 2636
rect 754 2553 765 2556
rect 754 2523 757 2553
rect 730 2503 741 2506
rect 738 2446 741 2503
rect 762 2493 765 2526
rect 818 2456 821 2613
rect 866 2576 869 2623
rect 866 2573 877 2576
rect 858 2523 861 2546
rect 866 2533 869 2556
rect 874 2526 877 2573
rect 882 2546 885 2616
rect 922 2613 925 2633
rect 898 2593 901 2606
rect 882 2543 909 2546
rect 882 2533 893 2536
rect 866 2483 869 2526
rect 874 2523 893 2526
rect 898 2523 901 2536
rect 906 2523 909 2543
rect 914 2533 917 2586
rect 818 2453 825 2456
rect 734 2443 741 2446
rect 642 2393 645 2406
rect 626 2323 629 2336
rect 682 2333 685 2416
rect 722 2413 725 2436
rect 690 2323 693 2336
rect 634 2296 637 2316
rect 714 2313 717 2346
rect 634 2293 645 2296
rect 538 1976 541 2006
rect 514 1973 541 1976
rect 546 2003 557 2006
rect 562 2143 569 2146
rect 514 1923 517 1946
rect 522 1923 525 1936
rect 530 1906 533 1926
rect 538 1913 541 1936
rect 502 1903 509 1906
rect 506 1836 509 1903
rect 522 1903 533 1906
rect 522 1846 525 1903
rect 522 1843 533 1846
rect 498 1833 509 1836
rect 490 1763 493 1816
rect 490 1733 493 1746
rect 498 1673 501 1833
rect 530 1823 533 1843
rect 506 1803 509 1816
rect 514 1803 517 1816
rect 522 1763 525 1806
rect 506 1646 509 1746
rect 514 1723 517 1746
rect 522 1723 525 1736
rect 530 1716 533 1816
rect 538 1743 541 1896
rect 546 1763 549 2003
rect 554 1923 557 1976
rect 562 1923 565 2143
rect 570 2083 573 2126
rect 570 2013 573 2026
rect 570 1993 573 2006
rect 570 1933 573 1946
rect 578 1913 581 2136
rect 586 2123 589 2206
rect 602 2193 605 2216
rect 594 2043 597 2136
rect 602 2133 605 2166
rect 602 2093 605 2126
rect 586 1926 589 2016
rect 602 2013 605 2086
rect 594 1943 597 1986
rect 586 1923 593 1926
rect 602 1923 605 1956
rect 554 1813 557 1896
rect 562 1796 565 1856
rect 570 1803 573 1816
rect 578 1813 581 1876
rect 590 1816 593 1923
rect 602 1823 605 1876
rect 590 1813 605 1816
rect 558 1793 565 1796
rect 522 1713 533 1716
rect 522 1656 525 1713
rect 538 1673 541 1726
rect 558 1716 561 1793
rect 570 1723 573 1766
rect 586 1733 589 1806
rect 594 1733 597 1806
rect 602 1726 605 1813
rect 546 1713 561 1716
rect 490 1643 509 1646
rect 514 1653 525 1656
rect 474 1503 477 1546
rect 474 1423 477 1456
rect 474 1223 477 1416
rect 482 1306 485 1606
rect 490 1543 493 1643
rect 514 1636 517 1653
rect 506 1633 517 1636
rect 506 1603 509 1633
rect 514 1623 533 1626
rect 490 1473 493 1526
rect 498 1453 501 1596
rect 490 1323 493 1416
rect 498 1403 501 1426
rect 506 1416 509 1526
rect 514 1426 517 1623
rect 522 1433 525 1616
rect 530 1603 533 1616
rect 530 1483 533 1536
rect 538 1523 541 1646
rect 546 1623 549 1713
rect 554 1686 557 1706
rect 554 1683 561 1686
rect 558 1616 561 1683
rect 558 1613 565 1616
rect 570 1613 573 1696
rect 546 1516 549 1586
rect 554 1523 557 1606
rect 542 1513 549 1516
rect 514 1423 525 1426
rect 506 1413 517 1416
rect 530 1413 533 1466
rect 542 1456 545 1513
rect 538 1453 545 1456
rect 514 1403 517 1413
rect 514 1346 517 1396
rect 506 1343 517 1346
rect 498 1306 501 1336
rect 506 1323 509 1343
rect 482 1303 489 1306
rect 498 1303 509 1306
rect 486 1246 489 1303
rect 486 1243 493 1246
rect 474 1213 485 1216
rect 442 1193 453 1196
rect 426 1123 433 1126
rect 418 1096 421 1116
rect 402 1093 421 1096
rect 402 993 405 1006
rect 394 973 401 976
rect 386 943 389 956
rect 378 923 381 936
rect 370 813 373 836
rect 378 806 381 886
rect 374 803 381 806
rect 374 736 377 803
rect 370 733 377 736
rect 370 703 373 733
rect 378 703 381 716
rect 370 613 373 696
rect 378 606 381 696
rect 370 603 381 606
rect 370 503 373 603
rect 378 513 381 596
rect 362 426 365 466
rect 386 436 389 936
rect 398 816 401 973
rect 394 813 401 816
rect 394 763 397 813
rect 402 783 405 796
rect 410 753 413 1093
rect 418 806 421 1076
rect 430 946 433 1123
rect 442 1023 445 1166
rect 450 1133 453 1193
rect 458 1193 469 1196
rect 474 1193 477 1206
rect 458 1116 461 1193
rect 482 1186 485 1213
rect 490 1193 493 1243
rect 466 1183 485 1186
rect 466 1123 469 1183
rect 458 1113 469 1116
rect 442 993 445 1016
rect 450 973 453 1006
rect 426 943 433 946
rect 426 913 429 943
rect 426 813 429 856
rect 418 803 429 806
rect 434 803 437 926
rect 458 923 461 966
rect 442 823 445 906
rect 458 903 461 916
rect 466 903 469 1113
rect 474 953 477 996
rect 482 936 485 1086
rect 478 933 485 936
rect 450 816 453 866
rect 442 813 453 816
rect 458 813 461 826
rect 410 726 413 736
rect 394 723 413 726
rect 394 713 405 716
rect 418 713 421 796
rect 394 646 397 713
rect 426 706 429 803
rect 434 713 437 736
rect 442 706 445 813
rect 450 733 453 796
rect 422 703 429 706
rect 434 703 445 706
rect 450 703 453 716
rect 394 643 405 646
rect 394 523 397 606
rect 402 573 405 643
rect 410 483 413 686
rect 422 556 425 703
rect 434 613 437 703
rect 458 686 461 806
rect 466 783 469 816
rect 478 776 481 933
rect 490 823 493 1176
rect 498 1163 501 1216
rect 498 1146 501 1156
rect 506 1153 509 1296
rect 514 1233 517 1336
rect 498 1143 509 1146
rect 498 1073 501 1136
rect 498 1003 501 1066
rect 506 1053 509 1143
rect 514 1123 517 1216
rect 522 1183 525 1386
rect 538 1366 541 1453
rect 546 1383 549 1436
rect 530 1363 541 1366
rect 522 1056 525 1156
rect 530 1063 533 1363
rect 546 1323 549 1376
rect 554 1316 557 1506
rect 542 1313 557 1316
rect 542 1206 545 1313
rect 562 1286 565 1613
rect 570 1503 573 1556
rect 578 1503 581 1726
rect 598 1723 605 1726
rect 586 1613 589 1716
rect 598 1656 601 1723
rect 594 1653 601 1656
rect 570 1443 573 1496
rect 578 1416 581 1476
rect 586 1423 589 1606
rect 594 1583 597 1653
rect 602 1576 605 1636
rect 594 1573 605 1576
rect 594 1546 597 1573
rect 602 1553 605 1566
rect 594 1543 605 1546
rect 594 1513 597 1536
rect 602 1496 605 1543
rect 594 1493 605 1496
rect 594 1473 597 1493
rect 570 1393 573 1416
rect 578 1413 589 1416
rect 578 1373 581 1406
rect 586 1346 589 1413
rect 578 1343 589 1346
rect 570 1303 573 1326
rect 542 1203 549 1206
rect 522 1053 533 1056
rect 506 1013 517 1016
rect 506 1003 525 1006
rect 498 803 501 916
rect 506 813 509 1003
rect 530 996 533 1053
rect 514 993 533 996
rect 514 876 517 993
rect 522 926 525 946
rect 522 923 533 926
rect 538 906 541 1146
rect 546 1073 549 1203
rect 546 923 549 1056
rect 554 1026 557 1286
rect 562 1283 569 1286
rect 566 1226 569 1283
rect 566 1223 573 1226
rect 562 1203 565 1216
rect 562 1043 565 1146
rect 570 1133 573 1223
rect 578 1153 581 1343
rect 586 1203 589 1336
rect 594 1323 597 1426
rect 594 1273 597 1316
rect 586 1126 589 1166
rect 570 1106 573 1126
rect 578 1123 589 1126
rect 594 1113 597 1176
rect 570 1103 581 1106
rect 578 1036 581 1103
rect 570 1033 581 1036
rect 554 1023 561 1026
rect 558 946 561 1023
rect 554 943 561 946
rect 538 903 545 906
rect 514 873 533 876
rect 466 773 481 776
rect 466 733 469 773
rect 474 763 509 766
rect 474 706 477 763
rect 442 683 461 686
rect 470 703 477 706
rect 442 613 445 683
rect 470 636 473 703
rect 482 693 485 756
rect 470 633 477 636
rect 442 593 445 606
rect 458 556 461 616
rect 418 553 425 556
rect 434 553 461 556
rect 418 533 421 553
rect 434 536 437 553
rect 442 543 461 546
rect 426 526 429 536
rect 434 533 445 536
rect 418 523 429 526
rect 442 436 445 526
rect 458 523 461 543
rect 466 523 469 616
rect 474 613 477 633
rect 474 516 477 586
rect 346 423 365 426
rect 378 433 389 436
rect 378 416 381 433
rect 410 423 413 436
rect 418 433 445 436
rect 458 513 477 516
rect 458 423 461 513
rect 482 483 485 656
rect 490 603 493 726
rect 498 723 501 736
rect 506 733 509 763
rect 498 676 501 696
rect 498 673 505 676
rect 502 596 505 673
rect 514 603 517 826
rect 522 773 525 816
rect 530 813 533 873
rect 542 826 545 903
rect 538 823 545 826
rect 522 723 525 746
rect 530 706 533 766
rect 526 703 533 706
rect 526 606 529 703
rect 526 603 533 606
rect 498 593 505 596
rect 498 546 501 593
rect 490 543 501 546
rect 490 476 493 543
rect 498 506 501 536
rect 514 523 517 596
rect 530 583 533 603
rect 538 593 541 823
rect 546 733 549 806
rect 554 726 557 943
rect 562 823 565 926
rect 562 793 565 806
rect 546 723 557 726
rect 546 613 549 723
rect 562 713 565 736
rect 570 696 573 1033
rect 594 1023 597 1106
rect 578 826 581 1006
rect 586 923 589 1016
rect 594 833 597 1016
rect 578 823 589 826
rect 578 803 581 816
rect 562 693 573 696
rect 562 636 565 693
rect 562 633 573 636
rect 570 613 573 633
rect 546 573 549 606
rect 538 546 541 566
rect 538 543 549 546
rect 554 536 557 606
rect 578 583 581 776
rect 586 723 589 823
rect 594 773 597 826
rect 594 706 597 736
rect 590 703 597 706
rect 590 636 593 703
rect 586 633 593 636
rect 522 533 541 536
rect 498 503 517 506
rect 466 473 493 476
rect 302 293 309 296
rect 314 313 325 316
rect 330 353 337 356
rect 374 413 381 416
rect 302 226 305 293
rect 302 223 309 226
rect 306 206 309 223
rect 314 213 317 313
rect 330 256 333 353
rect 374 346 377 413
rect 386 373 389 416
rect 410 403 413 416
rect 374 343 381 346
rect 338 263 341 336
rect 362 323 365 336
rect 378 323 381 343
rect 386 323 389 336
rect 394 316 397 326
rect 354 313 397 316
rect 330 253 373 256
rect 330 223 333 253
rect 346 243 365 246
rect 346 233 349 243
rect 338 213 349 216
rect 306 203 317 206
rect 250 193 285 196
rect 226 183 237 186
rect 226 123 229 136
rect 234 133 237 183
rect 258 133 261 193
rect 162 103 165 123
rect 226 113 237 116
rect 234 76 237 113
rect 250 76 253 126
rect 314 106 317 203
rect 322 123 325 136
rect 330 133 333 166
rect 354 133 357 236
rect 362 183 365 243
rect 370 223 373 253
rect 410 223 413 336
rect 434 323 437 336
rect 442 263 445 416
rect 450 323 453 346
rect 458 333 461 376
rect 466 333 469 473
rect 482 413 485 436
rect 474 343 477 406
rect 490 373 493 406
rect 498 336 501 416
rect 506 393 509 446
rect 514 403 517 503
rect 538 493 541 533
rect 546 533 557 536
rect 474 323 477 336
rect 482 333 501 336
rect 482 313 485 333
rect 498 313 501 326
rect 514 323 517 336
rect 522 316 525 456
rect 546 446 549 533
rect 554 503 557 526
rect 538 443 549 446
rect 538 366 541 443
rect 562 436 565 566
rect 570 536 573 556
rect 586 543 589 633
rect 602 613 605 1486
rect 610 1356 613 2186
rect 618 1993 621 2256
rect 642 2226 645 2293
rect 626 2143 629 2226
rect 634 2223 645 2226
rect 626 2073 629 2126
rect 618 1553 621 1936
rect 626 1833 629 2006
rect 626 1613 629 1826
rect 634 1626 637 2223
rect 674 2213 677 2286
rect 682 2213 685 2246
rect 722 2213 725 2386
rect 734 2346 737 2443
rect 754 2393 757 2406
rect 730 2343 737 2346
rect 730 2326 733 2343
rect 778 2333 781 2416
rect 822 2376 825 2453
rect 834 2413 837 2456
rect 890 2446 893 2523
rect 954 2493 957 2526
rect 890 2443 901 2446
rect 866 2393 869 2406
rect 898 2396 901 2443
rect 890 2393 901 2396
rect 818 2373 825 2376
rect 730 2323 749 2326
rect 778 2313 781 2326
rect 786 2233 789 2336
rect 810 2273 813 2316
rect 818 2313 821 2373
rect 834 2333 837 2356
rect 834 2246 837 2266
rect 842 2253 845 2336
rect 866 2333 869 2346
rect 882 2333 885 2346
rect 834 2243 845 2246
rect 738 2223 805 2226
rect 738 2213 741 2223
rect 642 2166 645 2206
rect 658 2173 661 2196
rect 642 2163 653 2166
rect 666 2153 669 2206
rect 642 2123 645 2136
rect 666 2123 669 2146
rect 674 2133 677 2166
rect 682 2133 685 2196
rect 642 2103 645 2116
rect 642 1983 645 2016
rect 650 2003 653 2036
rect 642 1823 645 1926
rect 650 1893 653 1936
rect 658 1923 661 2016
rect 666 2003 669 2016
rect 674 1996 677 2116
rect 682 2103 685 2126
rect 682 2013 685 2046
rect 690 2003 693 2126
rect 674 1993 693 1996
rect 666 1926 669 1936
rect 666 1923 677 1926
rect 650 1816 653 1836
rect 642 1813 653 1816
rect 650 1756 653 1813
rect 642 1753 653 1756
rect 642 1636 645 1736
rect 650 1723 653 1746
rect 650 1643 653 1716
rect 642 1633 653 1636
rect 634 1623 645 1626
rect 626 1583 629 1606
rect 634 1556 637 1616
rect 626 1553 637 1556
rect 618 1513 621 1546
rect 618 1406 621 1506
rect 626 1483 629 1553
rect 642 1546 645 1623
rect 650 1603 653 1633
rect 658 1596 661 1906
rect 666 1853 669 1886
rect 666 1813 669 1826
rect 666 1743 669 1776
rect 666 1643 669 1736
rect 674 1733 677 1806
rect 682 1776 685 1936
rect 690 1933 693 1993
rect 690 1873 693 1926
rect 690 1826 693 1856
rect 698 1833 701 2156
rect 706 2083 709 2196
rect 690 1823 701 1826
rect 698 1812 701 1823
rect 690 1786 693 1796
rect 690 1783 701 1786
rect 682 1773 693 1776
rect 682 1733 685 1766
rect 674 1723 685 1726
rect 682 1703 685 1723
rect 690 1626 693 1773
rect 698 1693 701 1783
rect 698 1673 701 1686
rect 666 1623 693 1626
rect 666 1613 669 1623
rect 674 1606 677 1616
rect 634 1543 645 1546
rect 650 1593 661 1596
rect 626 1433 629 1446
rect 618 1403 629 1406
rect 618 1383 621 1396
rect 610 1353 621 1356
rect 610 763 613 1346
rect 618 1323 621 1353
rect 626 1343 629 1403
rect 626 1313 629 1336
rect 618 1173 621 1236
rect 618 1013 621 1146
rect 626 1123 629 1226
rect 634 1216 637 1543
rect 642 1443 645 1536
rect 650 1523 653 1593
rect 666 1586 669 1606
rect 674 1603 693 1606
rect 658 1583 669 1586
rect 666 1523 669 1536
rect 658 1446 661 1496
rect 654 1443 661 1446
rect 642 1413 645 1426
rect 654 1356 657 1443
rect 654 1353 661 1356
rect 642 1333 653 1336
rect 658 1326 661 1353
rect 650 1323 661 1326
rect 650 1256 653 1323
rect 642 1253 653 1256
rect 642 1233 645 1253
rect 666 1243 669 1436
rect 634 1213 641 1216
rect 650 1213 653 1226
rect 638 1146 641 1213
rect 634 1143 641 1146
rect 626 1103 629 1116
rect 634 1026 637 1143
rect 658 1133 661 1216
rect 666 1203 669 1236
rect 642 1123 661 1126
rect 642 1103 645 1123
rect 666 1113 669 1126
rect 674 1096 677 1546
rect 682 1523 685 1596
rect 690 1506 693 1603
rect 686 1503 693 1506
rect 686 1426 689 1503
rect 682 1423 689 1426
rect 682 1296 685 1423
rect 690 1393 693 1416
rect 690 1353 693 1386
rect 690 1313 693 1346
rect 682 1293 689 1296
rect 686 1196 689 1293
rect 626 1023 637 1026
rect 666 1093 677 1096
rect 682 1193 689 1196
rect 666 1026 669 1093
rect 682 1033 685 1193
rect 690 1123 693 1146
rect 690 1033 693 1106
rect 698 1083 701 1646
rect 706 1603 709 2056
rect 714 1963 717 2186
rect 722 2113 725 2206
rect 722 1993 725 2096
rect 706 1533 709 1556
rect 706 1403 709 1456
rect 706 1323 709 1336
rect 714 1306 717 1936
rect 722 1823 725 1896
rect 730 1813 733 2026
rect 738 2016 741 2156
rect 746 2093 749 2206
rect 754 2123 757 2216
rect 786 2186 789 2206
rect 802 2203 805 2216
rect 810 2213 813 2226
rect 818 2213 829 2216
rect 778 2183 789 2186
rect 818 2183 821 2213
rect 778 2136 781 2183
rect 778 2133 789 2136
rect 738 2013 749 2016
rect 722 1803 733 1806
rect 722 1686 725 1803
rect 738 1746 741 2006
rect 746 1826 749 2013
rect 754 1946 757 2116
rect 762 2096 765 2116
rect 762 2093 769 2096
rect 766 2026 769 2093
rect 762 2023 769 2026
rect 762 1953 765 2023
rect 754 1943 765 1946
rect 754 1903 757 1936
rect 746 1823 757 1826
rect 746 1773 749 1816
rect 738 1743 749 1746
rect 730 1703 733 1726
rect 738 1723 741 1736
rect 746 1723 749 1743
rect 722 1683 729 1686
rect 726 1586 729 1683
rect 722 1583 729 1586
rect 722 1543 725 1583
rect 730 1513 733 1566
rect 738 1543 741 1606
rect 746 1603 749 1616
rect 754 1546 757 1823
rect 762 1673 765 1943
rect 770 1806 773 2006
rect 778 1993 781 2066
rect 778 1813 781 1946
rect 786 1883 789 2133
rect 786 1833 789 1856
rect 794 1813 797 2146
rect 802 2073 805 2166
rect 810 2103 813 2126
rect 818 2036 821 2136
rect 826 2116 829 2126
rect 834 2123 837 2136
rect 842 2123 845 2243
rect 850 2226 853 2326
rect 858 2313 869 2316
rect 858 2243 861 2313
rect 874 2306 877 2326
rect 890 2323 893 2393
rect 914 2376 917 2416
rect 946 2413 949 2486
rect 970 2436 973 2676
rect 1050 2673 1053 2713
rect 978 2533 981 2556
rect 986 2543 989 2616
rect 1050 2613 1053 2626
rect 1002 2593 1005 2606
rect 1018 2523 1021 2546
rect 1082 2543 1085 2616
rect 1098 2586 1101 2773
rect 1106 2743 1109 2756
rect 1130 2703 1133 2746
rect 1138 2743 1141 2816
rect 1146 2803 1149 2903
rect 1098 2583 1105 2586
rect 1034 2456 1037 2536
rect 1102 2526 1105 2583
rect 1114 2573 1117 2616
rect 1138 2613 1141 2736
rect 1146 2623 1149 2736
rect 1154 2713 1157 2806
rect 1162 2776 1165 2886
rect 1194 2866 1197 3016
rect 1202 3003 1205 3046
rect 1210 2973 1213 3016
rect 1218 3003 1221 3016
rect 1234 3013 1245 3016
rect 1234 3003 1237 3013
rect 1250 3006 1253 3026
rect 1266 3013 1269 3036
rect 1274 3023 1277 3046
rect 1242 3003 1253 3006
rect 1234 2926 1237 2936
rect 1186 2863 1197 2866
rect 1186 2823 1189 2863
rect 1202 2836 1205 2926
rect 1226 2923 1237 2926
rect 1242 2923 1245 3003
rect 1266 2993 1269 3006
rect 1274 3003 1277 3016
rect 1250 2933 1253 2986
rect 1250 2923 1261 2926
rect 1274 2923 1277 2976
rect 1282 2923 1285 2936
rect 1298 2933 1301 3103
rect 1330 3073 1333 3116
rect 1338 3093 1341 3126
rect 1306 2993 1309 3006
rect 1322 2923 1325 3016
rect 1330 3003 1333 3026
rect 1346 3003 1349 3086
rect 1354 3073 1357 3126
rect 1374 3116 1377 3163
rect 1386 3123 1389 3326
rect 1374 3113 1381 3116
rect 1394 3113 1397 3216
rect 1354 2956 1357 3016
rect 1370 2973 1373 3016
rect 1378 3003 1381 3113
rect 1402 3096 1405 3256
rect 1410 3233 1421 3236
rect 1410 3213 1413 3233
rect 1418 3156 1421 3226
rect 1398 3093 1405 3096
rect 1410 3153 1421 3156
rect 1426 3153 1429 3316
rect 1474 3226 1477 3340
rect 1554 3313 1557 3340
rect 1514 3263 1541 3266
rect 1458 3223 1477 3226
rect 1506 3223 1509 3236
rect 1458 3183 1461 3223
rect 1474 3213 1509 3216
rect 1398 3026 1401 3093
rect 1398 3023 1405 3026
rect 1410 3023 1413 3153
rect 1418 3116 1421 3146
rect 1418 3113 1429 3116
rect 1426 3056 1429 3113
rect 1442 3083 1445 3136
rect 1450 3133 1453 3146
rect 1458 3123 1461 3166
rect 1466 3133 1469 3146
rect 1450 3103 1453 3116
rect 1474 3113 1477 3213
rect 1482 3163 1485 3206
rect 1482 3106 1485 3136
rect 1482 3103 1493 3106
rect 1418 3053 1429 3056
rect 1338 2953 1357 2956
rect 1226 2896 1229 2923
rect 1250 2916 1253 2923
rect 1234 2913 1253 2916
rect 1330 2913 1333 2936
rect 1226 2893 1237 2896
rect 1194 2833 1205 2836
rect 1170 2793 1173 2806
rect 1162 2773 1173 2776
rect 1170 2666 1173 2773
rect 1194 2766 1197 2833
rect 1234 2813 1237 2893
rect 1338 2823 1341 2953
rect 1346 2836 1349 2926
rect 1346 2833 1357 2836
rect 1210 2783 1213 2806
rect 1194 2763 1205 2766
rect 1202 2723 1205 2763
rect 1226 2733 1229 2756
rect 1290 2753 1293 2816
rect 1298 2803 1301 2816
rect 1322 2813 1341 2816
rect 1322 2743 1325 2813
rect 1338 2783 1341 2806
rect 1346 2803 1349 2826
rect 1354 2786 1357 2833
rect 1346 2783 1357 2786
rect 1362 2786 1365 2936
rect 1386 2903 1389 3016
rect 1394 2856 1397 3006
rect 1402 2906 1405 3023
rect 1418 3013 1421 3053
rect 1410 3003 1429 3006
rect 1434 3003 1437 3036
rect 1442 3023 1469 3026
rect 1410 2923 1413 3003
rect 1442 2993 1445 3016
rect 1466 3013 1469 3023
rect 1474 3003 1477 3066
rect 1490 3026 1493 3103
rect 1490 3023 1501 3026
rect 1482 2973 1485 3016
rect 1498 2986 1501 3023
rect 1506 2996 1509 3206
rect 1514 3203 1517 3263
rect 1538 3216 1541 3263
rect 1538 3213 1549 3216
rect 1554 3213 1557 3226
rect 1538 3116 1541 3136
rect 1554 3133 1557 3206
rect 1562 3163 1565 3236
rect 1586 3233 1613 3236
rect 1586 3213 1589 3233
rect 1578 3173 1581 3206
rect 1594 3183 1597 3216
rect 1618 3166 1621 3316
rect 1610 3163 1621 3166
rect 1562 3143 1589 3146
rect 1530 3113 1541 3116
rect 1546 3113 1549 3126
rect 1530 3066 1533 3113
rect 1554 3093 1557 3126
rect 1530 3063 1541 3066
rect 1514 3013 1525 3016
rect 1530 3013 1533 3046
rect 1538 3033 1541 3063
rect 1546 3026 1549 3046
rect 1562 3036 1565 3143
rect 1570 3133 1581 3136
rect 1586 3133 1589 3143
rect 1570 3103 1573 3126
rect 1538 3023 1549 3026
rect 1554 3033 1565 3036
rect 1538 3003 1541 3023
rect 1554 3006 1557 3033
rect 1546 3003 1557 3006
rect 1546 2996 1549 3003
rect 1506 2993 1549 2996
rect 1498 2983 1509 2986
rect 1506 2966 1509 2983
rect 1442 2913 1445 2926
rect 1450 2923 1453 2936
rect 1402 2903 1409 2906
rect 1386 2853 1397 2856
rect 1386 2813 1389 2853
rect 1406 2846 1409 2903
rect 1406 2843 1421 2846
rect 1386 2786 1389 2806
rect 1362 2783 1389 2786
rect 1410 2783 1413 2816
rect 1346 2743 1349 2783
rect 1418 2776 1421 2843
rect 1402 2773 1421 2776
rect 1402 2756 1405 2773
rect 1394 2753 1405 2756
rect 1410 2763 1453 2766
rect 1162 2663 1173 2666
rect 1162 2646 1165 2663
rect 1158 2643 1165 2646
rect 1158 2576 1161 2643
rect 1158 2573 1165 2576
rect 1114 2533 1125 2536
rect 962 2433 973 2436
rect 1018 2453 1037 2456
rect 914 2373 925 2376
rect 866 2303 877 2306
rect 850 2223 857 2226
rect 854 2156 857 2223
rect 866 2213 869 2303
rect 866 2163 869 2206
rect 854 2153 861 2156
rect 850 2123 853 2136
rect 858 2123 861 2153
rect 826 2113 869 2116
rect 850 2083 853 2106
rect 874 2096 877 2236
rect 866 2093 877 2096
rect 810 2033 821 2036
rect 826 2026 829 2056
rect 866 2026 869 2093
rect 818 2023 829 2026
rect 858 2023 869 2026
rect 802 2003 805 2016
rect 802 1943 805 1956
rect 802 1923 805 1936
rect 770 1803 781 1806
rect 770 1733 773 1796
rect 770 1656 773 1696
rect 778 1663 781 1803
rect 786 1723 789 1736
rect 770 1653 781 1656
rect 762 1583 765 1616
rect 778 1603 781 1653
rect 786 1583 789 1596
rect 794 1576 797 1806
rect 802 1723 805 1876
rect 810 1863 813 1936
rect 818 1923 821 2023
rect 826 1913 829 1926
rect 802 1703 805 1716
rect 802 1603 805 1616
rect 778 1573 797 1576
rect 754 1543 761 1546
rect 738 1466 741 1516
rect 730 1463 741 1466
rect 746 1446 749 1536
rect 758 1446 761 1543
rect 722 1443 749 1446
rect 754 1443 761 1446
rect 722 1373 725 1443
rect 730 1426 733 1436
rect 738 1433 749 1436
rect 730 1423 749 1426
rect 730 1406 733 1416
rect 754 1406 757 1443
rect 770 1426 773 1526
rect 778 1503 781 1573
rect 786 1526 789 1546
rect 786 1523 793 1526
rect 802 1523 805 1576
rect 730 1403 741 1406
rect 730 1333 733 1396
rect 738 1343 741 1403
rect 750 1403 757 1406
rect 762 1423 773 1426
rect 722 1313 725 1326
rect 706 1293 709 1306
rect 714 1303 725 1306
rect 730 1303 733 1326
rect 706 1076 709 1206
rect 714 1156 717 1246
rect 722 1203 725 1303
rect 738 1213 741 1336
rect 750 1246 753 1403
rect 746 1243 753 1246
rect 746 1196 749 1243
rect 730 1193 749 1196
rect 714 1153 725 1156
rect 714 1123 717 1136
rect 698 1073 709 1076
rect 698 1026 701 1073
rect 722 1066 725 1153
rect 730 1093 733 1193
rect 738 1133 749 1136
rect 746 1086 749 1126
rect 754 1113 757 1236
rect 746 1083 757 1086
rect 666 1023 677 1026
rect 618 933 621 956
rect 618 756 621 866
rect 610 753 621 756
rect 626 753 629 1023
rect 650 973 653 1006
rect 666 926 669 936
rect 642 923 669 926
rect 634 893 637 916
rect 642 913 661 916
rect 666 913 669 923
rect 642 903 645 913
rect 650 856 653 906
rect 642 853 653 856
rect 642 833 645 853
rect 650 823 653 846
rect 658 816 661 826
rect 650 813 661 816
rect 610 683 613 753
rect 618 723 621 746
rect 626 646 629 736
rect 634 723 637 806
rect 642 703 645 726
rect 650 713 653 813
rect 658 726 661 806
rect 666 793 669 826
rect 666 733 669 776
rect 658 723 669 726
rect 610 643 629 646
rect 594 593 597 606
rect 570 533 577 536
rect 574 466 577 533
rect 602 473 605 536
rect 554 433 565 436
rect 570 463 577 466
rect 538 363 549 366
rect 538 333 541 346
rect 546 326 549 363
rect 514 313 525 316
rect 530 313 533 326
rect 538 323 549 326
rect 554 316 557 433
rect 562 413 565 426
rect 570 406 573 463
rect 578 413 581 446
rect 610 443 613 643
rect 618 556 621 606
rect 626 593 629 616
rect 642 613 645 626
rect 650 603 653 686
rect 618 553 629 556
rect 594 406 597 436
rect 602 413 605 426
rect 562 386 565 406
rect 570 403 581 406
rect 586 403 597 406
rect 562 383 569 386
rect 546 313 557 316
rect 498 293 509 296
rect 498 223 501 293
rect 514 223 517 313
rect 546 296 549 313
rect 566 306 569 383
rect 538 293 549 296
rect 562 303 569 306
rect 394 206 397 216
rect 394 203 421 206
rect 338 113 341 126
rect 354 106 357 126
rect 314 103 357 106
rect 410 93 413 136
rect 418 123 421 203
rect 426 133 429 216
rect 434 123 437 206
rect 458 193 461 216
rect 498 163 501 206
rect 538 176 541 293
rect 562 233 565 303
rect 578 253 581 403
rect 610 376 613 406
rect 538 173 549 176
rect 546 153 549 173
rect 418 113 429 116
rect 498 103 501 126
rect 506 123 509 146
rect 514 143 549 146
rect 514 133 517 143
rect 522 93 525 126
rect 538 113 541 126
rect 546 123 549 143
rect 554 133 557 226
rect 562 213 565 226
rect 570 193 573 206
rect 562 133 565 156
rect 586 113 589 376
rect 606 373 613 376
rect 594 293 597 316
rect 606 286 609 373
rect 618 296 621 546
rect 626 496 629 553
rect 634 513 637 526
rect 642 513 653 516
rect 626 493 633 496
rect 630 336 633 493
rect 626 333 633 336
rect 642 333 645 513
rect 658 443 661 666
rect 666 533 669 723
rect 674 706 677 1023
rect 682 1016 685 1026
rect 690 1023 701 1026
rect 706 1063 725 1066
rect 706 1023 709 1063
rect 714 1016 717 1026
rect 682 1013 717 1016
rect 730 1013 733 1076
rect 682 783 685 836
rect 682 733 685 746
rect 682 713 685 726
rect 674 703 685 706
rect 682 633 685 703
rect 674 596 677 626
rect 690 603 693 986
rect 706 923 709 1006
rect 730 933 733 946
rect 706 913 725 916
rect 706 903 709 913
rect 730 906 733 926
rect 714 903 733 906
rect 738 853 741 1006
rect 706 803 709 836
rect 698 653 701 786
rect 674 593 693 596
rect 674 533 685 536
rect 690 533 693 593
rect 698 563 701 636
rect 706 616 709 766
rect 730 743 733 766
rect 714 623 717 736
rect 730 703 733 726
rect 706 613 717 616
rect 722 613 725 696
rect 738 686 741 806
rect 746 776 749 1036
rect 754 1003 757 1083
rect 754 893 757 996
rect 754 793 757 856
rect 746 773 753 776
rect 750 706 753 773
rect 762 733 765 1423
rect 770 1393 773 1416
rect 770 1213 773 1386
rect 770 1103 773 1126
rect 770 803 773 1076
rect 778 973 781 1466
rect 790 1446 793 1523
rect 810 1493 813 1816
rect 818 1813 821 1856
rect 834 1823 837 1956
rect 842 1933 845 1986
rect 850 1916 853 2006
rect 858 1943 861 2023
rect 866 2013 877 2016
rect 846 1913 853 1916
rect 846 1826 849 1913
rect 846 1823 853 1826
rect 818 1693 821 1786
rect 834 1756 837 1816
rect 850 1803 853 1823
rect 858 1813 861 1926
rect 858 1783 861 1806
rect 826 1753 837 1756
rect 826 1616 829 1753
rect 834 1733 837 1746
rect 842 1743 853 1746
rect 834 1633 837 1726
rect 826 1613 833 1616
rect 818 1593 821 1606
rect 818 1533 821 1566
rect 818 1503 821 1516
rect 830 1486 833 1613
rect 826 1483 833 1486
rect 826 1463 829 1483
rect 786 1443 793 1446
rect 786 1126 789 1443
rect 794 1403 797 1426
rect 794 1256 797 1336
rect 802 1273 805 1446
rect 810 1433 829 1436
rect 810 1323 813 1433
rect 818 1416 821 1426
rect 826 1423 829 1433
rect 842 1426 845 1736
rect 858 1616 861 1736
rect 866 1703 869 1866
rect 874 1786 877 1946
rect 882 1913 885 2146
rect 890 2126 893 2226
rect 898 2183 901 2216
rect 914 2193 917 2356
rect 922 2333 925 2373
rect 930 2333 933 2346
rect 954 2303 957 2316
rect 962 2313 965 2433
rect 978 2373 981 2406
rect 1002 2376 1005 2416
rect 1018 2396 1021 2453
rect 1058 2413 1061 2496
rect 1082 2406 1085 2526
rect 1102 2523 1109 2526
rect 1106 2413 1109 2523
rect 1138 2503 1141 2526
rect 1122 2413 1125 2426
rect 1146 2423 1149 2526
rect 1162 2513 1165 2573
rect 1170 2493 1173 2536
rect 1194 2533 1197 2616
rect 1202 2586 1205 2616
rect 1250 2613 1253 2736
rect 1346 2733 1357 2736
rect 1322 2723 1341 2726
rect 1338 2713 1341 2723
rect 1298 2616 1301 2636
rect 1290 2613 1301 2616
rect 1218 2593 1221 2606
rect 1202 2583 1213 2586
rect 1210 2533 1213 2583
rect 1186 2503 1189 2526
rect 1202 2523 1221 2526
rect 1242 2523 1245 2566
rect 1290 2556 1293 2613
rect 1306 2563 1309 2616
rect 1354 2613 1357 2733
rect 1362 2713 1365 2726
rect 1394 2706 1397 2753
rect 1410 2733 1413 2763
rect 1394 2703 1405 2706
rect 1402 2633 1405 2703
rect 1330 2593 1333 2606
rect 1290 2553 1297 2556
rect 1250 2533 1253 2546
rect 1202 2446 1205 2523
rect 1266 2503 1269 2536
rect 1198 2443 1205 2446
rect 1018 2393 1029 2396
rect 986 2373 1005 2376
rect 1026 2373 1029 2393
rect 978 2326 981 2366
rect 986 2333 989 2373
rect 978 2323 989 2326
rect 986 2313 989 2323
rect 922 2223 933 2226
rect 922 2203 925 2223
rect 930 2213 949 2216
rect 930 2146 933 2213
rect 938 2193 941 2206
rect 954 2203 957 2226
rect 962 2196 965 2296
rect 946 2193 965 2196
rect 922 2143 933 2146
rect 938 2143 941 2156
rect 922 2126 925 2143
rect 930 2133 941 2136
rect 890 2123 909 2126
rect 890 2013 893 2096
rect 890 1983 893 2006
rect 898 2003 901 2116
rect 906 2093 909 2123
rect 918 2123 925 2126
rect 906 1996 909 2086
rect 918 2046 921 2123
rect 914 2043 921 2046
rect 914 2006 917 2043
rect 922 2013 925 2036
rect 914 2003 925 2006
rect 890 1943 893 1976
rect 898 1953 901 1996
rect 906 1993 917 1996
rect 914 1936 917 1993
rect 898 1933 917 1936
rect 898 1863 901 1926
rect 906 1923 917 1926
rect 882 1793 885 1826
rect 906 1823 909 1923
rect 922 1913 925 2003
rect 930 1983 933 2126
rect 946 2116 949 2193
rect 954 2133 957 2146
rect 946 2113 953 2116
rect 938 1993 941 2096
rect 950 2046 953 2113
rect 962 2056 965 2186
rect 970 2143 973 2216
rect 978 2186 981 2236
rect 994 2223 997 2336
rect 1002 2216 1005 2326
rect 1010 2296 1013 2316
rect 1010 2293 1021 2296
rect 1018 2226 1021 2293
rect 994 2213 1005 2216
rect 1010 2223 1021 2226
rect 994 2193 997 2213
rect 1002 2186 1005 2206
rect 978 2183 1005 2186
rect 978 2133 981 2176
rect 1002 2156 1005 2176
rect 994 2153 1005 2156
rect 994 2086 997 2153
rect 994 2083 1005 2086
rect 962 2053 981 2056
rect 946 2043 953 2046
rect 922 1846 925 1886
rect 930 1853 933 1936
rect 938 1923 941 1966
rect 938 1893 941 1916
rect 922 1843 933 1846
rect 890 1813 909 1816
rect 890 1786 893 1813
rect 874 1783 893 1786
rect 874 1723 877 1776
rect 890 1723 893 1746
rect 898 1716 901 1806
rect 890 1713 901 1716
rect 850 1613 861 1616
rect 850 1566 853 1613
rect 858 1586 861 1606
rect 866 1593 869 1616
rect 882 1603 885 1676
rect 890 1613 893 1713
rect 906 1696 909 1813
rect 914 1793 917 1836
rect 922 1803 925 1826
rect 930 1813 933 1843
rect 938 1836 941 1876
rect 946 1853 949 2043
rect 954 2006 957 2026
rect 962 2013 965 2036
rect 970 2013 973 2046
rect 978 2023 981 2053
rect 954 2003 965 2006
rect 954 1946 957 1996
rect 962 1953 965 2003
rect 954 1943 973 1946
rect 938 1833 949 1836
rect 946 1813 949 1833
rect 954 1796 957 1816
rect 946 1793 957 1796
rect 902 1693 909 1696
rect 902 1636 905 1693
rect 902 1633 909 1636
rect 890 1586 893 1606
rect 858 1583 893 1586
rect 890 1573 893 1583
rect 850 1563 861 1566
rect 850 1513 853 1526
rect 842 1423 849 1426
rect 818 1413 829 1416
rect 818 1363 821 1406
rect 826 1313 829 1413
rect 834 1393 837 1416
rect 834 1343 837 1376
rect 846 1346 849 1423
rect 842 1343 849 1346
rect 834 1306 837 1336
rect 818 1303 837 1306
rect 794 1253 829 1256
rect 794 1223 797 1253
rect 794 1183 797 1216
rect 802 1153 805 1236
rect 810 1223 813 1236
rect 786 1123 797 1126
rect 778 933 781 956
rect 786 926 789 1116
rect 782 923 789 926
rect 782 846 785 923
rect 778 843 785 846
rect 734 683 741 686
rect 746 703 753 706
rect 770 703 773 726
rect 746 683 749 703
rect 666 506 669 526
rect 682 513 685 526
rect 698 506 701 516
rect 666 503 701 506
rect 706 486 709 606
rect 626 313 629 333
rect 658 326 661 336
rect 642 323 661 326
rect 618 293 629 296
rect 606 283 613 286
rect 594 203 597 226
rect 610 213 613 283
rect 626 226 629 293
rect 618 223 629 226
rect 618 206 621 223
rect 618 203 637 206
rect 642 203 645 323
rect 650 313 661 316
rect 666 313 669 406
rect 674 343 677 416
rect 682 376 685 486
rect 702 483 709 486
rect 690 383 693 416
rect 702 396 705 483
rect 702 393 709 396
rect 682 373 693 376
rect 706 373 709 393
rect 714 376 717 613
rect 722 493 725 586
rect 734 576 737 683
rect 762 676 765 686
rect 746 673 765 676
rect 746 603 749 673
rect 730 573 737 576
rect 730 513 733 573
rect 754 566 757 626
rect 778 576 781 843
rect 794 833 797 1123
rect 810 1013 813 1216
rect 802 993 805 1006
rect 802 923 805 946
rect 810 913 813 1006
rect 818 833 821 1246
rect 826 1146 829 1253
rect 834 1163 837 1226
rect 826 1143 833 1146
rect 830 966 833 1143
rect 826 963 833 966
rect 826 943 829 963
rect 826 833 829 936
rect 834 903 837 916
rect 842 866 845 1343
rect 858 1336 861 1563
rect 898 1546 901 1616
rect 906 1583 909 1633
rect 914 1623 917 1766
rect 922 1716 925 1786
rect 930 1723 933 1776
rect 946 1763 949 1793
rect 954 1746 957 1786
rect 938 1743 957 1746
rect 938 1733 941 1743
rect 938 1723 949 1726
rect 954 1723 957 1736
rect 962 1723 965 1886
rect 922 1713 933 1716
rect 922 1603 925 1626
rect 866 1543 901 1546
rect 866 1446 869 1543
rect 874 1493 877 1526
rect 890 1513 893 1536
rect 898 1506 901 1536
rect 906 1533 909 1546
rect 882 1503 901 1506
rect 922 1483 925 1546
rect 874 1446 877 1456
rect 866 1443 877 1446
rect 866 1423 869 1436
rect 858 1333 865 1336
rect 850 1313 853 1326
rect 850 1153 853 1296
rect 862 1256 865 1333
rect 858 1253 865 1256
rect 858 1233 861 1253
rect 866 1183 869 1216
rect 858 1133 861 1156
rect 850 1113 853 1126
rect 850 953 853 1016
rect 850 913 853 946
rect 858 933 861 1006
rect 866 993 869 1166
rect 874 1156 877 1443
rect 882 1386 885 1446
rect 890 1403 893 1416
rect 914 1413 917 1426
rect 922 1413 925 1436
rect 898 1403 909 1406
rect 930 1403 933 1713
rect 970 1706 973 1943
rect 986 1926 989 2026
rect 994 1993 997 2066
rect 1002 2043 1005 2083
rect 1002 2003 1005 2016
rect 994 1933 997 1966
rect 978 1903 981 1926
rect 986 1923 997 1926
rect 986 1903 989 1916
rect 978 1723 981 1856
rect 986 1793 989 1806
rect 994 1786 997 1923
rect 1002 1813 1005 1986
rect 1010 1896 1013 2223
rect 1018 2133 1021 2196
rect 1026 2173 1029 2206
rect 1018 2013 1021 2126
rect 1026 1956 1029 2126
rect 1034 2003 1037 2356
rect 1066 2343 1069 2406
rect 1082 2403 1125 2406
rect 1162 2393 1165 2406
rect 1198 2386 1201 2443
rect 1294 2436 1297 2553
rect 1294 2433 1301 2436
rect 1210 2393 1213 2416
rect 1242 2413 1245 2426
rect 1198 2383 1205 2386
rect 1082 2333 1085 2366
rect 1082 2316 1085 2326
rect 1090 2323 1093 2346
rect 1106 2323 1109 2336
rect 1114 2316 1117 2336
rect 1162 2333 1165 2346
rect 1146 2323 1165 2326
rect 1082 2313 1117 2316
rect 1090 2296 1093 2313
rect 1082 2293 1093 2296
rect 1066 2226 1069 2236
rect 1042 2223 1069 2226
rect 1082 2226 1085 2293
rect 1082 2223 1093 2226
rect 1042 2213 1045 2223
rect 1050 2203 1053 2216
rect 1042 2123 1045 2136
rect 1050 2123 1061 2126
rect 1066 2123 1069 2196
rect 1074 2133 1077 2156
rect 1082 2123 1085 2206
rect 1018 1953 1029 1956
rect 1018 1913 1021 1953
rect 1010 1893 1017 1896
rect 1014 1826 1017 1893
rect 1026 1873 1029 1946
rect 1034 1923 1037 1986
rect 1042 1933 1045 2116
rect 1050 1983 1053 2076
rect 1058 2053 1085 2056
rect 1042 1913 1045 1926
rect 1010 1823 1017 1826
rect 986 1783 997 1786
rect 962 1703 973 1706
rect 962 1636 965 1703
rect 962 1633 973 1636
rect 946 1603 957 1606
rect 938 1526 941 1596
rect 946 1543 949 1603
rect 938 1523 945 1526
rect 882 1383 889 1386
rect 886 1246 889 1383
rect 882 1243 889 1246
rect 882 1223 885 1243
rect 898 1226 901 1336
rect 906 1323 909 1403
rect 922 1383 925 1396
rect 942 1376 945 1523
rect 938 1373 945 1376
rect 894 1223 901 1226
rect 894 1156 897 1223
rect 874 1153 885 1156
rect 894 1153 901 1156
rect 874 1123 877 1146
rect 882 1106 885 1153
rect 878 1103 885 1106
rect 878 1036 881 1103
rect 890 1083 893 1126
rect 898 1066 901 1153
rect 906 1073 909 1256
rect 898 1063 909 1066
rect 878 1033 885 1036
rect 874 993 877 1016
rect 882 986 885 1033
rect 890 1013 893 1056
rect 898 1003 901 1016
rect 874 983 885 986
rect 834 863 845 866
rect 850 853 853 906
rect 858 893 861 926
rect 866 903 869 956
rect 786 783 789 826
rect 842 823 845 846
rect 786 723 789 736
rect 794 706 797 726
rect 790 703 797 706
rect 790 626 793 703
rect 790 623 797 626
rect 786 593 789 606
rect 794 596 797 623
rect 802 613 805 816
rect 826 796 829 816
rect 826 793 837 796
rect 810 733 813 766
rect 826 733 829 746
rect 810 723 821 726
rect 826 723 837 726
rect 810 663 813 723
rect 842 676 845 766
rect 850 753 853 816
rect 858 736 861 836
rect 866 803 869 846
rect 834 673 845 676
rect 854 733 861 736
rect 810 613 813 636
rect 794 593 805 596
rect 778 573 785 576
rect 754 563 773 566
rect 738 523 741 556
rect 754 546 757 563
rect 746 543 757 546
rect 746 516 749 543
rect 738 513 749 516
rect 738 496 741 513
rect 754 496 757 536
rect 770 533 773 563
rect 762 513 765 526
rect 738 493 745 496
rect 754 493 769 496
rect 714 373 725 376
rect 690 333 693 373
rect 698 363 717 366
rect 690 303 693 316
rect 698 276 701 346
rect 698 273 709 276
rect 666 213 677 216
rect 666 203 669 213
rect 674 196 677 206
rect 682 203 685 226
rect 690 196 693 216
rect 706 213 709 273
rect 674 193 693 196
rect 666 123 669 186
rect 698 163 701 206
rect 706 193 709 206
rect 714 133 717 363
rect 722 203 725 373
rect 730 306 733 446
rect 742 426 745 493
rect 742 423 749 426
rect 746 403 749 423
rect 754 413 757 486
rect 766 426 769 493
rect 782 486 785 573
rect 802 526 805 593
rect 778 483 785 486
rect 766 423 773 426
rect 770 403 773 423
rect 770 333 773 366
rect 730 303 741 306
rect 738 216 741 303
rect 770 273 773 326
rect 770 223 773 266
rect 730 213 741 216
rect 778 213 781 483
rect 794 426 797 526
rect 802 523 809 526
rect 786 423 797 426
rect 806 426 809 523
rect 818 446 821 586
rect 826 463 829 606
rect 834 533 837 673
rect 854 666 857 733
rect 854 663 861 666
rect 842 593 845 606
rect 850 586 853 646
rect 858 603 861 663
rect 842 583 853 586
rect 834 493 837 526
rect 842 523 845 583
rect 850 533 853 566
rect 850 523 861 526
rect 850 483 853 523
rect 818 443 829 446
rect 806 423 813 426
rect 786 353 789 423
rect 786 223 789 326
rect 794 273 797 416
rect 802 316 805 406
rect 810 393 813 423
rect 818 413 821 436
rect 826 423 829 443
rect 810 343 821 346
rect 810 333 813 343
rect 826 333 829 366
rect 834 343 837 356
rect 802 313 813 316
rect 794 216 797 256
rect 810 246 813 313
rect 834 263 837 316
rect 842 303 845 426
rect 850 386 853 426
rect 858 403 861 466
rect 850 383 857 386
rect 854 316 857 383
rect 866 333 869 726
rect 874 613 877 983
rect 882 786 885 966
rect 890 933 893 956
rect 898 943 901 996
rect 890 903 893 916
rect 898 823 901 926
rect 890 803 901 806
rect 882 783 889 786
rect 886 636 889 783
rect 898 723 901 746
rect 906 743 909 1063
rect 914 993 917 1276
rect 922 1153 925 1356
rect 914 803 917 976
rect 922 796 925 1146
rect 930 1113 933 1326
rect 938 1243 941 1373
rect 954 1343 957 1596
rect 962 1463 965 1616
rect 970 1516 973 1633
rect 978 1623 981 1636
rect 978 1603 981 1616
rect 978 1533 981 1576
rect 986 1523 989 1783
rect 994 1733 1005 1736
rect 994 1603 997 1696
rect 1010 1616 1013 1823
rect 1018 1723 1021 1806
rect 1018 1693 1021 1716
rect 1026 1673 1029 1736
rect 1034 1646 1037 1836
rect 1042 1813 1045 1856
rect 1050 1803 1053 1976
rect 1058 1796 1061 2053
rect 1074 2016 1077 2046
rect 1082 2023 1085 2053
rect 1066 1983 1069 2016
rect 1074 2013 1085 2016
rect 1090 2013 1093 2223
rect 1098 2186 1101 2276
rect 1114 2243 1117 2306
rect 1170 2286 1173 2336
rect 1202 2326 1205 2383
rect 1258 2333 1261 2346
rect 1202 2323 1209 2326
rect 1154 2283 1173 2286
rect 1114 2223 1117 2236
rect 1106 2203 1117 2206
rect 1122 2196 1125 2276
rect 1114 2193 1125 2196
rect 1098 2183 1105 2186
rect 1102 2036 1105 2183
rect 1114 2143 1117 2193
rect 1130 2186 1133 2266
rect 1138 2213 1141 2226
rect 1130 2183 1141 2186
rect 1098 2033 1105 2036
rect 1114 2036 1117 2046
rect 1122 2043 1125 2176
rect 1138 2166 1141 2183
rect 1146 2173 1149 2246
rect 1154 2203 1157 2283
rect 1162 2223 1165 2236
rect 1170 2213 1173 2266
rect 1162 2166 1165 2206
rect 1170 2193 1173 2206
rect 1138 2163 1149 2166
rect 1130 2133 1133 2156
rect 1114 2033 1125 2036
rect 1082 2003 1085 2013
rect 1098 1966 1101 2033
rect 1114 2016 1117 2026
rect 1106 2013 1117 2016
rect 1106 1983 1109 2013
rect 1114 1996 1117 2006
rect 1122 2003 1125 2033
rect 1130 1996 1133 2116
rect 1138 2043 1141 2126
rect 1146 2086 1149 2163
rect 1154 2163 1165 2166
rect 1154 2153 1157 2163
rect 1162 2153 1173 2156
rect 1154 2133 1157 2146
rect 1154 2093 1157 2126
rect 1162 2113 1165 2153
rect 1170 2086 1173 2126
rect 1146 2083 1173 2086
rect 1146 2056 1149 2076
rect 1146 2053 1153 2056
rect 1114 1993 1133 1996
rect 1098 1963 1109 1966
rect 1066 1883 1069 1936
rect 1082 1883 1085 1926
rect 1066 1813 1069 1826
rect 1050 1793 1061 1796
rect 1066 1803 1077 1806
rect 1050 1706 1053 1793
rect 1066 1723 1069 1803
rect 1082 1793 1085 1816
rect 1074 1733 1085 1736
rect 1026 1643 1037 1646
rect 1042 1703 1053 1706
rect 1010 1613 1017 1616
rect 1002 1593 1005 1606
rect 970 1513 977 1516
rect 974 1446 977 1513
rect 970 1443 977 1446
rect 946 1293 949 1336
rect 962 1333 965 1426
rect 970 1373 973 1443
rect 978 1413 981 1426
rect 978 1393 981 1406
rect 954 1213 957 1326
rect 962 1323 973 1326
rect 970 1303 973 1323
rect 978 1296 981 1336
rect 966 1293 981 1296
rect 966 1226 969 1293
rect 978 1273 981 1293
rect 962 1223 969 1226
rect 962 1206 965 1223
rect 986 1206 989 1466
rect 946 1163 949 1206
rect 954 1203 965 1206
rect 954 1146 957 1156
rect 938 1143 957 1146
rect 914 793 925 796
rect 914 656 917 793
rect 922 723 925 746
rect 930 666 933 1086
rect 938 993 941 1006
rect 946 983 949 1143
rect 954 1103 957 1136
rect 962 1036 965 1186
rect 970 1123 973 1206
rect 978 1203 989 1206
rect 978 1143 981 1203
rect 994 1196 997 1546
rect 1002 1533 1005 1586
rect 1002 1423 1005 1526
rect 1014 1456 1017 1613
rect 1026 1596 1029 1643
rect 1034 1623 1037 1636
rect 1034 1603 1037 1616
rect 1026 1593 1037 1596
rect 1026 1483 1029 1546
rect 1034 1473 1037 1593
rect 1042 1566 1045 1703
rect 1074 1676 1077 1733
rect 1082 1703 1085 1726
rect 1074 1673 1085 1676
rect 1050 1613 1053 1626
rect 1066 1613 1069 1636
rect 1042 1563 1061 1566
rect 1042 1463 1045 1536
rect 1010 1453 1017 1456
rect 1002 1403 1005 1416
rect 1002 1253 1005 1366
rect 1010 1306 1013 1453
rect 1018 1403 1021 1436
rect 1050 1433 1053 1526
rect 1058 1426 1061 1563
rect 1066 1496 1069 1556
rect 1074 1513 1077 1646
rect 1066 1493 1073 1496
rect 1050 1423 1061 1426
rect 1070 1426 1073 1493
rect 1070 1423 1077 1426
rect 1018 1326 1021 1346
rect 1026 1333 1029 1416
rect 1042 1396 1045 1416
rect 1050 1403 1053 1423
rect 1058 1403 1061 1416
rect 1066 1396 1069 1416
rect 1042 1393 1069 1396
rect 1034 1333 1037 1386
rect 1066 1333 1069 1386
rect 1018 1323 1029 1326
rect 1010 1303 1017 1306
rect 1014 1246 1017 1303
rect 1010 1243 1017 1246
rect 986 1046 989 1196
rect 994 1193 1005 1196
rect 994 1123 997 1193
rect 1002 1053 1005 1136
rect 986 1043 997 1046
rect 958 1033 965 1036
rect 958 986 961 1033
rect 970 1013 973 1026
rect 978 1013 989 1016
rect 958 983 965 986
rect 962 963 965 983
rect 938 843 941 946
rect 946 943 981 946
rect 946 883 949 943
rect 954 903 957 936
rect 978 933 981 943
rect 986 926 989 1006
rect 962 923 989 926
rect 986 896 989 916
rect 978 893 989 896
rect 954 813 957 856
rect 978 846 981 893
rect 978 843 989 846
rect 938 733 941 786
rect 954 733 965 736
rect 938 716 941 726
rect 946 723 965 726
rect 938 713 965 716
rect 970 696 973 806
rect 978 763 981 826
rect 986 803 989 843
rect 994 726 997 1043
rect 1002 913 1005 966
rect 1002 803 1005 846
rect 1010 813 1013 1243
rect 1018 1163 1021 1196
rect 1018 1113 1021 1126
rect 1026 1116 1029 1323
rect 1042 1246 1045 1326
rect 1074 1293 1077 1423
rect 1082 1383 1085 1673
rect 1090 1533 1093 1926
rect 1098 1923 1101 1956
rect 1106 1916 1109 1963
rect 1114 1933 1117 1993
rect 1106 1913 1113 1916
rect 1098 1833 1101 1896
rect 1110 1846 1113 1913
rect 1106 1843 1113 1846
rect 1098 1703 1101 1766
rect 1106 1696 1109 1843
rect 1114 1763 1117 1826
rect 1122 1756 1125 1936
rect 1130 1833 1133 1926
rect 1138 1896 1141 2026
rect 1150 1976 1153 2053
rect 1162 2036 1165 2046
rect 1178 2043 1181 2216
rect 1186 2073 1189 2256
rect 1194 2123 1197 2316
rect 1206 2206 1209 2323
rect 1266 2316 1269 2416
rect 1290 2403 1293 2416
rect 1298 2413 1301 2433
rect 1306 2406 1309 2526
rect 1354 2523 1357 2606
rect 1426 2593 1429 2736
rect 1450 2723 1453 2763
rect 1458 2743 1461 2966
rect 1506 2963 1517 2966
rect 1466 2913 1469 2956
rect 1482 2923 1485 2936
rect 1514 2896 1517 2963
rect 1562 2936 1565 3026
rect 1570 3013 1573 3066
rect 1578 3046 1581 3133
rect 1586 3113 1589 3126
rect 1610 3076 1613 3163
rect 1610 3073 1621 3076
rect 1578 3043 1597 3046
rect 1586 3003 1589 3016
rect 1594 3003 1597 3043
rect 1618 3013 1621 3073
rect 1626 3043 1629 3126
rect 1634 3073 1637 3340
rect 1650 3323 1653 3340
rect 1858 3326 1861 3340
rect 1650 3223 1653 3246
rect 1650 3203 1653 3216
rect 1666 3206 1669 3226
rect 1666 3203 1677 3206
rect 1682 3156 1685 3216
rect 1690 3213 1693 3246
rect 1754 3223 1757 3236
rect 1770 3226 1773 3256
rect 1802 3246 1805 3326
rect 1850 3323 1861 3326
rect 1802 3243 1809 3246
rect 1778 3233 1797 3236
rect 1770 3223 1781 3226
rect 1690 3193 1693 3206
rect 1706 3176 1709 3196
rect 1746 3186 1749 3216
rect 1762 3213 1773 3216
rect 1698 3173 1709 3176
rect 1738 3183 1749 3186
rect 1754 3183 1757 3206
rect 1674 3146 1677 3156
rect 1682 3153 1693 3156
rect 1642 3133 1645 3146
rect 1674 3143 1685 3146
rect 1650 3133 1661 3136
rect 1642 3123 1653 3126
rect 1666 3106 1669 3136
rect 1682 3133 1685 3143
rect 1674 3123 1685 3126
rect 1690 3123 1693 3153
rect 1738 3133 1741 3183
rect 1746 3143 1757 3146
rect 1778 3136 1781 3223
rect 1786 3213 1789 3226
rect 1794 3203 1797 3233
rect 1786 3193 1797 3196
rect 1806 3186 1809 3243
rect 1850 3216 1853 3323
rect 1802 3183 1809 3186
rect 1746 3133 1757 3136
rect 1778 3133 1785 3136
rect 1746 3126 1749 3133
rect 1730 3123 1749 3126
rect 1650 3103 1669 3106
rect 1626 3013 1629 3026
rect 1530 2923 1533 2936
rect 1554 2933 1565 2936
rect 1570 2936 1573 2946
rect 1570 2933 1597 2936
rect 1602 2933 1613 2936
rect 1554 2916 1557 2933
rect 1506 2893 1517 2896
rect 1550 2913 1557 2916
rect 1466 2813 1469 2826
rect 1498 2803 1501 2816
rect 1506 2746 1509 2893
rect 1550 2856 1553 2913
rect 1550 2853 1557 2856
rect 1514 2753 1517 2816
rect 1530 2793 1533 2806
rect 1506 2743 1517 2746
rect 1514 2726 1517 2743
rect 1506 2723 1517 2726
rect 1506 2636 1509 2723
rect 1434 2613 1437 2626
rect 1442 2603 1445 2616
rect 1458 2613 1461 2636
rect 1506 2633 1517 2636
rect 1474 2613 1477 2626
rect 1450 2593 1453 2606
rect 1314 2416 1317 2516
rect 1370 2503 1373 2536
rect 1410 2506 1413 2526
rect 1402 2503 1413 2506
rect 1402 2446 1405 2503
rect 1418 2476 1421 2526
rect 1458 2523 1461 2606
rect 1466 2553 1469 2606
rect 1474 2593 1477 2606
rect 1482 2603 1485 2616
rect 1474 2503 1477 2536
rect 1418 2473 1429 2476
rect 1314 2413 1325 2416
rect 1306 2403 1317 2406
rect 1322 2386 1325 2413
rect 1318 2383 1325 2386
rect 1218 2313 1237 2316
rect 1258 2313 1269 2316
rect 1218 2213 1221 2313
rect 1258 2226 1261 2313
rect 1282 2293 1285 2316
rect 1290 2303 1293 2336
rect 1202 2203 1209 2206
rect 1162 2033 1189 2036
rect 1146 1973 1153 1976
rect 1146 1953 1149 1973
rect 1154 1923 1157 1936
rect 1162 1906 1165 2016
rect 1178 1966 1181 2026
rect 1186 2003 1189 2033
rect 1194 2023 1197 2116
rect 1194 1973 1197 2016
rect 1170 1963 1181 1966
rect 1170 1913 1173 1963
rect 1186 1923 1189 1946
rect 1162 1903 1181 1906
rect 1138 1893 1173 1896
rect 1138 1823 1141 1856
rect 1102 1693 1109 1696
rect 1114 1753 1125 1756
rect 1102 1636 1105 1693
rect 1098 1633 1105 1636
rect 1098 1596 1101 1633
rect 1106 1603 1109 1616
rect 1114 1613 1117 1753
rect 1122 1686 1125 1726
rect 1130 1693 1133 1736
rect 1138 1723 1141 1796
rect 1146 1723 1149 1886
rect 1154 1716 1157 1856
rect 1162 1793 1165 1886
rect 1170 1746 1173 1893
rect 1162 1743 1173 1746
rect 1162 1733 1165 1743
rect 1146 1713 1157 1716
rect 1122 1683 1133 1686
rect 1122 1606 1125 1676
rect 1114 1603 1125 1606
rect 1098 1593 1117 1596
rect 1082 1303 1085 1376
rect 1034 1243 1045 1246
rect 1034 1176 1037 1243
rect 1042 1213 1045 1236
rect 1058 1213 1061 1246
rect 1082 1213 1085 1226
rect 1042 1186 1045 1206
rect 1050 1203 1085 1206
rect 1082 1186 1085 1203
rect 1042 1183 1069 1186
rect 1034 1173 1061 1176
rect 1050 1116 1053 1136
rect 1058 1123 1061 1173
rect 1066 1123 1069 1183
rect 1078 1183 1085 1186
rect 1026 1113 1033 1116
rect 1018 1023 1021 1106
rect 1030 1026 1033 1113
rect 1026 1023 1033 1026
rect 1018 933 1021 946
rect 1026 926 1029 1023
rect 1018 923 1029 926
rect 1018 733 1021 923
rect 966 693 973 696
rect 930 663 937 666
rect 914 653 925 656
rect 882 633 889 636
rect 882 606 885 633
rect 874 603 885 606
rect 874 523 877 603
rect 890 593 893 616
rect 882 523 885 546
rect 890 533 893 576
rect 898 523 901 636
rect 914 613 917 626
rect 906 516 909 606
rect 898 513 909 516
rect 882 383 885 416
rect 890 413 893 436
rect 854 313 861 316
rect 858 266 861 313
rect 850 263 861 266
rect 786 213 797 216
rect 802 243 813 246
rect 850 243 853 263
rect 730 183 733 213
rect 738 123 741 146
rect 746 133 749 196
rect 754 116 757 126
rect 770 123 773 206
rect 786 153 789 213
rect 794 133 797 206
rect 802 123 805 243
rect 810 143 813 216
rect 818 203 821 226
rect 826 203 829 216
rect 866 213 869 226
rect 834 123 837 136
rect 874 133 877 216
rect 882 203 885 326
rect 890 323 893 336
rect 898 256 901 513
rect 914 506 917 606
rect 922 603 925 653
rect 934 596 937 663
rect 946 613 949 626
rect 930 593 937 596
rect 922 523 925 536
rect 906 483 909 506
rect 914 503 921 506
rect 906 403 909 476
rect 918 446 921 503
rect 930 463 933 593
rect 938 513 941 526
rect 918 443 925 446
rect 922 396 925 443
rect 914 393 925 396
rect 914 276 917 393
rect 914 273 921 276
rect 890 253 901 256
rect 890 223 893 253
rect 898 223 901 246
rect 906 233 909 266
rect 898 213 909 216
rect 918 206 921 273
rect 914 203 921 206
rect 882 116 885 126
rect 730 113 757 116
rect 858 113 885 116
rect 898 93 901 126
rect 906 123 909 146
rect 234 73 253 76
rect 914 73 917 203
rect 930 153 933 336
rect 938 323 941 426
rect 946 396 949 606
rect 954 443 957 636
rect 966 586 969 693
rect 978 593 981 726
rect 994 723 1005 726
rect 986 623 989 716
rect 1002 656 1005 723
rect 994 653 1005 656
rect 994 633 997 653
rect 986 613 997 616
rect 966 583 973 586
rect 962 533 965 546
rect 954 403 957 426
rect 962 413 965 466
rect 970 453 973 583
rect 986 533 989 606
rect 994 583 997 613
rect 1002 556 1005 626
rect 1010 606 1013 636
rect 1010 603 1017 606
rect 994 553 1005 556
rect 994 533 997 553
rect 1014 536 1017 603
rect 1026 583 1029 886
rect 1034 813 1037 1006
rect 1042 986 1045 1116
rect 1050 1113 1061 1116
rect 1050 1013 1053 1026
rect 1058 993 1061 1113
rect 1042 983 1061 986
rect 1042 923 1045 936
rect 1034 763 1037 806
rect 1042 803 1045 846
rect 1050 746 1053 946
rect 1058 923 1061 983
rect 1066 863 1069 1036
rect 1078 1016 1081 1183
rect 1090 1023 1093 1496
rect 1098 1343 1101 1546
rect 1098 1273 1101 1336
rect 1106 1243 1109 1536
rect 1114 1523 1117 1593
rect 1122 1526 1125 1536
rect 1130 1533 1133 1683
rect 1146 1636 1149 1713
rect 1154 1693 1165 1696
rect 1170 1693 1173 1736
rect 1146 1633 1153 1636
rect 1122 1523 1133 1526
rect 1122 1493 1125 1516
rect 1114 1256 1117 1466
rect 1122 1403 1125 1416
rect 1130 1403 1133 1523
rect 1138 1493 1141 1626
rect 1150 1586 1153 1633
rect 1146 1583 1153 1586
rect 1146 1526 1149 1583
rect 1154 1533 1157 1566
rect 1162 1533 1165 1693
rect 1170 1583 1173 1596
rect 1178 1586 1181 1903
rect 1186 1813 1189 1916
rect 1194 1813 1197 1946
rect 1202 1853 1205 2203
rect 1210 2183 1221 2186
rect 1210 2123 1213 2183
rect 1226 2146 1229 2226
rect 1258 2223 1269 2226
rect 1234 2183 1237 2216
rect 1242 2193 1245 2206
rect 1266 2176 1269 2223
rect 1282 2213 1285 2286
rect 1290 2243 1301 2246
rect 1290 2206 1293 2243
rect 1298 2213 1301 2236
rect 1282 2203 1293 2206
rect 1250 2173 1269 2176
rect 1218 2143 1229 2146
rect 1218 2116 1221 2143
rect 1210 2113 1221 2116
rect 1210 1933 1213 2113
rect 1218 2093 1221 2106
rect 1218 2013 1221 2026
rect 1218 1923 1221 1986
rect 1226 1943 1229 2136
rect 1234 2133 1237 2166
rect 1234 2076 1237 2116
rect 1242 2083 1245 2146
rect 1234 2073 1245 2076
rect 1234 2013 1237 2036
rect 1242 2013 1245 2073
rect 1242 1973 1245 2006
rect 1226 1906 1229 1926
rect 1234 1923 1245 1926
rect 1222 1903 1229 1906
rect 1210 1806 1213 1876
rect 1222 1836 1225 1903
rect 1222 1833 1229 1836
rect 1226 1813 1229 1833
rect 1186 1796 1189 1806
rect 1194 1803 1221 1806
rect 1186 1793 1197 1796
rect 1194 1726 1197 1793
rect 1202 1733 1205 1786
rect 1210 1733 1213 1796
rect 1186 1623 1189 1726
rect 1194 1723 1205 1726
rect 1202 1713 1205 1723
rect 1210 1693 1213 1726
rect 1186 1603 1189 1616
rect 1194 1603 1197 1616
rect 1178 1583 1185 1586
rect 1170 1533 1173 1556
rect 1182 1526 1185 1583
rect 1146 1523 1157 1526
rect 1122 1363 1125 1386
rect 1122 1273 1125 1346
rect 1114 1253 1121 1256
rect 1098 1066 1101 1206
rect 1106 1073 1109 1196
rect 1118 1156 1121 1253
rect 1130 1173 1133 1346
rect 1138 1333 1141 1426
rect 1114 1153 1121 1156
rect 1098 1063 1109 1066
rect 1078 1013 1085 1016
rect 1074 923 1077 946
rect 1058 823 1069 826
rect 1058 793 1061 816
rect 1050 743 1069 746
rect 1042 713 1045 736
rect 1074 726 1077 836
rect 1066 723 1077 726
rect 1042 623 1045 646
rect 1042 576 1045 616
rect 1034 573 1045 576
rect 1014 533 1025 536
rect 978 473 981 526
rect 994 516 997 526
rect 986 513 997 516
rect 986 493 989 513
rect 1002 506 1005 526
rect 994 503 1005 506
rect 946 393 965 396
rect 946 333 949 386
rect 954 333 957 346
rect 946 323 957 326
rect 962 286 965 393
rect 970 333 973 446
rect 978 403 981 416
rect 994 413 997 503
rect 1002 413 1005 426
rect 986 383 989 406
rect 994 393 997 406
rect 1010 383 1013 526
rect 1022 416 1025 533
rect 1022 413 1029 416
rect 1026 396 1029 413
rect 1034 403 1037 573
rect 1042 523 1045 566
rect 1050 453 1053 676
rect 1066 646 1069 723
rect 1066 643 1073 646
rect 1058 546 1061 626
rect 1070 576 1073 643
rect 1070 573 1077 576
rect 1074 553 1077 573
rect 1082 553 1085 1013
rect 1098 1003 1101 1016
rect 1106 996 1109 1063
rect 1098 993 1109 996
rect 1098 976 1101 993
rect 1098 973 1105 976
rect 1114 973 1117 1153
rect 1138 1136 1141 1296
rect 1146 1213 1149 1486
rect 1154 1423 1157 1523
rect 1162 1506 1165 1526
rect 1178 1523 1185 1526
rect 1162 1503 1169 1506
rect 1166 1436 1169 1503
rect 1162 1433 1169 1436
rect 1162 1416 1165 1433
rect 1154 1413 1165 1416
rect 1154 1356 1157 1413
rect 1162 1393 1165 1406
rect 1154 1353 1165 1356
rect 1146 1143 1149 1156
rect 1090 933 1093 966
rect 1090 763 1093 926
rect 1102 836 1105 973
rect 1098 833 1105 836
rect 1098 813 1101 833
rect 1114 813 1117 956
rect 1106 773 1109 806
rect 1122 746 1125 1136
rect 1138 1133 1149 1136
rect 1130 1093 1133 1126
rect 1138 1113 1141 1126
rect 1146 1053 1149 1133
rect 1154 1093 1157 1336
rect 1162 1323 1165 1353
rect 1162 1213 1165 1306
rect 1170 1213 1173 1416
rect 1178 1363 1181 1523
rect 1186 1393 1189 1416
rect 1194 1383 1197 1596
rect 1202 1473 1205 1646
rect 1210 1563 1213 1616
rect 1210 1523 1213 1556
rect 1210 1376 1213 1406
rect 1186 1373 1213 1376
rect 1178 1333 1181 1346
rect 1178 1316 1181 1326
rect 1186 1323 1189 1373
rect 1194 1333 1197 1356
rect 1202 1316 1205 1326
rect 1178 1313 1205 1316
rect 1162 1186 1165 1206
rect 1162 1183 1169 1186
rect 1166 1086 1169 1183
rect 1178 1123 1181 1256
rect 1162 1083 1169 1086
rect 1162 1036 1165 1083
rect 1186 1046 1189 1313
rect 1194 1113 1197 1296
rect 1202 1243 1205 1313
rect 1202 1106 1205 1236
rect 1210 1116 1213 1366
rect 1218 1293 1221 1803
rect 1226 1743 1229 1806
rect 1234 1733 1237 1906
rect 1242 1803 1245 1816
rect 1250 1776 1253 2173
rect 1258 2096 1261 2166
rect 1274 2133 1277 2196
rect 1282 2193 1285 2203
rect 1290 2143 1293 2196
rect 1266 2106 1269 2126
rect 1282 2113 1293 2116
rect 1282 2106 1285 2113
rect 1298 2106 1301 2206
rect 1306 2143 1309 2336
rect 1318 2296 1321 2383
rect 1330 2306 1333 2426
rect 1338 2403 1341 2446
rect 1402 2443 1413 2446
rect 1362 2393 1365 2406
rect 1370 2403 1373 2416
rect 1402 2393 1405 2426
rect 1410 2376 1413 2443
rect 1426 2416 1429 2473
rect 1426 2413 1437 2416
rect 1434 2403 1437 2413
rect 1442 2403 1445 2416
rect 1410 2373 1429 2376
rect 1346 2326 1349 2346
rect 1362 2333 1365 2356
rect 1338 2323 1357 2326
rect 1330 2303 1341 2306
rect 1318 2293 1325 2296
rect 1266 2103 1285 2106
rect 1290 2103 1301 2106
rect 1258 2093 1277 2096
rect 1258 1983 1261 2046
rect 1266 2013 1269 2026
rect 1258 1933 1261 1946
rect 1258 1883 1261 1926
rect 1266 1893 1269 1926
rect 1258 1823 1269 1826
rect 1258 1793 1261 1823
rect 1274 1816 1277 2093
rect 1290 2013 1293 2103
rect 1266 1813 1277 1816
rect 1250 1773 1257 1776
rect 1242 1716 1245 1766
rect 1234 1713 1245 1716
rect 1234 1646 1237 1713
rect 1254 1706 1257 1773
rect 1250 1703 1257 1706
rect 1234 1643 1245 1646
rect 1250 1643 1253 1703
rect 1226 1613 1229 1626
rect 1226 1506 1229 1546
rect 1234 1536 1237 1626
rect 1242 1603 1245 1643
rect 1266 1583 1269 1813
rect 1282 1803 1285 1996
rect 1290 1786 1293 1966
rect 1298 1886 1301 2096
rect 1306 2013 1309 2136
rect 1314 2083 1317 2206
rect 1322 2133 1325 2293
rect 1338 2236 1341 2303
rect 1338 2233 1357 2236
rect 1338 2216 1341 2226
rect 1330 2213 1341 2216
rect 1330 2146 1333 2213
rect 1338 2193 1341 2206
rect 1346 2173 1349 2196
rect 1354 2166 1357 2233
rect 1362 2203 1365 2256
rect 1370 2213 1373 2286
rect 1378 2213 1381 2316
rect 1378 2183 1381 2206
rect 1354 2163 1381 2166
rect 1362 2146 1365 2156
rect 1330 2143 1357 2146
rect 1362 2143 1373 2146
rect 1330 2113 1333 2143
rect 1338 2113 1341 2126
rect 1306 1893 1309 2006
rect 1314 1933 1317 1996
rect 1338 1946 1341 2026
rect 1346 2013 1349 2126
rect 1354 2116 1357 2143
rect 1370 2123 1373 2136
rect 1378 2116 1381 2163
rect 1386 2133 1389 2336
rect 1410 2333 1413 2366
rect 1426 2356 1429 2373
rect 1426 2353 1433 2356
rect 1402 2323 1413 2326
rect 1394 2133 1397 2266
rect 1418 2243 1421 2336
rect 1430 2256 1433 2353
rect 1450 2326 1453 2426
rect 1466 2413 1469 2426
rect 1450 2323 1461 2326
rect 1426 2253 1433 2256
rect 1426 2236 1429 2253
rect 1410 2233 1429 2236
rect 1442 2236 1445 2316
rect 1458 2266 1461 2323
rect 1450 2263 1461 2266
rect 1450 2243 1453 2263
rect 1442 2233 1461 2236
rect 1402 2126 1405 2216
rect 1410 2136 1413 2233
rect 1418 2223 1453 2226
rect 1418 2203 1421 2223
rect 1426 2203 1429 2216
rect 1434 2213 1445 2216
rect 1450 2213 1453 2223
rect 1434 2163 1437 2206
rect 1410 2133 1421 2136
rect 1402 2123 1413 2126
rect 1354 2113 1365 2116
rect 1378 2113 1385 2116
rect 1362 1973 1365 2016
rect 1370 1946 1373 2076
rect 1338 1943 1357 1946
rect 1330 1933 1341 1936
rect 1322 1913 1325 1926
rect 1298 1883 1317 1886
rect 1298 1813 1301 1856
rect 1306 1813 1309 1826
rect 1282 1783 1293 1786
rect 1242 1543 1245 1566
rect 1234 1533 1245 1536
rect 1242 1523 1245 1533
rect 1226 1503 1237 1506
rect 1234 1436 1237 1503
rect 1250 1493 1253 1556
rect 1274 1553 1277 1596
rect 1258 1543 1269 1546
rect 1266 1533 1277 1536
rect 1282 1533 1285 1783
rect 1290 1733 1293 1746
rect 1298 1683 1301 1756
rect 1298 1623 1301 1666
rect 1306 1633 1309 1786
rect 1314 1623 1317 1883
rect 1322 1803 1325 1906
rect 1330 1853 1333 1933
rect 1338 1906 1341 1926
rect 1346 1913 1349 1936
rect 1338 1903 1349 1906
rect 1330 1786 1333 1846
rect 1326 1783 1333 1786
rect 1326 1686 1329 1783
rect 1326 1683 1333 1686
rect 1330 1663 1333 1683
rect 1338 1656 1341 1896
rect 1346 1826 1349 1903
rect 1354 1873 1357 1943
rect 1362 1943 1373 1946
rect 1382 1946 1385 2113
rect 1382 1943 1389 1946
rect 1362 1923 1365 1943
rect 1370 1886 1373 1926
rect 1362 1883 1373 1886
rect 1370 1833 1373 1876
rect 1378 1826 1381 1936
rect 1346 1823 1357 1826
rect 1346 1803 1349 1816
rect 1354 1783 1357 1823
rect 1362 1823 1381 1826
rect 1362 1753 1365 1823
rect 1346 1663 1349 1736
rect 1370 1733 1373 1806
rect 1378 1763 1381 1816
rect 1386 1806 1389 1943
rect 1394 1906 1397 2036
rect 1402 2013 1405 2116
rect 1410 2013 1413 2123
rect 1402 1913 1413 1916
rect 1418 1913 1421 2133
rect 1426 1953 1429 2126
rect 1434 2083 1437 2136
rect 1442 2123 1445 2206
rect 1450 2183 1453 2206
rect 1458 2176 1461 2233
rect 1450 2173 1461 2176
rect 1466 2203 1477 2206
rect 1434 1996 1437 2006
rect 1442 2003 1445 2026
rect 1450 2013 1453 2173
rect 1458 2093 1461 2126
rect 1466 2123 1469 2203
rect 1474 2113 1477 2136
rect 1458 2003 1461 2016
rect 1466 2013 1469 2036
rect 1474 2013 1477 2026
rect 1466 1996 1469 2006
rect 1434 1993 1469 1996
rect 1394 1903 1405 1906
rect 1394 1813 1397 1866
rect 1386 1803 1393 1806
rect 1402 1803 1405 1903
rect 1410 1813 1413 1913
rect 1426 1903 1429 1936
rect 1434 1923 1437 1993
rect 1442 1916 1445 1976
rect 1434 1913 1445 1916
rect 1418 1803 1421 1876
rect 1390 1746 1393 1803
rect 1426 1776 1429 1896
rect 1434 1843 1437 1913
rect 1450 1896 1453 1966
rect 1442 1893 1453 1896
rect 1434 1786 1437 1816
rect 1442 1793 1445 1893
rect 1466 1886 1469 1926
rect 1454 1883 1469 1886
rect 1434 1783 1445 1786
rect 1426 1773 1437 1776
rect 1390 1743 1397 1746
rect 1354 1723 1381 1726
rect 1330 1653 1341 1656
rect 1226 1433 1237 1436
rect 1226 1286 1229 1433
rect 1234 1363 1237 1416
rect 1222 1283 1229 1286
rect 1222 1176 1225 1283
rect 1234 1233 1237 1356
rect 1242 1313 1245 1416
rect 1250 1306 1253 1476
rect 1274 1456 1277 1533
rect 1274 1453 1285 1456
rect 1258 1406 1261 1426
rect 1266 1413 1269 1436
rect 1258 1403 1269 1406
rect 1282 1403 1285 1453
rect 1290 1433 1293 1616
rect 1290 1396 1293 1426
rect 1258 1393 1293 1396
rect 1258 1353 1261 1393
rect 1258 1316 1261 1346
rect 1266 1333 1269 1386
rect 1274 1323 1277 1336
rect 1282 1333 1293 1336
rect 1282 1316 1285 1326
rect 1258 1313 1285 1316
rect 1250 1303 1277 1306
rect 1242 1213 1245 1226
rect 1258 1213 1261 1246
rect 1274 1236 1277 1303
rect 1274 1233 1285 1236
rect 1218 1173 1225 1176
rect 1218 1123 1221 1173
rect 1210 1113 1221 1116
rect 1202 1103 1209 1106
rect 1186 1043 1197 1046
rect 1130 1033 1165 1036
rect 1130 853 1133 1033
rect 1138 1023 1173 1026
rect 1138 926 1141 1016
rect 1146 983 1149 1006
rect 1154 1003 1157 1016
rect 1146 933 1149 966
rect 1162 933 1165 996
rect 1170 956 1173 1006
rect 1178 963 1181 1006
rect 1186 983 1189 996
rect 1170 953 1189 956
rect 1194 953 1197 1043
rect 1206 1006 1209 1103
rect 1218 1013 1221 1113
rect 1226 1096 1229 1136
rect 1234 1113 1237 1206
rect 1242 1133 1245 1166
rect 1242 1113 1245 1126
rect 1226 1093 1233 1096
rect 1230 1026 1233 1093
rect 1226 1023 1233 1026
rect 1206 1003 1213 1006
rect 1210 953 1213 1003
rect 1138 923 1149 926
rect 1146 906 1149 923
rect 1154 913 1157 926
rect 1162 923 1173 926
rect 1178 923 1181 946
rect 1162 906 1165 923
rect 1142 903 1149 906
rect 1154 903 1165 906
rect 1130 803 1133 846
rect 1142 836 1145 903
rect 1142 833 1149 836
rect 1138 803 1141 816
rect 1146 796 1149 833
rect 1090 743 1125 746
rect 1138 793 1149 796
rect 1138 743 1141 793
rect 1090 613 1093 743
rect 1122 716 1125 736
rect 1114 713 1125 716
rect 1114 656 1117 713
rect 1114 653 1125 656
rect 1106 613 1109 636
rect 1114 603 1117 616
rect 1058 543 1109 546
rect 1058 533 1061 543
rect 1058 463 1061 526
rect 1066 516 1069 536
rect 1106 533 1109 543
rect 1066 513 1077 516
rect 1074 456 1077 513
rect 1058 453 1077 456
rect 1050 396 1053 406
rect 1026 393 1053 396
rect 1010 346 1013 366
rect 1002 336 1005 346
rect 1010 343 1021 346
rect 978 333 1005 336
rect 938 283 965 286
rect 938 233 941 283
rect 970 223 973 246
rect 978 213 981 333
rect 994 246 997 326
rect 1018 296 1021 343
rect 1010 293 1021 296
rect 1042 293 1045 316
rect 1058 313 1061 453
rect 994 243 1005 246
rect 994 176 997 226
rect 1002 193 1005 243
rect 1010 213 1013 293
rect 1018 256 1021 276
rect 1018 253 1029 256
rect 1026 206 1029 253
rect 946 173 997 176
rect 946 133 949 173
rect 954 83 957 136
rect 970 133 973 166
rect 962 113 965 126
rect 986 103 989 136
rect 1010 123 1013 206
rect 1018 203 1029 206
rect 1018 123 1021 203
rect 1042 196 1045 216
rect 1050 203 1053 256
rect 1058 213 1061 226
rect 1058 196 1061 206
rect 1042 193 1061 196
rect 1066 186 1069 326
rect 1074 293 1077 426
rect 1082 253 1085 416
rect 1090 313 1093 396
rect 1098 323 1101 526
rect 1106 473 1109 526
rect 1122 516 1125 653
rect 1130 613 1133 726
rect 1138 713 1141 736
rect 1146 723 1149 786
rect 1154 733 1157 903
rect 1162 723 1165 896
rect 1138 533 1141 616
rect 1146 596 1149 706
rect 1154 676 1157 716
rect 1162 703 1165 716
rect 1170 703 1173 856
rect 1178 816 1181 916
rect 1186 853 1189 953
rect 1194 933 1205 936
rect 1194 876 1197 933
rect 1218 913 1221 936
rect 1194 873 1213 876
rect 1194 816 1197 836
rect 1178 813 1189 816
rect 1194 813 1205 816
rect 1178 763 1181 806
rect 1154 673 1173 676
rect 1154 603 1157 666
rect 1170 636 1173 673
rect 1178 643 1181 716
rect 1186 636 1189 813
rect 1194 663 1197 806
rect 1210 803 1213 873
rect 1218 853 1221 886
rect 1218 786 1221 826
rect 1214 783 1221 786
rect 1170 633 1189 636
rect 1146 593 1157 596
rect 1114 443 1117 516
rect 1122 513 1133 516
rect 1130 446 1133 513
rect 1122 443 1133 446
rect 1146 446 1149 526
rect 1154 513 1157 593
rect 1162 493 1165 586
rect 1170 533 1173 633
rect 1194 603 1197 626
rect 1202 613 1205 746
rect 1214 686 1217 783
rect 1214 683 1221 686
rect 1186 533 1189 566
rect 1210 553 1213 666
rect 1202 533 1213 536
rect 1218 533 1221 683
rect 1226 556 1229 1023
rect 1234 803 1237 1006
rect 1242 913 1245 1096
rect 1250 1063 1253 1206
rect 1242 813 1245 826
rect 1242 773 1245 806
rect 1234 733 1237 756
rect 1242 703 1245 726
rect 1234 566 1237 696
rect 1242 613 1245 686
rect 1250 613 1253 1026
rect 1258 943 1261 1146
rect 1266 1123 1269 1206
rect 1258 623 1261 936
rect 1266 823 1269 1116
rect 1274 1013 1277 1216
rect 1282 1023 1285 1233
rect 1274 983 1277 1006
rect 1282 976 1285 1016
rect 1274 973 1285 976
rect 1274 943 1277 973
rect 1282 936 1285 956
rect 1278 933 1285 936
rect 1278 846 1281 933
rect 1274 843 1281 846
rect 1266 713 1269 796
rect 1274 743 1277 843
rect 1282 756 1285 826
rect 1290 793 1293 1333
rect 1298 1253 1301 1596
rect 1314 1576 1317 1616
rect 1322 1603 1325 1636
rect 1306 1573 1317 1576
rect 1306 1393 1309 1573
rect 1314 1376 1317 1566
rect 1330 1533 1333 1653
rect 1338 1593 1341 1606
rect 1346 1583 1349 1626
rect 1370 1613 1373 1646
rect 1322 1433 1325 1526
rect 1338 1506 1341 1536
rect 1346 1523 1349 1536
rect 1354 1513 1357 1606
rect 1378 1596 1381 1723
rect 1386 1713 1389 1726
rect 1386 1613 1389 1636
rect 1362 1593 1381 1596
rect 1338 1503 1349 1506
rect 1310 1373 1317 1376
rect 1310 1316 1313 1373
rect 1322 1323 1325 1366
rect 1310 1313 1317 1316
rect 1298 1033 1301 1206
rect 1298 943 1301 1016
rect 1306 936 1309 1286
rect 1314 1083 1317 1313
rect 1322 1213 1325 1226
rect 1322 1123 1325 1156
rect 1330 1123 1333 1436
rect 1338 1283 1341 1496
rect 1346 1483 1349 1503
rect 1346 1423 1357 1426
rect 1346 1413 1357 1416
rect 1362 1406 1365 1593
rect 1394 1563 1397 1743
rect 1402 1736 1405 1756
rect 1402 1733 1409 1736
rect 1406 1636 1409 1733
rect 1418 1723 1421 1766
rect 1418 1703 1421 1716
rect 1402 1633 1409 1636
rect 1402 1603 1405 1633
rect 1410 1586 1413 1616
rect 1406 1583 1413 1586
rect 1370 1533 1373 1546
rect 1386 1536 1389 1556
rect 1382 1533 1389 1536
rect 1354 1403 1365 1406
rect 1362 1336 1365 1396
rect 1346 1266 1349 1336
rect 1342 1263 1349 1266
rect 1354 1333 1365 1336
rect 1342 1186 1345 1263
rect 1354 1203 1357 1333
rect 1362 1213 1365 1326
rect 1342 1183 1349 1186
rect 1322 993 1325 1106
rect 1338 1016 1341 1166
rect 1346 1153 1349 1183
rect 1362 1116 1365 1136
rect 1346 1103 1349 1116
rect 1358 1113 1365 1116
rect 1358 1046 1361 1113
rect 1358 1043 1365 1046
rect 1362 1023 1365 1043
rect 1338 1013 1357 1016
rect 1314 943 1317 986
rect 1298 843 1301 936
rect 1306 933 1317 936
rect 1314 923 1317 933
rect 1322 903 1325 936
rect 1298 813 1301 836
rect 1314 813 1317 826
rect 1282 753 1293 756
rect 1274 723 1277 736
rect 1282 716 1285 736
rect 1274 713 1285 716
rect 1290 713 1293 753
rect 1274 693 1277 713
rect 1250 603 1261 606
rect 1234 563 1261 566
rect 1226 553 1245 556
rect 1210 526 1213 533
rect 1202 446 1205 526
rect 1210 523 1221 526
rect 1210 513 1221 516
rect 1218 493 1221 513
rect 1226 506 1229 526
rect 1226 503 1233 506
rect 1146 443 1165 446
rect 1202 443 1209 446
rect 1122 423 1125 443
rect 1130 423 1157 426
rect 1122 306 1125 406
rect 1130 373 1133 423
rect 1138 413 1157 416
rect 1114 303 1125 306
rect 1114 246 1117 303
rect 1114 243 1125 246
rect 1098 223 1117 226
rect 1050 183 1069 186
rect 1034 113 1045 116
rect 1050 83 1053 183
rect 1058 116 1061 136
rect 1074 123 1077 136
rect 1082 116 1085 186
rect 1098 123 1101 223
rect 1122 213 1125 243
rect 1130 233 1133 296
rect 1138 223 1141 396
rect 1154 393 1157 406
rect 1162 403 1165 443
rect 1146 213 1149 296
rect 1162 283 1165 336
rect 1170 333 1173 356
rect 1178 323 1181 406
rect 1186 333 1189 416
rect 1194 413 1197 436
rect 1194 306 1197 406
rect 1206 356 1209 443
rect 1218 396 1221 466
rect 1230 436 1233 503
rect 1226 433 1233 436
rect 1226 403 1229 433
rect 1242 416 1245 553
rect 1234 413 1245 416
rect 1218 393 1229 396
rect 1186 303 1197 306
rect 1202 353 1209 356
rect 1162 206 1165 256
rect 1186 226 1189 303
rect 1158 203 1165 206
rect 1170 223 1189 226
rect 1058 113 1085 116
rect 1114 93 1117 126
rect 1122 123 1125 156
rect 1158 146 1161 203
rect 1154 143 1161 146
rect 1154 133 1157 143
rect 1170 93 1173 223
rect 1178 133 1181 176
rect 1194 173 1197 216
rect 1178 116 1181 126
rect 1186 123 1189 166
rect 1194 116 1197 126
rect 1202 123 1205 353
rect 1210 303 1213 336
rect 1218 323 1221 336
rect 1226 306 1229 393
rect 1222 303 1229 306
rect 1222 236 1225 303
rect 1222 233 1229 236
rect 1210 193 1213 206
rect 1218 123 1221 216
rect 1226 153 1229 233
rect 1178 113 1197 116
rect 1226 93 1229 136
rect 1234 43 1237 413
rect 1242 383 1245 406
rect 1250 393 1253 406
rect 1258 386 1261 563
rect 1266 533 1269 566
rect 1274 446 1277 666
rect 1282 633 1285 706
rect 1282 603 1285 616
rect 1290 603 1293 656
rect 1298 586 1301 776
rect 1306 753 1309 806
rect 1314 803 1325 806
rect 1330 786 1333 1006
rect 1338 993 1357 996
rect 1362 976 1365 1006
rect 1354 973 1365 976
rect 1338 813 1341 836
rect 1354 796 1357 973
rect 1370 956 1373 1486
rect 1382 1436 1385 1533
rect 1406 1526 1409 1583
rect 1418 1533 1421 1666
rect 1426 1636 1429 1706
rect 1434 1643 1437 1773
rect 1442 1706 1445 1783
rect 1454 1756 1457 1883
rect 1466 1813 1469 1846
rect 1474 1833 1477 1996
rect 1482 1826 1485 2426
rect 1498 2403 1501 2526
rect 1514 2523 1517 2633
rect 1530 2613 1533 2726
rect 1546 2706 1549 2736
rect 1554 2723 1557 2853
rect 1562 2813 1565 2926
rect 1570 2906 1573 2926
rect 1570 2903 1577 2906
rect 1574 2836 1577 2903
rect 1594 2886 1597 2933
rect 1618 2923 1621 2986
rect 1626 2933 1629 2996
rect 1642 2933 1645 3016
rect 1650 3003 1653 3103
rect 1658 3013 1661 3036
rect 1714 3023 1717 3036
rect 1666 3013 1677 3016
rect 1634 2916 1637 2926
rect 1650 2923 1653 2976
rect 1666 2923 1669 2986
rect 1682 2983 1685 3006
rect 1690 2973 1693 3006
rect 1698 2956 1701 3016
rect 1714 2993 1717 3006
rect 1722 2986 1725 3056
rect 1730 3003 1733 3026
rect 1714 2983 1725 2986
rect 1698 2953 1709 2956
rect 1698 2933 1701 2946
rect 1706 2933 1709 2953
rect 1610 2913 1637 2916
rect 1594 2883 1621 2886
rect 1570 2833 1577 2836
rect 1570 2806 1573 2833
rect 1562 2803 1573 2806
rect 1562 2743 1565 2803
rect 1578 2783 1581 2816
rect 1578 2713 1581 2726
rect 1546 2703 1557 2706
rect 1554 2646 1557 2703
rect 1546 2643 1557 2646
rect 1522 2543 1525 2606
rect 1522 2486 1525 2506
rect 1546 2486 1549 2643
rect 1602 2613 1605 2736
rect 1610 2733 1613 2816
rect 1618 2803 1621 2883
rect 1706 2856 1709 2926
rect 1714 2906 1717 2983
rect 1722 2933 1725 2976
rect 1754 2973 1757 3126
rect 1770 3103 1773 3126
rect 1782 3086 1785 3133
rect 1802 3106 1805 3183
rect 1810 3133 1813 3146
rect 1802 3103 1809 3106
rect 1818 3103 1821 3206
rect 1826 3203 1829 3216
rect 1842 3213 1853 3216
rect 1866 3213 1869 3246
rect 1842 3176 1845 3213
rect 1858 3183 1861 3206
rect 1842 3173 1861 3176
rect 1834 3133 1845 3136
rect 1778 3083 1785 3086
rect 1730 2923 1733 2966
rect 1714 2903 1725 2906
rect 1674 2853 1709 2856
rect 1674 2823 1677 2853
rect 1722 2836 1725 2903
rect 1754 2883 1757 2926
rect 1762 2916 1765 3016
rect 1778 3013 1781 3083
rect 1770 2983 1773 3006
rect 1786 3003 1789 3026
rect 1770 2933 1773 2946
rect 1762 2913 1773 2916
rect 1778 2913 1781 2926
rect 1718 2833 1725 2836
rect 1642 2743 1645 2816
rect 1658 2783 1661 2806
rect 1690 2793 1693 2806
rect 1718 2776 1721 2833
rect 1738 2793 1741 2816
rect 1714 2773 1721 2776
rect 1714 2753 1717 2773
rect 1770 2746 1773 2816
rect 1666 2743 1717 2746
rect 1666 2733 1669 2743
rect 1666 2713 1669 2726
rect 1562 2533 1565 2596
rect 1578 2583 1581 2606
rect 1610 2533 1613 2556
rect 1658 2533 1661 2616
rect 1666 2533 1669 2596
rect 1522 2483 1533 2486
rect 1546 2483 1557 2486
rect 1530 2403 1533 2483
rect 1554 2423 1557 2483
rect 1498 2333 1501 2356
rect 1522 2323 1525 2346
rect 1530 2333 1533 2396
rect 1562 2366 1565 2436
rect 1578 2393 1581 2416
rect 1554 2363 1565 2366
rect 1490 2296 1493 2316
rect 1490 2293 1501 2296
rect 1522 2293 1525 2316
rect 1498 2226 1501 2293
rect 1490 2223 1501 2226
rect 1490 2203 1493 2223
rect 1506 2193 1509 2206
rect 1490 2003 1493 2136
rect 1498 1996 1501 2106
rect 1490 1993 1501 1996
rect 1490 1893 1493 1993
rect 1482 1823 1493 1826
rect 1466 1763 1469 1806
rect 1450 1753 1457 1756
rect 1450 1733 1453 1753
rect 1474 1733 1477 1806
rect 1450 1713 1453 1726
rect 1482 1723 1485 1816
rect 1442 1703 1453 1706
rect 1426 1633 1437 1636
rect 1426 1613 1429 1626
rect 1434 1596 1437 1633
rect 1430 1593 1437 1596
rect 1430 1526 1433 1593
rect 1382 1433 1389 1436
rect 1378 1403 1381 1416
rect 1386 1393 1389 1433
rect 1378 1343 1381 1366
rect 1386 1336 1389 1386
rect 1378 1333 1389 1336
rect 1394 1333 1397 1526
rect 1406 1523 1413 1526
rect 1410 1443 1413 1523
rect 1426 1523 1433 1526
rect 1426 1506 1429 1523
rect 1422 1503 1429 1506
rect 1422 1426 1425 1503
rect 1434 1443 1437 1516
rect 1442 1436 1445 1686
rect 1450 1653 1453 1703
rect 1490 1666 1493 1823
rect 1458 1663 1493 1666
rect 1450 1523 1453 1626
rect 1458 1586 1461 1663
rect 1466 1603 1469 1616
rect 1474 1603 1477 1656
rect 1498 1646 1501 1956
rect 1506 1946 1509 2136
rect 1514 2123 1517 2176
rect 1522 2133 1525 2276
rect 1554 2266 1557 2363
rect 1570 2276 1573 2336
rect 1578 2326 1581 2386
rect 1594 2333 1597 2356
rect 1578 2323 1593 2326
rect 1570 2273 1581 2276
rect 1554 2263 1573 2266
rect 1530 2213 1533 2226
rect 1546 2196 1549 2246
rect 1554 2213 1557 2226
rect 1530 2123 1533 2146
rect 1538 2083 1541 2196
rect 1546 2193 1553 2196
rect 1550 2076 1553 2193
rect 1562 2106 1565 2216
rect 1570 2153 1573 2263
rect 1570 2123 1573 2136
rect 1578 2123 1581 2273
rect 1590 2246 1593 2323
rect 1590 2243 1597 2246
rect 1586 2203 1589 2226
rect 1586 2133 1589 2146
rect 1562 2103 1573 2106
rect 1514 1993 1517 2076
rect 1546 2073 1553 2076
rect 1522 1973 1525 2056
rect 1506 1943 1517 1946
rect 1506 1933 1533 1936
rect 1530 1923 1533 1933
rect 1506 1813 1509 1846
rect 1506 1763 1509 1806
rect 1506 1703 1509 1726
rect 1506 1663 1509 1696
rect 1490 1643 1501 1646
rect 1482 1613 1485 1636
rect 1490 1626 1493 1643
rect 1498 1633 1509 1636
rect 1490 1623 1501 1626
rect 1498 1613 1501 1623
rect 1458 1583 1477 1586
rect 1434 1433 1445 1436
rect 1378 1233 1381 1333
rect 1386 1306 1389 1326
rect 1386 1303 1393 1306
rect 1390 1226 1393 1303
rect 1378 1213 1381 1226
rect 1386 1223 1393 1226
rect 1378 1113 1381 1126
rect 1378 983 1381 1036
rect 1386 1003 1389 1223
rect 1394 1183 1397 1206
rect 1402 1123 1405 1426
rect 1422 1423 1429 1426
rect 1418 1393 1421 1406
rect 1410 1293 1413 1336
rect 1418 1303 1421 1326
rect 1426 1236 1429 1423
rect 1434 1323 1437 1433
rect 1450 1423 1453 1516
rect 1458 1503 1461 1576
rect 1474 1526 1477 1583
rect 1490 1533 1493 1606
rect 1474 1523 1485 1526
rect 1442 1403 1445 1416
rect 1450 1413 1461 1416
rect 1450 1323 1453 1336
rect 1450 1286 1453 1306
rect 1446 1283 1453 1286
rect 1426 1233 1437 1236
rect 1418 1213 1421 1226
rect 1410 1163 1413 1206
rect 1394 1013 1397 1076
rect 1410 1046 1413 1136
rect 1402 1043 1413 1046
rect 1366 953 1373 956
rect 1366 876 1369 953
rect 1378 933 1389 936
rect 1378 886 1381 926
rect 1386 903 1389 926
rect 1394 893 1397 926
rect 1378 883 1385 886
rect 1402 883 1405 1043
rect 1418 1036 1421 1196
rect 1434 1176 1437 1233
rect 1446 1206 1449 1283
rect 1458 1253 1461 1406
rect 1466 1403 1469 1496
rect 1474 1393 1477 1416
rect 1482 1356 1485 1523
rect 1506 1516 1509 1546
rect 1498 1513 1509 1516
rect 1498 1446 1501 1513
rect 1514 1456 1517 1916
rect 1522 1893 1525 1916
rect 1522 1813 1525 1856
rect 1522 1793 1525 1806
rect 1522 1723 1525 1766
rect 1522 1703 1525 1716
rect 1530 1683 1533 1916
rect 1538 1903 1541 1936
rect 1546 1913 1549 2073
rect 1570 2056 1573 2103
rect 1562 2053 1573 2056
rect 1594 2053 1597 2243
rect 1562 2033 1565 2053
rect 1554 2023 1597 2026
rect 1554 2013 1557 2023
rect 1562 2013 1573 2016
rect 1570 1973 1573 2006
rect 1554 1923 1557 1936
rect 1562 1906 1565 1936
rect 1578 1926 1581 2016
rect 1594 2013 1597 2023
rect 1578 1923 1597 1926
rect 1558 1903 1565 1906
rect 1538 1813 1541 1896
rect 1538 1656 1541 1716
rect 1530 1653 1541 1656
rect 1546 1636 1549 1866
rect 1558 1836 1561 1903
rect 1558 1833 1565 1836
rect 1554 1733 1557 1816
rect 1530 1623 1533 1636
rect 1542 1633 1549 1636
rect 1522 1613 1533 1616
rect 1522 1533 1525 1556
rect 1542 1546 1545 1633
rect 1530 1533 1533 1546
rect 1542 1543 1549 1546
rect 1522 1473 1525 1526
rect 1538 1503 1541 1526
rect 1546 1496 1549 1543
rect 1554 1533 1557 1636
rect 1562 1613 1565 1833
rect 1562 1583 1565 1606
rect 1530 1493 1549 1496
rect 1514 1453 1521 1456
rect 1498 1443 1509 1446
rect 1474 1353 1485 1356
rect 1458 1213 1461 1226
rect 1446 1203 1453 1206
rect 1426 1173 1437 1176
rect 1426 1043 1429 1173
rect 1434 1036 1437 1126
rect 1442 1043 1445 1156
rect 1450 1106 1453 1203
rect 1466 1146 1469 1326
rect 1474 1286 1477 1353
rect 1490 1346 1493 1426
rect 1482 1343 1493 1346
rect 1482 1303 1485 1343
rect 1474 1283 1481 1286
rect 1478 1216 1481 1283
rect 1478 1213 1485 1216
rect 1490 1213 1493 1336
rect 1498 1313 1501 1416
rect 1506 1263 1509 1443
rect 1518 1386 1521 1453
rect 1514 1383 1521 1386
rect 1466 1143 1477 1146
rect 1458 1113 1461 1126
rect 1450 1103 1461 1106
rect 1410 1033 1421 1036
rect 1426 1033 1453 1036
rect 1410 1013 1413 1033
rect 1410 936 1413 1006
rect 1418 1003 1421 1026
rect 1426 1013 1429 1033
rect 1450 1023 1453 1033
rect 1442 963 1445 1016
rect 1450 993 1453 1016
rect 1458 986 1461 1103
rect 1450 983 1461 986
rect 1410 933 1417 936
rect 1366 873 1373 876
rect 1354 793 1365 796
rect 1326 783 1333 786
rect 1290 583 1301 586
rect 1290 536 1293 583
rect 1290 533 1301 536
rect 1306 533 1309 616
rect 1298 513 1301 533
rect 1306 463 1309 526
rect 1250 383 1261 386
rect 1270 443 1277 446
rect 1270 386 1273 443
rect 1282 413 1285 436
rect 1282 393 1285 406
rect 1270 383 1277 386
rect 1242 213 1245 356
rect 1250 306 1253 383
rect 1258 323 1261 376
rect 1266 343 1269 356
rect 1250 303 1257 306
rect 1254 236 1257 303
rect 1250 233 1257 236
rect 1250 213 1253 233
rect 1242 193 1245 206
rect 1258 193 1261 216
rect 1266 173 1269 336
rect 1274 283 1277 383
rect 1290 353 1293 406
rect 1298 393 1301 456
rect 1282 333 1293 336
rect 1298 326 1301 386
rect 1306 343 1309 416
rect 1314 393 1317 776
rect 1326 626 1329 783
rect 1362 773 1365 793
rect 1370 776 1373 873
rect 1382 796 1385 883
rect 1414 866 1417 933
rect 1414 863 1421 866
rect 1402 813 1405 826
rect 1394 803 1405 806
rect 1410 803 1413 846
rect 1418 803 1421 863
rect 1426 846 1429 936
rect 1442 863 1445 956
rect 1426 843 1437 846
rect 1434 796 1437 843
rect 1382 793 1397 796
rect 1370 773 1377 776
rect 1326 623 1333 626
rect 1330 603 1333 623
rect 1338 616 1341 756
rect 1346 683 1349 726
rect 1354 623 1357 636
rect 1362 633 1365 746
rect 1374 676 1377 773
rect 1370 673 1377 676
rect 1370 626 1373 673
rect 1378 633 1381 656
rect 1386 646 1389 736
rect 1394 713 1397 793
rect 1426 793 1437 796
rect 1402 723 1405 776
rect 1426 733 1429 793
rect 1450 766 1453 983
rect 1458 923 1461 936
rect 1466 916 1469 1126
rect 1474 1103 1477 1143
rect 1474 1003 1477 1096
rect 1482 1086 1485 1213
rect 1498 1193 1501 1206
rect 1490 1093 1493 1116
rect 1506 1103 1509 1186
rect 1482 1083 1509 1086
rect 1482 986 1485 1006
rect 1458 913 1469 916
rect 1478 983 1485 986
rect 1478 916 1481 983
rect 1490 923 1493 1016
rect 1498 993 1501 1026
rect 1498 933 1501 966
rect 1478 913 1485 916
rect 1458 903 1461 913
rect 1458 813 1461 896
rect 1450 763 1457 766
rect 1442 716 1445 756
rect 1402 713 1421 716
rect 1434 713 1445 716
rect 1402 703 1405 713
rect 1410 693 1413 706
rect 1418 646 1421 666
rect 1386 643 1397 646
rect 1362 616 1365 626
rect 1370 623 1381 626
rect 1386 623 1389 636
rect 1338 613 1365 616
rect 1322 516 1325 576
rect 1330 533 1333 566
rect 1346 546 1349 606
rect 1342 543 1349 546
rect 1322 513 1333 516
rect 1330 426 1333 513
rect 1322 423 1333 426
rect 1342 426 1345 543
rect 1342 423 1349 426
rect 1282 286 1285 326
rect 1290 293 1293 326
rect 1298 323 1309 326
rect 1314 286 1317 336
rect 1322 333 1325 423
rect 1346 406 1349 423
rect 1338 403 1349 406
rect 1282 283 1317 286
rect 1330 286 1333 336
rect 1330 283 1349 286
rect 1282 203 1285 246
rect 1298 223 1317 226
rect 1298 216 1301 223
rect 1290 213 1301 216
rect 1242 126 1245 166
rect 1298 153 1301 206
rect 1314 146 1317 223
rect 1330 213 1333 256
rect 1338 223 1341 276
rect 1314 143 1325 146
rect 1330 143 1333 206
rect 1346 203 1349 283
rect 1354 213 1357 536
rect 1362 533 1365 613
rect 1370 516 1373 536
rect 1366 513 1373 516
rect 1366 436 1369 513
rect 1378 453 1381 623
rect 1394 533 1397 643
rect 1402 603 1405 646
rect 1418 643 1425 646
rect 1394 513 1397 526
rect 1410 523 1413 626
rect 1422 566 1425 643
rect 1434 636 1437 713
rect 1454 706 1457 763
rect 1466 723 1469 866
rect 1474 823 1477 856
rect 1482 813 1485 913
rect 1498 893 1501 916
rect 1450 703 1457 706
rect 1450 643 1453 703
rect 1434 633 1445 636
rect 1418 563 1425 566
rect 1418 533 1421 563
rect 1434 506 1437 616
rect 1442 606 1445 633
rect 1458 613 1461 626
rect 1466 606 1469 686
rect 1474 663 1477 806
rect 1490 803 1493 826
rect 1482 733 1485 776
rect 1490 743 1493 766
rect 1506 756 1509 1083
rect 1514 903 1517 1383
rect 1522 1333 1525 1366
rect 1522 1213 1525 1256
rect 1522 1133 1525 1196
rect 1522 1073 1525 1116
rect 1522 1013 1525 1036
rect 1522 923 1525 1006
rect 1530 863 1533 1493
rect 1554 1463 1557 1516
rect 1538 1403 1541 1446
rect 1562 1426 1565 1516
rect 1570 1473 1573 1916
rect 1586 1913 1597 1916
rect 1578 1803 1581 1846
rect 1586 1813 1589 1896
rect 1578 1683 1581 1786
rect 1586 1733 1589 1806
rect 1594 1776 1597 1913
rect 1602 1863 1605 2526
rect 1618 2523 1629 2526
rect 1618 2413 1621 2523
rect 1642 2403 1645 2506
rect 1666 2396 1669 2416
rect 1658 2393 1669 2396
rect 1618 2323 1621 2376
rect 1634 2333 1637 2346
rect 1658 2333 1661 2393
rect 1674 2386 1677 2736
rect 1714 2613 1717 2743
rect 1722 2743 1773 2746
rect 1722 2733 1725 2743
rect 1778 2736 1781 2816
rect 1786 2803 1789 2816
rect 1794 2796 1797 3076
rect 1806 3036 1809 3103
rect 1842 3066 1845 3126
rect 1802 3033 1809 3036
rect 1834 3063 1845 3066
rect 1802 3016 1805 3033
rect 1802 3013 1821 3016
rect 1802 2933 1805 2946
rect 1818 2933 1821 3013
rect 1826 2993 1829 3016
rect 1834 2983 1837 3063
rect 1850 3056 1853 3106
rect 1842 3053 1853 3056
rect 1842 3013 1845 3053
rect 1850 3003 1853 3026
rect 1858 3013 1861 3173
rect 1866 3086 1869 3146
rect 1874 3123 1877 3340
rect 1938 3253 1941 3340
rect 1906 3233 1933 3236
rect 1906 3213 1909 3233
rect 1930 3216 1933 3226
rect 1882 3193 1893 3196
rect 1882 3093 1885 3106
rect 1890 3103 1893 3116
rect 1866 3083 1893 3086
rect 1866 3013 1869 3076
rect 1890 3046 1893 3083
rect 1898 3053 1901 3136
rect 1906 3096 1909 3126
rect 1914 3113 1917 3216
rect 1922 3213 1933 3216
rect 1938 3213 1941 3236
rect 1954 3223 1957 3236
rect 1922 3193 1925 3206
rect 1930 3166 1933 3213
rect 1962 3193 1965 3236
rect 1930 3163 1941 3166
rect 1938 3123 1941 3163
rect 1970 3153 1973 3340
rect 1978 3183 1981 3226
rect 1986 3213 1989 3246
rect 2002 3236 2005 3340
rect 2290 3266 2293 3340
rect 2330 3286 2333 3340
rect 2330 3283 2341 3286
rect 2234 3263 2293 3266
rect 2090 3253 2117 3256
rect 1998 3233 2005 3236
rect 1998 3186 2001 3233
rect 1998 3183 2005 3186
rect 2002 3163 2005 3183
rect 2010 3153 2013 3226
rect 2018 3183 2021 3206
rect 2026 3203 2029 3216
rect 2034 3176 2037 3216
rect 2042 3206 2045 3226
rect 2066 3216 2069 3236
rect 2066 3213 2085 3216
rect 2090 3213 2093 3253
rect 2098 3213 2101 3246
rect 2114 3223 2117 3253
rect 2162 3236 2165 3256
rect 2154 3233 2165 3236
rect 2122 3213 2125 3226
rect 2042 3203 2053 3206
rect 2018 3173 2037 3176
rect 1978 3133 1981 3146
rect 1994 3133 2013 3136
rect 2018 3133 2021 3173
rect 2050 3156 2053 3203
rect 2042 3153 2053 3156
rect 2010 3126 2013 3133
rect 1954 3123 1973 3126
rect 2010 3123 2021 3126
rect 1906 3093 1917 3096
rect 1914 3046 1917 3093
rect 1890 3043 1901 3046
rect 1882 3013 1885 3036
rect 1898 3016 1901 3043
rect 1906 3043 1917 3046
rect 1906 3023 1909 3043
rect 1898 3013 1909 3016
rect 1930 3013 1933 3026
rect 1946 3023 1949 3036
rect 1954 3013 1957 3066
rect 1890 2986 1893 3006
rect 1882 2983 1893 2986
rect 1810 2823 1813 2926
rect 1826 2903 1829 2966
rect 1842 2836 1845 2936
rect 1858 2933 1861 2976
rect 1898 2973 1901 3006
rect 1906 2963 1909 3013
rect 1930 3003 1949 3006
rect 1962 3003 1973 3006
rect 1906 2933 1909 2946
rect 1890 2893 1893 2926
rect 1914 2913 1917 2996
rect 1922 2923 1925 2956
rect 1930 2933 1933 3003
rect 1826 2833 1845 2836
rect 1754 2656 1757 2736
rect 1762 2733 1781 2736
rect 1786 2793 1797 2796
rect 1810 2793 1813 2806
rect 1762 2723 1765 2733
rect 1786 2726 1789 2793
rect 1818 2743 1821 2766
rect 1778 2723 1789 2726
rect 1754 2653 1761 2656
rect 1690 2583 1693 2606
rect 1682 2533 1685 2546
rect 1714 2523 1717 2606
rect 1758 2596 1761 2653
rect 1802 2623 1805 2736
rect 1818 2703 1821 2726
rect 1826 2716 1829 2833
rect 1938 2826 1941 2926
rect 1946 2913 1949 2936
rect 1954 2903 1957 2976
rect 1970 2836 1973 3003
rect 1978 2983 1981 3116
rect 2026 3113 2029 3136
rect 2034 3123 2037 3136
rect 2042 3123 2045 3153
rect 2050 3093 2053 3136
rect 2066 3113 2069 3146
rect 1986 2953 1989 3016
rect 2002 2993 2005 3006
rect 2010 2976 2013 3016
rect 2018 3003 2021 3076
rect 2002 2973 2013 2976
rect 2026 2973 2029 3016
rect 2034 3003 2037 3056
rect 2074 3023 2077 3206
rect 2082 3133 2085 3213
rect 2090 3193 2093 3206
rect 2082 3016 2085 3126
rect 2090 3106 2093 3166
rect 2154 3156 2157 3233
rect 2170 3223 2181 3226
rect 2170 3193 2173 3206
rect 2178 3183 2181 3206
rect 2098 3123 2101 3136
rect 2114 3123 2117 3156
rect 2154 3153 2181 3156
rect 2186 3153 2189 3216
rect 2202 3163 2205 3206
rect 2210 3186 2213 3216
rect 2234 3196 2237 3263
rect 2258 3203 2261 3246
rect 2234 3193 2245 3196
rect 2210 3183 2229 3186
rect 2090 3103 2101 3106
rect 2098 3026 2101 3103
rect 2130 3053 2133 3126
rect 2146 3123 2149 3136
rect 2162 3116 2165 3136
rect 2170 3133 2173 3146
rect 2178 3136 2181 3153
rect 2178 3133 2185 3136
rect 2146 3113 2165 3116
rect 2146 3036 2149 3113
rect 2170 3096 2173 3116
rect 2042 3003 2045 3016
rect 2058 3013 2069 3016
rect 2074 3013 2085 3016
rect 2090 3023 2101 3026
rect 2122 3033 2149 3036
rect 2162 3093 2173 3096
rect 2066 2993 2069 3006
rect 1966 2833 1973 2836
rect 1938 2823 1957 2826
rect 1842 2783 1845 2806
rect 1890 2793 1893 2816
rect 1834 2723 1837 2736
rect 1842 2723 1845 2736
rect 1850 2733 1853 2756
rect 1858 2723 1861 2766
rect 1922 2753 1925 2816
rect 1930 2803 1933 2816
rect 1938 2763 1941 2816
rect 1954 2793 1957 2806
rect 1966 2786 1969 2833
rect 1986 2813 1989 2936
rect 1994 2903 1997 2926
rect 2002 2916 2005 2973
rect 2074 2966 2077 3013
rect 2090 2996 2093 3023
rect 2090 2993 2101 2996
rect 2042 2963 2077 2966
rect 2018 2933 2029 2936
rect 2002 2913 2013 2916
rect 2018 2913 2021 2926
rect 2026 2856 2029 2926
rect 2042 2906 2045 2963
rect 2042 2903 2053 2906
rect 2018 2853 2029 2856
rect 1966 2783 1973 2786
rect 1986 2783 1989 2806
rect 1970 2766 1973 2783
rect 1970 2763 1981 2766
rect 1826 2713 1853 2716
rect 1850 2656 1853 2713
rect 1906 2686 1909 2736
rect 1906 2683 1917 2686
rect 1846 2653 1853 2656
rect 1770 2603 1773 2616
rect 1834 2613 1837 2626
rect 1758 2593 1773 2596
rect 1706 2456 1709 2476
rect 1706 2453 1713 2456
rect 1666 2383 1677 2386
rect 1610 2213 1613 2306
rect 1618 2213 1629 2216
rect 1634 2213 1637 2226
rect 1618 2193 1621 2206
rect 1626 2183 1629 2206
rect 1610 2003 1613 2116
rect 1618 2106 1621 2136
rect 1626 2123 1629 2146
rect 1618 2103 1625 2106
rect 1622 2036 1625 2103
rect 1618 2033 1625 2036
rect 1618 2013 1621 2033
rect 1634 2006 1637 2156
rect 1610 1896 1613 1986
rect 1618 1903 1621 2006
rect 1626 2003 1637 2006
rect 1642 2003 1645 2266
rect 1650 2203 1653 2236
rect 1650 2123 1653 2146
rect 1650 2013 1653 2026
rect 1626 1933 1629 2003
rect 1634 1923 1637 1996
rect 1658 1956 1661 2226
rect 1666 2056 1669 2383
rect 1682 2333 1685 2396
rect 1690 2383 1693 2416
rect 1710 2376 1713 2453
rect 1722 2406 1725 2526
rect 1730 2523 1749 2526
rect 1730 2506 1733 2523
rect 1730 2503 1741 2506
rect 1754 2503 1757 2536
rect 1762 2533 1765 2566
rect 1770 2526 1773 2593
rect 1802 2583 1805 2606
rect 1778 2533 1781 2556
rect 1770 2523 1805 2526
rect 1826 2523 1829 2606
rect 1846 2586 1849 2653
rect 1846 2583 1853 2586
rect 1738 2436 1741 2503
rect 1730 2433 1741 2436
rect 1730 2413 1733 2433
rect 1738 2406 1741 2416
rect 1722 2403 1741 2406
rect 1706 2373 1713 2376
rect 1674 2103 1677 2236
rect 1682 2143 1685 2206
rect 1690 2153 1693 2256
rect 1698 2133 1701 2316
rect 1706 2146 1709 2373
rect 1722 2333 1733 2336
rect 1714 2313 1717 2326
rect 1746 2323 1749 2406
rect 1754 2393 1757 2426
rect 1762 2386 1765 2416
rect 1778 2403 1781 2416
rect 1762 2383 1773 2386
rect 1714 2223 1749 2226
rect 1714 2213 1717 2223
rect 1722 2173 1725 2216
rect 1730 2183 1733 2206
rect 1738 2193 1741 2216
rect 1746 2203 1749 2223
rect 1706 2143 1717 2146
rect 1682 2123 1701 2126
rect 1706 2106 1709 2136
rect 1698 2103 1709 2106
rect 1666 2053 1677 2056
rect 1666 1963 1669 2046
rect 1658 1953 1669 1956
rect 1626 1913 1653 1916
rect 1610 1893 1617 1896
rect 1614 1836 1617 1893
rect 1614 1833 1621 1836
rect 1602 1783 1605 1816
rect 1618 1813 1621 1833
rect 1594 1773 1605 1776
rect 1610 1773 1613 1806
rect 1602 1733 1605 1773
rect 1626 1753 1629 1913
rect 1634 1803 1637 1836
rect 1610 1733 1621 1736
rect 1586 1703 1589 1726
rect 1602 1723 1613 1726
rect 1618 1663 1621 1733
rect 1626 1723 1637 1726
rect 1626 1646 1629 1723
rect 1634 1703 1637 1716
rect 1586 1643 1629 1646
rect 1578 1623 1581 1636
rect 1578 1606 1581 1616
rect 1586 1613 1589 1643
rect 1602 1633 1629 1636
rect 1602 1613 1605 1633
rect 1578 1603 1597 1606
rect 1594 1536 1597 1603
rect 1586 1533 1597 1536
rect 1586 1476 1589 1533
rect 1586 1473 1597 1476
rect 1546 1423 1565 1426
rect 1538 1133 1541 1396
rect 1538 963 1541 1096
rect 1538 893 1541 916
rect 1546 846 1549 1423
rect 1562 1413 1573 1416
rect 1554 1356 1557 1406
rect 1578 1403 1581 1436
rect 1586 1396 1589 1456
rect 1594 1426 1597 1473
rect 1602 1446 1605 1526
rect 1610 1503 1613 1556
rect 1618 1513 1621 1606
rect 1626 1553 1629 1626
rect 1634 1613 1637 1686
rect 1642 1546 1645 1906
rect 1650 1816 1653 1906
rect 1658 1833 1661 1926
rect 1666 1883 1669 1953
rect 1658 1823 1669 1826
rect 1650 1813 1669 1816
rect 1658 1773 1661 1806
rect 1666 1743 1669 1806
rect 1650 1613 1653 1736
rect 1658 1716 1661 1736
rect 1658 1713 1665 1716
rect 1662 1646 1665 1713
rect 1658 1643 1665 1646
rect 1658 1583 1661 1643
rect 1666 1593 1669 1626
rect 1642 1543 1653 1546
rect 1626 1513 1629 1526
rect 1634 1503 1637 1536
rect 1650 1496 1653 1543
rect 1666 1533 1669 1556
rect 1674 1516 1677 2053
rect 1682 2013 1685 2066
rect 1698 2026 1701 2103
rect 1714 2073 1717 2143
rect 1690 2023 1701 2026
rect 1682 1933 1685 1956
rect 1682 1726 1685 1836
rect 1690 1763 1693 2023
rect 1698 2003 1701 2016
rect 1714 2013 1717 2036
rect 1706 1973 1709 2006
rect 1722 2003 1725 2156
rect 1730 2013 1733 2066
rect 1730 1983 1733 2006
rect 1714 1866 1717 1936
rect 1722 1933 1733 1936
rect 1722 1906 1725 1933
rect 1730 1913 1733 1926
rect 1738 1923 1741 2146
rect 1746 2133 1749 2166
rect 1746 2053 1749 2126
rect 1746 2003 1749 2026
rect 1722 1903 1749 1906
rect 1690 1733 1693 1756
rect 1698 1733 1701 1866
rect 1714 1863 1733 1866
rect 1706 1793 1709 1856
rect 1682 1723 1701 1726
rect 1690 1703 1693 1723
rect 1706 1716 1709 1776
rect 1698 1713 1709 1716
rect 1682 1603 1685 1616
rect 1682 1573 1685 1596
rect 1642 1493 1653 1496
rect 1666 1513 1677 1516
rect 1682 1513 1685 1536
rect 1602 1443 1621 1446
rect 1594 1423 1605 1426
rect 1578 1393 1589 1396
rect 1554 1353 1573 1356
rect 1562 1333 1565 1346
rect 1554 1213 1557 1326
rect 1562 1213 1565 1236
rect 1554 1153 1557 1206
rect 1554 1083 1557 1136
rect 1562 1123 1565 1136
rect 1562 1076 1565 1116
rect 1570 1106 1573 1353
rect 1578 1333 1581 1393
rect 1586 1333 1589 1376
rect 1586 1316 1589 1326
rect 1578 1313 1589 1316
rect 1578 1243 1581 1313
rect 1578 1123 1581 1206
rect 1570 1103 1577 1106
rect 1554 1073 1565 1076
rect 1554 1003 1557 1073
rect 1562 996 1565 1066
rect 1574 1036 1577 1103
rect 1558 993 1565 996
rect 1570 1033 1577 1036
rect 1558 876 1561 993
rect 1502 753 1509 756
rect 1522 843 1549 846
rect 1554 873 1561 876
rect 1522 756 1525 843
rect 1554 836 1557 873
rect 1530 833 1541 836
rect 1546 833 1557 836
rect 1530 803 1533 833
rect 1538 813 1541 826
rect 1546 796 1549 833
rect 1542 793 1549 796
rect 1522 753 1533 756
rect 1482 676 1485 716
rect 1490 693 1493 736
rect 1482 673 1493 676
rect 1442 603 1453 606
rect 1458 603 1469 606
rect 1474 596 1477 646
rect 1490 626 1493 673
rect 1482 623 1493 626
rect 1482 603 1485 623
rect 1502 616 1505 753
rect 1514 623 1517 746
rect 1502 613 1509 616
rect 1522 613 1525 626
rect 1466 593 1477 596
rect 1442 523 1445 536
rect 1458 533 1461 546
rect 1466 526 1469 593
rect 1506 586 1509 613
rect 1482 526 1485 586
rect 1506 583 1513 586
rect 1490 533 1493 566
rect 1426 503 1437 506
rect 1366 433 1373 436
rect 1362 403 1365 416
rect 1370 413 1373 433
rect 1378 316 1381 416
rect 1394 393 1397 406
rect 1402 403 1405 496
rect 1426 436 1429 503
rect 1450 473 1453 526
rect 1462 523 1469 526
rect 1462 466 1465 523
rect 1458 463 1465 466
rect 1426 433 1437 436
rect 1410 323 1413 356
rect 1418 323 1421 336
rect 1426 333 1429 416
rect 1434 316 1437 433
rect 1442 416 1445 436
rect 1442 413 1449 416
rect 1378 313 1413 316
rect 1430 313 1437 316
rect 1378 236 1381 313
rect 1362 233 1381 236
rect 1370 173 1373 226
rect 1386 223 1389 276
rect 1402 196 1405 216
rect 1410 196 1413 216
rect 1418 213 1421 296
rect 1430 246 1433 313
rect 1446 306 1449 413
rect 1442 303 1449 306
rect 1430 243 1437 246
rect 1402 193 1413 196
rect 1426 193 1429 226
rect 1402 176 1405 193
rect 1434 186 1437 243
rect 1394 173 1405 176
rect 1410 183 1437 186
rect 1242 123 1253 126
rect 1258 113 1261 126
rect 1282 113 1285 136
rect 1290 126 1293 136
rect 1290 123 1317 126
rect 1290 93 1293 123
rect 1314 53 1317 123
rect 1322 113 1325 143
rect 1338 126 1341 146
rect 1346 133 1349 166
rect 1354 143 1381 146
rect 1338 123 1373 126
rect 1378 123 1381 143
rect 1394 116 1397 173
rect 1394 113 1405 116
rect 1402 93 1405 113
rect 1410 63 1413 183
rect 1442 173 1445 303
rect 1458 226 1461 463
rect 1474 406 1477 526
rect 1482 523 1493 526
rect 1498 473 1501 576
rect 1482 423 1501 426
rect 1466 403 1477 406
rect 1482 326 1485 366
rect 1490 333 1493 406
rect 1498 383 1501 423
rect 1510 416 1513 583
rect 1522 506 1525 606
rect 1530 573 1533 753
rect 1542 716 1545 793
rect 1542 713 1549 716
rect 1546 693 1549 713
rect 1554 636 1557 806
rect 1562 716 1565 856
rect 1570 783 1573 1033
rect 1578 1003 1581 1016
rect 1578 933 1581 976
rect 1586 896 1589 1306
rect 1594 1203 1597 1336
rect 1602 1323 1605 1423
rect 1618 1346 1621 1416
rect 1626 1363 1629 1406
rect 1634 1353 1637 1406
rect 1618 1343 1625 1346
rect 1610 1306 1613 1336
rect 1602 1303 1613 1306
rect 1602 1203 1605 1303
rect 1622 1296 1625 1343
rect 1618 1293 1625 1296
rect 1634 1293 1637 1326
rect 1618 1236 1621 1293
rect 1618 1233 1637 1236
rect 1618 1223 1637 1226
rect 1618 1216 1621 1223
rect 1610 1213 1621 1216
rect 1602 1123 1605 1186
rect 1610 1063 1613 1146
rect 1594 943 1597 1006
rect 1582 893 1589 896
rect 1582 846 1585 893
rect 1602 886 1605 996
rect 1610 923 1613 1006
rect 1618 953 1621 1206
rect 1626 1076 1629 1216
rect 1634 1113 1637 1223
rect 1626 1073 1637 1076
rect 1626 943 1629 1066
rect 1634 953 1637 1073
rect 1618 916 1621 936
rect 1594 883 1605 886
rect 1582 843 1589 846
rect 1586 823 1589 843
rect 1594 813 1597 883
rect 1610 853 1613 916
rect 1618 913 1625 916
rect 1622 846 1625 913
rect 1618 843 1625 846
rect 1618 826 1621 843
rect 1602 823 1621 826
rect 1570 733 1573 776
rect 1586 726 1589 746
rect 1578 723 1589 726
rect 1594 716 1597 726
rect 1562 713 1597 716
rect 1554 633 1565 636
rect 1538 536 1541 626
rect 1554 613 1557 626
rect 1562 606 1565 633
rect 1546 603 1565 606
rect 1530 533 1541 536
rect 1530 513 1533 533
rect 1538 506 1541 526
rect 1522 503 1541 506
rect 1538 486 1541 503
rect 1530 483 1541 486
rect 1530 426 1533 483
rect 1522 423 1533 426
rect 1510 413 1517 416
rect 1514 403 1517 413
rect 1498 333 1501 366
rect 1514 333 1517 356
rect 1482 323 1493 326
rect 1498 323 1509 326
rect 1458 223 1465 226
rect 1450 183 1453 216
rect 1462 156 1465 223
rect 1474 213 1477 306
rect 1522 273 1525 423
rect 1530 333 1533 416
rect 1538 393 1541 406
rect 1546 396 1549 576
rect 1554 513 1557 546
rect 1562 506 1565 546
rect 1570 533 1573 616
rect 1578 533 1581 546
rect 1578 513 1581 526
rect 1562 503 1577 506
rect 1554 423 1557 436
rect 1562 413 1565 446
rect 1574 436 1577 503
rect 1574 433 1581 436
rect 1546 393 1557 396
rect 1482 193 1485 206
rect 1490 166 1493 216
rect 1498 213 1501 246
rect 1530 223 1533 326
rect 1538 323 1541 366
rect 1554 326 1557 393
rect 1570 366 1573 386
rect 1546 323 1557 326
rect 1566 363 1573 366
rect 1538 203 1541 246
rect 1458 153 1465 156
rect 1482 163 1493 166
rect 1426 76 1429 146
rect 1442 123 1445 136
rect 1458 133 1461 153
rect 1450 116 1453 126
rect 1442 113 1453 116
rect 1442 76 1445 113
rect 1482 103 1485 163
rect 1490 133 1493 156
rect 1530 143 1541 146
rect 1546 133 1549 323
rect 1554 213 1557 306
rect 1566 296 1569 363
rect 1578 306 1581 433
rect 1586 416 1589 456
rect 1594 423 1597 696
rect 1602 643 1605 823
rect 1626 816 1629 826
rect 1610 723 1613 816
rect 1622 813 1629 816
rect 1622 756 1625 813
rect 1634 773 1637 936
rect 1642 863 1645 1493
rect 1666 1446 1669 1513
rect 1666 1443 1677 1446
rect 1658 1406 1661 1426
rect 1658 1403 1665 1406
rect 1650 1333 1653 1396
rect 1662 1346 1665 1403
rect 1674 1386 1677 1443
rect 1682 1413 1685 1426
rect 1674 1383 1685 1386
rect 1662 1343 1669 1346
rect 1666 1326 1669 1343
rect 1650 1203 1653 1256
rect 1658 1223 1661 1326
rect 1666 1323 1677 1326
rect 1682 1316 1685 1383
rect 1678 1313 1685 1316
rect 1650 1143 1653 1196
rect 1658 1123 1661 1216
rect 1666 1116 1669 1266
rect 1678 1236 1681 1313
rect 1650 1113 1669 1116
rect 1674 1233 1681 1236
rect 1650 996 1653 1113
rect 1674 1096 1677 1233
rect 1690 1216 1693 1656
rect 1698 1623 1701 1713
rect 1714 1693 1717 1806
rect 1722 1803 1725 1816
rect 1730 1813 1733 1863
rect 1722 1733 1725 1786
rect 1738 1783 1741 1896
rect 1746 1816 1749 1903
rect 1754 1863 1757 2326
rect 1762 2303 1765 2336
rect 1770 2333 1773 2383
rect 1802 2366 1805 2523
rect 1834 2503 1837 2526
rect 1842 2523 1845 2566
rect 1850 2506 1853 2583
rect 1858 2533 1861 2546
rect 1882 2523 1885 2616
rect 1914 2583 1917 2683
rect 1938 2613 1941 2726
rect 1954 2723 1957 2746
rect 1978 2686 1981 2763
rect 1994 2733 1997 2746
rect 2018 2743 2021 2853
rect 2034 2793 2037 2816
rect 1970 2683 1981 2686
rect 1970 2656 1973 2683
rect 1970 2653 1981 2656
rect 1890 2513 1893 2526
rect 1846 2503 1853 2506
rect 1794 2363 1805 2366
rect 1794 2306 1797 2363
rect 1810 2333 1813 2386
rect 1826 2383 1829 2416
rect 1846 2406 1849 2503
rect 1858 2413 1861 2506
rect 1846 2403 1853 2406
rect 1882 2403 1885 2416
rect 1906 2413 1909 2536
rect 1914 2523 1917 2566
rect 1930 2516 1933 2536
rect 1922 2513 1933 2516
rect 1922 2426 1925 2476
rect 1918 2423 1925 2426
rect 1826 2333 1829 2346
rect 1786 2303 1797 2306
rect 1786 2246 1789 2303
rect 1810 2253 1813 2316
rect 1786 2243 1797 2246
rect 1762 2213 1765 2226
rect 1762 2193 1765 2206
rect 1770 2203 1773 2216
rect 1770 2133 1773 2146
rect 1778 2133 1781 2226
rect 1762 2113 1765 2126
rect 1762 2003 1765 2056
rect 1770 2013 1773 2026
rect 1754 1816 1757 1826
rect 1746 1813 1757 1816
rect 1730 1713 1733 1776
rect 1738 1703 1741 1726
rect 1698 1576 1701 1616
rect 1706 1593 1709 1656
rect 1698 1573 1705 1576
rect 1702 1496 1705 1573
rect 1714 1523 1717 1686
rect 1746 1683 1749 1813
rect 1754 1773 1757 1806
rect 1722 1593 1725 1606
rect 1698 1493 1705 1496
rect 1698 1473 1701 1493
rect 1714 1433 1717 1516
rect 1670 1093 1677 1096
rect 1682 1213 1693 1216
rect 1658 1013 1661 1046
rect 1670 1026 1673 1093
rect 1670 1023 1677 1026
rect 1650 993 1657 996
rect 1618 753 1625 756
rect 1618 723 1621 753
rect 1642 746 1645 856
rect 1654 846 1657 993
rect 1650 843 1657 846
rect 1666 843 1669 1006
rect 1650 806 1653 843
rect 1674 836 1677 1023
rect 1682 1006 1685 1213
rect 1698 1206 1701 1396
rect 1722 1366 1725 1556
rect 1730 1426 1733 1616
rect 1738 1613 1741 1636
rect 1754 1623 1757 1766
rect 1762 1733 1765 1936
rect 1738 1493 1741 1566
rect 1746 1513 1749 1606
rect 1754 1583 1757 1606
rect 1762 1523 1765 1726
rect 1770 1603 1773 1976
rect 1778 1803 1781 2126
rect 1786 2096 1789 2136
rect 1794 2123 1797 2243
rect 1802 2133 1805 2176
rect 1794 2113 1805 2116
rect 1786 2093 1805 2096
rect 1786 1923 1789 2076
rect 1786 1743 1789 1916
rect 1794 1763 1797 2086
rect 1802 2033 1805 2093
rect 1810 2073 1813 2246
rect 1834 2223 1837 2236
rect 1818 2123 1821 2216
rect 1826 2103 1829 2176
rect 1818 2016 1821 2036
rect 1802 1886 1805 2016
rect 1810 2013 1821 2016
rect 1826 2013 1829 2026
rect 1810 1903 1813 1926
rect 1802 1883 1809 1886
rect 1806 1816 1809 1883
rect 1818 1873 1821 2006
rect 1834 1946 1837 2166
rect 1842 2146 1845 2206
rect 1850 2203 1853 2403
rect 1874 2333 1877 2386
rect 1882 2333 1885 2346
rect 1898 2313 1901 2366
rect 1918 2346 1921 2423
rect 1930 2376 1933 2416
rect 1962 2413 1965 2526
rect 1970 2513 1973 2536
rect 1978 2473 1981 2653
rect 1986 2533 1989 2636
rect 2002 2626 2005 2726
rect 2034 2723 2037 2736
rect 2050 2666 2053 2903
rect 2066 2826 2069 2936
rect 2090 2913 2093 2926
rect 2058 2823 2069 2826
rect 2058 2783 2061 2823
rect 2066 2813 2085 2816
rect 2066 2743 2069 2813
rect 2090 2803 2093 2816
rect 2098 2796 2101 2993
rect 2114 2953 2117 3006
rect 2122 3003 2125 3033
rect 2162 3026 2165 3093
rect 2182 3086 2185 3133
rect 2202 3123 2205 3136
rect 2226 3133 2229 3183
rect 2242 3146 2245 3193
rect 2266 3183 2269 3216
rect 2274 3193 2277 3206
rect 2290 3193 2293 3216
rect 2298 3213 2301 3236
rect 2234 3143 2245 3146
rect 2218 3116 2221 3126
rect 2194 3113 2221 3116
rect 2234 3116 2237 3143
rect 2274 3133 2277 3146
rect 2234 3113 2245 3116
rect 2234 3096 2237 3113
rect 2250 3103 2253 3126
rect 2266 3113 2269 3126
rect 2298 3123 2301 3156
rect 2306 3133 2309 3206
rect 2314 3203 2317 3216
rect 2322 3176 2325 3216
rect 2322 3173 2333 3176
rect 2330 3133 2333 3173
rect 2338 3133 2341 3283
rect 2346 3213 2349 3266
rect 2354 3133 2357 3186
rect 2362 3153 2365 3326
rect 2370 3183 2373 3236
rect 2378 3223 2381 3246
rect 2386 3233 2389 3340
rect 2434 3326 2437 3340
rect 2426 3323 2437 3326
rect 2426 3266 2429 3323
rect 2426 3263 2437 3266
rect 2386 3213 2389 3226
rect 2402 3216 2405 3256
rect 2410 3223 2413 3246
rect 2394 3213 2413 3216
rect 2394 3203 2397 3213
rect 2410 3173 2413 3206
rect 2434 3186 2437 3263
rect 2450 3236 2453 3340
rect 2482 3326 2485 3340
rect 2474 3323 2485 3326
rect 2474 3266 2477 3323
rect 2498 3276 2501 3340
rect 2498 3273 2509 3276
rect 2474 3263 2485 3266
rect 2426 3183 2437 3186
rect 2442 3233 2453 3236
rect 2370 3133 2373 3146
rect 2178 3083 2185 3086
rect 2226 3093 2237 3096
rect 2178 3026 2181 3083
rect 2162 3023 2173 3026
rect 2130 2966 2133 3016
rect 2138 3003 2141 3016
rect 2146 2973 2149 3016
rect 2170 3003 2173 3023
rect 2178 3023 2221 3026
rect 2178 3013 2181 3023
rect 2186 3013 2197 3016
rect 2130 2963 2137 2966
rect 2106 2926 2109 2946
rect 2106 2923 2113 2926
rect 2110 2826 2113 2923
rect 2134 2906 2137 2963
rect 2186 2953 2189 3013
rect 2194 2993 2197 3006
rect 2210 2946 2213 3016
rect 2218 3003 2221 3023
rect 2226 2996 2229 3093
rect 2194 2943 2213 2946
rect 2218 2993 2229 2996
rect 2146 2923 2149 2936
rect 2130 2903 2137 2906
rect 2130 2836 2133 2903
rect 2154 2886 2157 2926
rect 2090 2793 2101 2796
rect 2106 2823 2113 2826
rect 2122 2833 2133 2836
rect 2138 2883 2157 2886
rect 2122 2823 2125 2833
rect 2050 2663 2061 2666
rect 2002 2623 2013 2626
rect 1994 2603 1997 2616
rect 1994 2523 1997 2596
rect 2010 2546 2013 2623
rect 2034 2583 2037 2606
rect 2058 2576 2061 2663
rect 2066 2613 2069 2736
rect 2082 2703 2085 2726
rect 2090 2656 2093 2793
rect 2106 2776 2109 2823
rect 2114 2793 2117 2806
rect 2130 2803 2133 2826
rect 2106 2773 2117 2776
rect 2082 2653 2093 2656
rect 2002 2543 2013 2546
rect 2042 2573 2061 2576
rect 2042 2546 2045 2573
rect 2082 2563 2085 2653
rect 2114 2636 2117 2773
rect 2138 2746 2141 2883
rect 2178 2813 2181 2936
rect 2194 2926 2197 2943
rect 2202 2933 2213 2936
rect 2194 2923 2205 2926
rect 2202 2913 2205 2923
rect 2210 2856 2213 2926
rect 2218 2923 2221 2993
rect 2202 2853 2213 2856
rect 2202 2813 2205 2853
rect 2226 2836 2229 2986
rect 2234 2973 2237 3016
rect 2234 2923 2237 2966
rect 2242 2893 2245 3016
rect 2258 3003 2261 3106
rect 2266 3013 2269 3026
rect 2282 3013 2285 3116
rect 2250 2923 2253 2956
rect 2266 2916 2269 3006
rect 2298 2986 2301 3046
rect 2322 3023 2325 3126
rect 2338 3026 2341 3126
rect 2346 3113 2349 3126
rect 2362 3056 2365 3126
rect 2386 3123 2389 3136
rect 2410 3106 2413 3156
rect 2354 3053 2365 3056
rect 2402 3103 2413 3106
rect 2338 3023 2349 3026
rect 2354 3023 2357 3053
rect 2402 3036 2405 3103
rect 2418 3073 2421 3136
rect 2426 3103 2429 3183
rect 2434 3133 2437 3176
rect 2442 3156 2445 3233
rect 2450 3203 2453 3226
rect 2442 3153 2449 3156
rect 2402 3033 2413 3036
rect 2346 3016 2349 3023
rect 2322 2993 2325 3006
rect 2330 2986 2333 3006
rect 2298 2983 2333 2986
rect 2338 2983 2341 3016
rect 2346 3013 2357 3016
rect 2410 3013 2413 3033
rect 2282 2933 2285 2966
rect 2298 2933 2301 2946
rect 2266 2913 2277 2916
rect 2274 2866 2277 2913
rect 2290 2873 2293 2926
rect 2306 2923 2309 2976
rect 2354 2963 2357 3006
rect 2314 2913 2317 2936
rect 2322 2906 2325 2926
rect 2330 2923 2341 2926
rect 2298 2903 2309 2906
rect 2314 2903 2325 2906
rect 2274 2863 2285 2866
rect 2222 2833 2229 2836
rect 2154 2783 2157 2806
rect 2222 2786 2225 2833
rect 2234 2813 2237 2826
rect 2222 2783 2229 2786
rect 2250 2783 2253 2806
rect 2226 2766 2229 2783
rect 2282 2766 2285 2863
rect 2298 2813 2301 2903
rect 2314 2816 2317 2903
rect 2338 2873 2341 2916
rect 2346 2903 2349 2936
rect 2314 2813 2349 2816
rect 2226 2763 2253 2766
rect 2282 2763 2289 2766
rect 2138 2743 2165 2746
rect 2138 2703 2141 2726
rect 2106 2633 2117 2636
rect 2106 2616 2109 2633
rect 2102 2613 2109 2616
rect 2102 2546 2105 2613
rect 2042 2543 2053 2546
rect 2002 2523 2005 2543
rect 1978 2403 1981 2416
rect 1930 2373 1941 2376
rect 1918 2343 1925 2346
rect 1922 2323 1925 2343
rect 1938 2333 1941 2373
rect 1906 2313 1941 2316
rect 1906 2296 1909 2313
rect 1866 2173 1869 2216
rect 1842 2143 1853 2146
rect 1826 1943 1837 1946
rect 1842 1946 1845 2136
rect 1850 2006 1853 2143
rect 1858 2123 1861 2136
rect 1866 2043 1869 2136
rect 1874 2123 1877 2146
rect 1858 2013 1861 2026
rect 1850 2003 1861 2006
rect 1858 1953 1861 2003
rect 1866 1976 1869 2036
rect 1874 2003 1877 2106
rect 1882 2013 1885 2136
rect 1866 1973 1877 1976
rect 1842 1943 1869 1946
rect 1818 1833 1821 1866
rect 1826 1823 1829 1943
rect 1834 1933 1861 1936
rect 1834 1923 1845 1926
rect 1850 1903 1853 1916
rect 1806 1813 1829 1816
rect 1810 1756 1813 1806
rect 1818 1763 1821 1786
rect 1794 1753 1813 1756
rect 1794 1736 1797 1753
rect 1826 1746 1829 1813
rect 1834 1783 1837 1896
rect 1858 1886 1861 1933
rect 1850 1883 1861 1886
rect 1842 1833 1845 1866
rect 1842 1813 1845 1826
rect 1850 1796 1853 1883
rect 1866 1876 1869 1943
rect 1874 1923 1877 1966
rect 1858 1823 1861 1876
rect 1866 1873 1877 1876
rect 1842 1793 1853 1796
rect 1842 1776 1845 1793
rect 1866 1786 1869 1866
rect 1874 1826 1877 1873
rect 1882 1843 1885 1956
rect 1874 1823 1881 1826
rect 1778 1733 1797 1736
rect 1778 1586 1781 1716
rect 1770 1583 1781 1586
rect 1754 1493 1757 1516
rect 1762 1426 1765 1506
rect 1770 1463 1773 1583
rect 1730 1423 1741 1426
rect 1762 1423 1769 1426
rect 1714 1363 1725 1366
rect 1730 1363 1733 1416
rect 1690 1203 1701 1206
rect 1690 1093 1693 1203
rect 1698 1143 1701 1196
rect 1698 1063 1701 1126
rect 1706 1113 1709 1346
rect 1714 1263 1717 1363
rect 1722 1333 1725 1356
rect 1714 1223 1717 1256
rect 1714 1163 1717 1216
rect 1722 1123 1725 1326
rect 1738 1236 1741 1423
rect 1746 1313 1749 1406
rect 1754 1333 1757 1416
rect 1766 1326 1769 1423
rect 1762 1323 1769 1326
rect 1730 1233 1741 1236
rect 1730 1106 1733 1233
rect 1738 1173 1741 1216
rect 1726 1103 1733 1106
rect 1698 1013 1701 1026
rect 1714 1023 1717 1086
rect 1682 1003 1701 1006
rect 1706 1003 1717 1006
rect 1682 923 1685 956
rect 1666 833 1677 836
rect 1658 813 1661 826
rect 1666 813 1669 833
rect 1650 803 1661 806
rect 1634 743 1645 746
rect 1626 723 1629 736
rect 1626 636 1629 686
rect 1602 633 1629 636
rect 1602 603 1605 633
rect 1610 623 1621 626
rect 1626 576 1629 626
rect 1634 603 1637 743
rect 1642 613 1645 736
rect 1658 726 1661 803
rect 1674 743 1677 806
rect 1650 586 1653 726
rect 1658 723 1669 726
rect 1666 646 1669 723
rect 1682 713 1685 916
rect 1690 736 1693 946
rect 1698 866 1701 1003
rect 1726 966 1729 1103
rect 1738 973 1741 1136
rect 1726 963 1733 966
rect 1706 943 1725 946
rect 1706 886 1709 926
rect 1714 893 1717 936
rect 1722 933 1725 943
rect 1722 886 1725 926
rect 1706 883 1725 886
rect 1698 863 1705 866
rect 1702 796 1705 863
rect 1722 823 1725 856
rect 1698 793 1705 796
rect 1698 763 1701 793
rect 1714 776 1717 806
rect 1706 773 1717 776
rect 1690 733 1701 736
rect 1690 696 1693 726
rect 1658 643 1669 646
rect 1686 693 1693 696
rect 1658 613 1661 643
rect 1686 626 1689 693
rect 1698 646 1701 733
rect 1706 703 1709 773
rect 1722 663 1725 796
rect 1698 643 1709 646
rect 1642 583 1653 586
rect 1626 573 1637 576
rect 1618 486 1621 516
rect 1626 493 1629 526
rect 1634 523 1637 573
rect 1642 533 1645 583
rect 1666 576 1669 626
rect 1674 613 1677 626
rect 1686 623 1693 626
rect 1690 603 1693 623
rect 1706 613 1725 616
rect 1666 573 1677 576
rect 1618 483 1629 486
rect 1586 413 1597 416
rect 1586 373 1589 406
rect 1578 303 1585 306
rect 1566 293 1573 296
rect 1570 273 1573 293
rect 1582 236 1585 303
rect 1594 293 1597 413
rect 1602 383 1605 456
rect 1610 423 1621 426
rect 1602 333 1605 376
rect 1610 323 1613 423
rect 1618 333 1621 356
rect 1626 306 1629 483
rect 1634 373 1637 416
rect 1642 333 1645 476
rect 1650 403 1653 516
rect 1658 403 1661 506
rect 1666 366 1669 536
rect 1674 513 1677 573
rect 1682 513 1685 536
rect 1698 533 1701 546
rect 1722 536 1725 606
rect 1714 533 1725 536
rect 1714 516 1717 533
rect 1730 523 1733 963
rect 1738 743 1741 936
rect 1746 913 1749 1236
rect 1754 1213 1757 1226
rect 1754 906 1757 1136
rect 1762 1106 1765 1323
rect 1778 1296 1781 1576
rect 1786 1533 1789 1726
rect 1794 1713 1797 1733
rect 1786 1503 1789 1516
rect 1786 1393 1789 1426
rect 1794 1336 1797 1666
rect 1802 1613 1805 1746
rect 1810 1743 1829 1746
rect 1834 1773 1845 1776
rect 1850 1783 1869 1786
rect 1802 1413 1805 1606
rect 1810 1553 1813 1743
rect 1834 1736 1837 1773
rect 1818 1733 1837 1736
rect 1818 1613 1821 1733
rect 1826 1693 1829 1726
rect 1834 1613 1837 1686
rect 1826 1596 1829 1606
rect 1818 1593 1829 1596
rect 1818 1546 1821 1593
rect 1810 1543 1821 1546
rect 1826 1546 1829 1586
rect 1834 1553 1837 1606
rect 1826 1543 1837 1546
rect 1810 1523 1813 1543
rect 1810 1406 1813 1516
rect 1818 1513 1821 1536
rect 1834 1426 1837 1543
rect 1818 1423 1837 1426
rect 1842 1416 1845 1736
rect 1850 1583 1853 1783
rect 1858 1733 1861 1776
rect 1878 1756 1881 1823
rect 1874 1753 1881 1756
rect 1866 1723 1869 1746
rect 1874 1733 1877 1753
rect 1858 1623 1861 1716
rect 1866 1713 1877 1716
rect 1866 1616 1869 1696
rect 1862 1613 1869 1616
rect 1850 1543 1853 1576
rect 1862 1546 1865 1613
rect 1858 1543 1865 1546
rect 1850 1503 1853 1526
rect 1834 1413 1845 1416
rect 1850 1413 1853 1476
rect 1802 1403 1813 1406
rect 1802 1343 1805 1403
rect 1818 1346 1821 1406
rect 1834 1396 1837 1413
rect 1842 1403 1853 1406
rect 1834 1393 1845 1396
rect 1818 1343 1829 1346
rect 1794 1333 1821 1336
rect 1802 1303 1805 1316
rect 1818 1313 1821 1333
rect 1826 1323 1829 1343
rect 1778 1293 1805 1296
rect 1770 1223 1773 1236
rect 1778 1143 1781 1286
rect 1786 1223 1797 1226
rect 1770 1123 1781 1126
rect 1762 1103 1769 1106
rect 1766 986 1769 1103
rect 1786 1073 1789 1223
rect 1794 1123 1797 1136
rect 1802 1116 1805 1293
rect 1810 1156 1813 1306
rect 1818 1203 1821 1236
rect 1826 1223 1829 1256
rect 1818 1173 1829 1176
rect 1810 1153 1821 1156
rect 1794 1113 1805 1116
rect 1794 1066 1797 1113
rect 1746 903 1757 906
rect 1762 983 1769 986
rect 1778 1063 1797 1066
rect 1746 733 1749 903
rect 1754 803 1757 866
rect 1762 786 1765 983
rect 1770 906 1773 966
rect 1778 923 1781 1063
rect 1786 1013 1789 1026
rect 1794 993 1797 1016
rect 1802 993 1805 1096
rect 1810 1063 1813 1146
rect 1818 1073 1821 1153
rect 1826 1133 1829 1173
rect 1834 1093 1837 1386
rect 1810 1023 1829 1026
rect 1810 993 1813 1023
rect 1786 923 1789 956
rect 1810 916 1813 956
rect 1818 923 1821 1016
rect 1826 1013 1829 1023
rect 1834 1003 1837 1016
rect 1810 913 1821 916
rect 1770 903 1777 906
rect 1774 836 1777 903
rect 1818 876 1821 913
rect 1758 783 1765 786
rect 1770 833 1777 836
rect 1786 873 1821 876
rect 1738 623 1741 716
rect 1746 693 1749 726
rect 1758 656 1761 783
rect 1770 733 1773 833
rect 1778 783 1781 796
rect 1746 653 1761 656
rect 1746 623 1749 653
rect 1770 646 1773 686
rect 1754 643 1773 646
rect 1754 616 1757 643
rect 1742 613 1757 616
rect 1762 633 1773 636
rect 1762 613 1765 633
rect 1778 623 1781 726
rect 1742 546 1745 613
rect 1786 606 1789 873
rect 1802 796 1805 816
rect 1798 793 1805 796
rect 1798 706 1801 793
rect 1798 703 1805 706
rect 1794 623 1797 686
rect 1802 626 1805 703
rect 1810 686 1813 866
rect 1826 826 1829 996
rect 1834 893 1837 906
rect 1822 823 1829 826
rect 1822 766 1825 823
rect 1822 763 1829 766
rect 1818 723 1821 746
rect 1818 693 1821 706
rect 1810 683 1821 686
rect 1802 623 1813 626
rect 1738 543 1745 546
rect 1754 603 1789 606
rect 1794 613 1805 616
rect 1706 513 1717 516
rect 1706 466 1709 513
rect 1730 473 1733 516
rect 1738 513 1741 543
rect 1754 526 1757 603
rect 1794 596 1797 613
rect 1810 596 1813 623
rect 1778 593 1797 596
rect 1802 593 1813 596
rect 1746 523 1757 526
rect 1706 463 1717 466
rect 1674 386 1677 426
rect 1714 406 1717 463
rect 1746 416 1749 523
rect 1770 463 1773 526
rect 1770 423 1773 436
rect 1778 423 1781 576
rect 1786 463 1789 536
rect 1802 503 1805 593
rect 1818 533 1821 666
rect 1810 506 1813 526
rect 1810 503 1821 506
rect 1682 403 1717 406
rect 1722 413 1749 416
rect 1754 413 1789 416
rect 1794 413 1797 496
rect 1810 473 1813 496
rect 1818 456 1821 503
rect 1814 453 1821 456
rect 1722 396 1725 413
rect 1698 393 1725 396
rect 1674 383 1685 386
rect 1666 363 1677 366
rect 1674 306 1677 363
rect 1626 303 1637 306
rect 1610 256 1613 276
rect 1610 253 1617 256
rect 1582 233 1605 236
rect 1562 223 1597 226
rect 1562 203 1565 223
rect 1570 153 1573 216
rect 1578 173 1581 206
rect 1594 193 1597 223
rect 1514 83 1517 116
rect 1554 113 1557 126
rect 1562 123 1565 136
rect 1602 123 1605 233
rect 1614 146 1617 253
rect 1634 246 1637 303
rect 1626 243 1637 246
rect 1658 303 1677 306
rect 1658 246 1661 303
rect 1682 286 1685 383
rect 1698 306 1701 393
rect 1706 316 1709 376
rect 1722 363 1725 393
rect 1746 356 1749 406
rect 1786 396 1789 413
rect 1778 393 1789 396
rect 1746 353 1757 356
rect 1730 343 1749 346
rect 1714 323 1717 336
rect 1722 323 1725 336
rect 1730 323 1733 343
rect 1738 316 1741 336
rect 1746 333 1749 343
rect 1706 313 1741 316
rect 1698 303 1733 306
rect 1746 303 1749 326
rect 1754 323 1757 353
rect 1778 346 1781 393
rect 1778 343 1789 346
rect 1786 323 1789 343
rect 1794 316 1797 406
rect 1802 373 1805 426
rect 1814 356 1817 453
rect 1814 353 1821 356
rect 1818 333 1821 353
rect 1754 313 1789 316
rect 1794 313 1805 316
rect 1658 243 1669 246
rect 1626 203 1629 243
rect 1634 223 1661 226
rect 1610 143 1617 146
rect 1610 126 1613 143
rect 1634 136 1637 223
rect 1658 206 1661 216
rect 1642 203 1661 206
rect 1666 203 1669 243
rect 1626 133 1637 136
rect 1610 123 1621 126
rect 1426 73 1445 76
rect 1586 63 1589 116
rect 1626 93 1629 133
rect 1658 113 1661 136
rect 1634 103 1653 106
rect 1666 63 1669 116
rect 1674 93 1677 286
rect 1682 283 1693 286
rect 1690 216 1693 283
rect 1686 213 1693 216
rect 1686 126 1689 213
rect 1698 133 1701 196
rect 1682 123 1689 126
rect 1706 123 1709 186
rect 1730 126 1733 303
rect 1738 193 1741 226
rect 1746 203 1749 246
rect 1722 123 1733 126
rect 1754 123 1757 313
rect 1802 266 1805 313
rect 1762 213 1765 226
rect 1778 213 1781 266
rect 1794 263 1805 266
rect 1794 243 1797 263
rect 1826 246 1829 763
rect 1834 733 1837 816
rect 1834 513 1837 716
rect 1842 573 1845 1393
rect 1850 1213 1853 1366
rect 1850 1023 1853 1136
rect 1850 993 1853 1006
rect 1850 843 1853 936
rect 1850 733 1853 746
rect 1850 693 1853 726
rect 1850 603 1853 646
rect 1842 543 1845 566
rect 1858 536 1861 1543
rect 1866 1513 1869 1526
rect 1866 1393 1869 1426
rect 1866 1203 1869 1326
rect 1874 1316 1877 1713
rect 1882 1613 1885 1736
rect 1890 1733 1893 2206
rect 1898 2193 1901 2296
rect 1906 2293 1917 2296
rect 1914 2236 1917 2293
rect 1906 2233 1917 2236
rect 1906 2203 1909 2233
rect 1898 2133 1901 2146
rect 1906 2123 1909 2166
rect 1922 2133 1925 2206
rect 1930 2203 1933 2216
rect 1946 2213 1949 2226
rect 1914 2106 1917 2126
rect 1910 2103 1917 2106
rect 1898 1953 1901 2076
rect 1910 2026 1913 2103
rect 1910 2023 1917 2026
rect 1898 1893 1901 1946
rect 1906 1886 1909 2006
rect 1898 1883 1909 1886
rect 1898 1726 1901 1883
rect 1906 1833 1909 1876
rect 1906 1813 1909 1826
rect 1906 1783 1909 1806
rect 1906 1733 1909 1746
rect 1890 1723 1901 1726
rect 1882 1443 1885 1536
rect 1890 1506 1893 1616
rect 1898 1603 1901 1716
rect 1906 1683 1909 1726
rect 1914 1706 1917 2023
rect 1922 2013 1925 2116
rect 1930 2083 1933 2196
rect 1938 2133 1941 2206
rect 1946 2116 1949 2136
rect 1942 2113 1949 2116
rect 1942 2046 1945 2113
rect 1954 2083 1957 2116
rect 1962 2113 1965 2336
rect 2010 2326 2013 2476
rect 2034 2453 2037 2526
rect 2050 2466 2053 2543
rect 2098 2543 2105 2546
rect 2090 2523 2093 2536
rect 2098 2516 2101 2543
rect 2114 2536 2117 2616
rect 2106 2533 2117 2536
rect 2106 2523 2109 2533
rect 2122 2526 2125 2566
rect 2130 2533 2133 2596
rect 2154 2583 2157 2736
rect 2178 2713 2181 2726
rect 2186 2613 2189 2736
rect 2218 2723 2221 2736
rect 2250 2696 2253 2763
rect 2266 2723 2269 2746
rect 2242 2693 2253 2696
rect 2202 2666 2205 2686
rect 2198 2663 2205 2666
rect 2198 2576 2201 2663
rect 2242 2636 2245 2693
rect 2286 2686 2289 2763
rect 2306 2733 2309 2746
rect 2314 2743 2317 2813
rect 2362 2766 2365 3006
rect 2370 2933 2373 3006
rect 2418 3003 2421 3026
rect 2434 3003 2437 3126
rect 2446 3056 2449 3153
rect 2458 3143 2461 3246
rect 2466 3213 2469 3236
rect 2482 3233 2485 3263
rect 2506 3226 2509 3273
rect 2586 3246 2589 3340
rect 2586 3243 2597 3246
rect 2498 3223 2509 3226
rect 2466 3196 2469 3206
rect 2466 3193 2485 3196
rect 2466 3133 2469 3166
rect 2482 3126 2485 3193
rect 2498 3153 2501 3223
rect 2506 3183 2509 3206
rect 2538 3183 2541 3206
rect 2546 3176 2549 3236
rect 2554 3186 2557 3206
rect 2562 3203 2565 3216
rect 2554 3183 2581 3186
rect 2546 3173 2565 3176
rect 2458 3083 2461 3126
rect 2474 3106 2477 3126
rect 2482 3123 2493 3126
rect 2466 3103 2477 3106
rect 2446 3053 2453 3056
rect 2442 3003 2445 3016
rect 2450 3013 2453 3053
rect 2450 3003 2461 3006
rect 2450 2996 2453 3003
rect 2434 2993 2453 2996
rect 2466 2993 2469 3103
rect 2482 3086 2485 3116
rect 2490 3103 2493 3123
rect 2482 3083 2489 3086
rect 2474 3016 2477 3076
rect 2486 3026 2489 3083
rect 2486 3023 2493 3026
rect 2474 3013 2485 3016
rect 2386 2906 2389 2926
rect 2394 2913 2397 2936
rect 2418 2933 2429 2936
rect 2378 2903 2389 2906
rect 2378 2836 2381 2903
rect 2378 2833 2413 2836
rect 2418 2833 2421 2933
rect 2434 2923 2437 2993
rect 2442 2933 2445 2956
rect 2450 2916 2453 2926
rect 2466 2923 2469 2936
rect 2426 2913 2453 2916
rect 2474 2856 2477 3013
rect 2482 2953 2485 3006
rect 2490 2903 2493 3023
rect 2498 2916 2501 3026
rect 2506 2933 2509 3126
rect 2514 3123 2517 3146
rect 2554 3136 2557 3146
rect 2522 3036 2525 3136
rect 2538 3133 2557 3136
rect 2538 3036 2541 3133
rect 2554 3053 2557 3126
rect 2562 3113 2565 3173
rect 2570 3146 2573 3166
rect 2578 3153 2581 3183
rect 2570 3143 2581 3146
rect 2578 3113 2581 3143
rect 2586 3106 2589 3206
rect 2594 3203 2597 3243
rect 2602 3223 2605 3256
rect 2610 3213 2613 3236
rect 2618 3173 2621 3216
rect 2626 3163 2629 3226
rect 2634 3193 2637 3206
rect 2642 3183 2645 3256
rect 2658 3223 2661 3236
rect 2674 3183 2677 3206
rect 2594 3123 2597 3136
rect 2610 3116 2613 3126
rect 2618 3123 2621 3156
rect 2642 3143 2677 3146
rect 2642 3123 2645 3136
rect 2650 3133 2661 3136
rect 2674 3133 2677 3143
rect 2650 3116 2653 3126
rect 2610 3113 2653 3116
rect 2578 3086 2581 3106
rect 2586 3103 2597 3106
rect 2570 3083 2581 3086
rect 2570 3036 2573 3083
rect 2594 3036 2597 3103
rect 2610 3086 2613 3106
rect 2658 3096 2661 3133
rect 2682 3126 2685 3166
rect 2650 3093 2661 3096
rect 2674 3123 2685 3126
rect 2690 3123 2693 3326
rect 2874 3323 2877 3340
rect 2738 3176 2741 3216
rect 2738 3173 2757 3176
rect 2714 3163 2741 3166
rect 2610 3083 2621 3086
rect 2514 3033 2525 3036
rect 2530 3033 2541 3036
rect 2522 2983 2525 3016
rect 2530 2976 2533 3033
rect 2522 2973 2533 2976
rect 2522 2923 2525 2973
rect 2538 2946 2541 3016
rect 2554 3013 2557 3036
rect 2570 3033 2581 3036
rect 2578 3016 2581 3033
rect 2570 3013 2581 3016
rect 2586 3033 2597 3036
rect 2586 3013 2589 3033
rect 2618 3026 2621 3083
rect 2610 3023 2621 3026
rect 2650 3026 2653 3093
rect 2650 3023 2661 3026
rect 2546 2953 2549 3006
rect 2554 2983 2557 3006
rect 2562 2993 2565 3006
rect 2538 2943 2549 2946
rect 2498 2913 2509 2916
rect 2530 2913 2533 2936
rect 2546 2926 2549 2943
rect 2554 2933 2557 2946
rect 2570 2936 2573 3013
rect 2578 2953 2581 3006
rect 2466 2853 2477 2856
rect 2378 2793 2381 2833
rect 2362 2763 2381 2766
rect 2306 2706 2309 2726
rect 2330 2713 2333 2726
rect 2234 2633 2245 2636
rect 2282 2683 2289 2686
rect 2198 2573 2205 2576
rect 2146 2543 2173 2546
rect 2114 2523 2125 2526
rect 2098 2513 2117 2516
rect 2046 2463 2053 2466
rect 2026 2373 2029 2416
rect 2046 2406 2049 2463
rect 2058 2413 2061 2456
rect 2046 2403 2053 2406
rect 2082 2403 2085 2416
rect 1978 2213 1981 2326
rect 2010 2323 2021 2326
rect 1994 2313 2005 2316
rect 1994 2253 1997 2313
rect 2002 2246 2005 2286
rect 1994 2243 2005 2246
rect 1970 2193 1973 2206
rect 1986 2203 1989 2226
rect 1942 2043 1949 2046
rect 1946 2026 1949 2043
rect 1954 2033 1973 2036
rect 1922 1916 1925 1936
rect 1930 1923 1933 2026
rect 1938 2013 1941 2026
rect 1946 2023 1957 2026
rect 1954 2016 1957 2023
rect 1946 1976 1949 2016
rect 1954 2013 1965 2016
rect 1938 1933 1941 1976
rect 1946 1973 1957 1976
rect 1938 1923 1949 1926
rect 1954 1916 1957 1926
rect 1922 1913 1957 1916
rect 1922 1776 1925 1896
rect 1946 1856 1949 1876
rect 1954 1863 1957 1913
rect 1946 1853 1957 1856
rect 1930 1816 1933 1826
rect 1930 1813 1941 1816
rect 1930 1783 1933 1806
rect 1938 1793 1941 1813
rect 1922 1773 1933 1776
rect 1922 1723 1925 1756
rect 1930 1736 1933 1773
rect 1946 1746 1949 1826
rect 1954 1823 1957 1853
rect 1954 1763 1957 1816
rect 1962 1813 1965 2013
rect 1970 1816 1973 2033
rect 1978 2013 1981 2116
rect 1986 2023 1989 2136
rect 1978 1823 1981 1976
rect 1986 1923 1989 1936
rect 1970 1813 1981 1816
rect 1946 1743 1957 1746
rect 1930 1733 1949 1736
rect 1930 1723 1941 1726
rect 1954 1723 1957 1743
rect 1962 1716 1965 1736
rect 1938 1713 1965 1716
rect 1914 1703 1925 1706
rect 1906 1603 1909 1666
rect 1922 1636 1925 1703
rect 1938 1696 1941 1713
rect 1914 1633 1925 1636
rect 1934 1693 1941 1696
rect 1934 1636 1937 1693
rect 1934 1633 1941 1636
rect 1906 1566 1909 1586
rect 1914 1573 1917 1633
rect 1906 1563 1917 1566
rect 1898 1523 1901 1556
rect 1890 1503 1897 1506
rect 1882 1333 1885 1406
rect 1894 1386 1897 1503
rect 1890 1383 1897 1386
rect 1890 1363 1893 1383
rect 1906 1356 1909 1536
rect 1914 1423 1917 1563
rect 1922 1543 1925 1616
rect 1930 1593 1933 1616
rect 1938 1613 1941 1633
rect 1946 1613 1949 1666
rect 1954 1606 1957 1706
rect 1962 1683 1965 1706
rect 1962 1613 1965 1636
rect 1938 1573 1941 1606
rect 1950 1603 1957 1606
rect 1930 1533 1933 1556
rect 1950 1546 1953 1603
rect 1970 1596 1973 1806
rect 1978 1713 1981 1813
rect 1986 1723 1989 1796
rect 1922 1493 1925 1526
rect 1938 1473 1941 1546
rect 1946 1543 1953 1546
rect 1966 1593 1973 1596
rect 1914 1393 1917 1416
rect 1922 1366 1925 1436
rect 1930 1423 1933 1436
rect 1922 1363 1933 1366
rect 1898 1333 1901 1356
rect 1906 1353 1925 1356
rect 1874 1313 1881 1316
rect 1878 1256 1881 1313
rect 1874 1253 1881 1256
rect 1874 1196 1877 1253
rect 1890 1236 1893 1326
rect 1882 1233 1893 1236
rect 1882 1203 1885 1233
rect 1890 1196 1893 1226
rect 1898 1213 1901 1286
rect 1874 1193 1893 1196
rect 1866 1123 1869 1136
rect 1866 1003 1869 1076
rect 1866 923 1869 976
rect 1866 793 1869 836
rect 1866 706 1869 746
rect 1874 726 1877 1193
rect 1882 963 1885 1136
rect 1890 1063 1893 1146
rect 1898 1056 1901 1206
rect 1906 1136 1909 1346
rect 1922 1316 1925 1353
rect 1930 1333 1933 1363
rect 1938 1353 1941 1466
rect 1946 1376 1949 1543
rect 1966 1536 1969 1593
rect 1962 1533 1969 1536
rect 1954 1493 1957 1526
rect 1954 1396 1957 1466
rect 1962 1443 1965 1533
rect 1970 1426 1973 1526
rect 1962 1423 1973 1426
rect 1978 1423 1981 1706
rect 1986 1663 1989 1716
rect 1986 1533 1989 1576
rect 1986 1503 1989 1526
rect 1962 1403 1965 1423
rect 1954 1393 1965 1396
rect 1946 1373 1953 1376
rect 1914 1283 1917 1316
rect 1922 1313 1941 1316
rect 1914 1143 1917 1236
rect 1906 1133 1917 1136
rect 1906 1073 1909 1096
rect 1890 1053 1901 1056
rect 1890 1013 1893 1053
rect 1882 733 1885 916
rect 1874 723 1885 726
rect 1866 703 1873 706
rect 1870 636 1873 703
rect 1866 633 1873 636
rect 1866 613 1869 633
rect 1874 593 1877 606
rect 1842 533 1861 536
rect 1834 403 1837 506
rect 1842 416 1845 533
rect 1882 526 1885 723
rect 1890 716 1893 1006
rect 1898 863 1901 1026
rect 1914 956 1917 1133
rect 1922 1063 1925 1206
rect 1930 1106 1933 1166
rect 1938 1123 1941 1313
rect 1950 1156 1953 1373
rect 1946 1153 1953 1156
rect 1930 1103 1937 1106
rect 1934 1026 1937 1103
rect 1934 1023 1941 1026
rect 1930 973 1933 1016
rect 1914 953 1933 956
rect 1906 933 1909 946
rect 1914 926 1917 946
rect 1906 923 1917 926
rect 1906 823 1909 923
rect 1898 803 1901 816
rect 1914 796 1917 846
rect 1922 833 1925 936
rect 1930 923 1933 953
rect 1938 903 1941 1023
rect 1946 963 1949 1153
rect 1954 896 1957 1136
rect 1962 913 1965 1393
rect 1970 1363 1973 1416
rect 1986 1413 1989 1436
rect 1978 1403 1989 1406
rect 1986 1293 1989 1346
rect 1978 1223 1981 1266
rect 1970 1113 1973 1206
rect 1938 893 1957 896
rect 1938 813 1941 893
rect 1970 843 1973 1076
rect 1978 1013 1981 1216
rect 1986 1153 1989 1206
rect 1986 1123 1989 1146
rect 1994 1106 1997 2243
rect 2018 2236 2021 2323
rect 2034 2293 2037 2336
rect 2042 2333 2045 2346
rect 2050 2283 2053 2403
rect 2066 2333 2069 2376
rect 2082 2333 2085 2346
rect 2002 2233 2021 2236
rect 2002 1973 2005 2233
rect 2010 2203 2013 2226
rect 2010 2093 2013 2146
rect 2018 2133 2021 2166
rect 2026 2123 2029 2196
rect 2034 2106 2037 2216
rect 2050 2203 2053 2216
rect 2066 2213 2069 2246
rect 2058 2183 2061 2206
rect 2030 2103 2037 2106
rect 2010 2013 2013 2076
rect 2030 2036 2033 2103
rect 2042 2063 2045 2176
rect 2074 2146 2077 2316
rect 2058 2143 2077 2146
rect 2058 2056 2061 2143
rect 2074 2113 2077 2136
rect 2082 2133 2085 2256
rect 2090 2123 2093 2326
rect 2114 2323 2117 2513
rect 2138 2456 2141 2526
rect 2146 2513 2149 2543
rect 2162 2526 2165 2536
rect 2170 2533 2173 2543
rect 2178 2526 2181 2546
rect 2154 2493 2157 2526
rect 2162 2523 2181 2526
rect 2202 2523 2205 2573
rect 2218 2503 2221 2526
rect 2234 2456 2237 2633
rect 2242 2533 2245 2546
rect 2258 2523 2261 2626
rect 2266 2583 2269 2616
rect 2274 2563 2277 2616
rect 2282 2546 2285 2683
rect 2298 2616 2301 2706
rect 2306 2703 2317 2706
rect 2314 2646 2317 2703
rect 2306 2643 2317 2646
rect 2306 2623 2309 2643
rect 2298 2613 2325 2616
rect 2290 2593 2293 2606
rect 2314 2573 2317 2606
rect 2282 2543 2333 2546
rect 2266 2516 2269 2526
rect 2282 2523 2285 2536
rect 2290 2516 2293 2536
rect 2306 2526 2309 2543
rect 2266 2513 2293 2516
rect 2302 2523 2309 2526
rect 2138 2453 2165 2456
rect 2234 2453 2245 2456
rect 2050 2053 2061 2056
rect 2030 2033 2037 2036
rect 2018 2013 2021 2026
rect 2034 2016 2037 2033
rect 2042 2023 2045 2036
rect 2026 1996 2029 2016
rect 2034 2013 2045 2016
rect 2018 1993 2029 1996
rect 2010 1883 2013 1916
rect 2002 1813 2005 1826
rect 2010 1823 2013 1876
rect 2018 1796 2021 1993
rect 2026 1923 2029 1976
rect 2034 1893 2037 1986
rect 2002 1793 2021 1796
rect 2002 1593 2005 1793
rect 2026 1766 2029 1886
rect 2042 1856 2045 2006
rect 2050 1926 2053 2053
rect 2058 1933 2061 2016
rect 2066 2013 2069 2036
rect 2074 2003 2077 2106
rect 2082 2013 2085 2056
rect 2066 1933 2069 1986
rect 2050 1923 2061 1926
rect 2050 1883 2053 1916
rect 2058 1866 2061 1923
rect 2066 1893 2069 1926
rect 2034 1853 2045 1856
rect 2054 1863 2061 1866
rect 2034 1813 2037 1853
rect 2042 1823 2045 1846
rect 2054 1766 2057 1863
rect 2026 1763 2037 1766
rect 2054 1763 2061 1766
rect 2010 1713 2013 1756
rect 2018 1723 2021 1736
rect 2026 1733 2029 1756
rect 2034 1716 2037 1763
rect 2050 1733 2053 1746
rect 2058 1736 2061 1763
rect 2066 1743 2069 1886
rect 2074 1843 2077 1996
rect 2090 1956 2093 2036
rect 2082 1953 2093 1956
rect 2082 1896 2085 1953
rect 2090 1923 2093 1946
rect 2098 1933 2101 2206
rect 2114 2203 2117 2226
rect 2122 2213 2125 2336
rect 2130 2333 2133 2416
rect 2162 2413 2165 2453
rect 2242 2436 2245 2453
rect 2242 2433 2249 2436
rect 2178 2403 2181 2416
rect 2130 2293 2133 2316
rect 2146 2296 2149 2386
rect 2146 2293 2153 2296
rect 2138 2266 2141 2286
rect 2134 2263 2141 2266
rect 2134 2176 2137 2263
rect 2150 2236 2153 2293
rect 2162 2273 2165 2396
rect 2226 2353 2229 2416
rect 2246 2346 2249 2433
rect 2258 2413 2261 2506
rect 2302 2446 2305 2523
rect 2314 2456 2317 2526
rect 2330 2523 2333 2543
rect 2338 2533 2341 2636
rect 2354 2603 2357 2736
rect 2346 2523 2349 2586
rect 2378 2576 2381 2763
rect 2386 2723 2389 2806
rect 2394 2713 2397 2816
rect 2402 2803 2405 2826
rect 2410 2813 2413 2833
rect 2450 2813 2453 2836
rect 2426 2783 2429 2806
rect 2466 2796 2469 2853
rect 2466 2793 2477 2796
rect 2474 2773 2477 2793
rect 2434 2683 2437 2726
rect 2466 2723 2469 2736
rect 2386 2603 2389 2616
rect 2394 2603 2397 2616
rect 2402 2576 2405 2616
rect 2410 2603 2413 2636
rect 2362 2573 2405 2576
rect 2314 2453 2357 2456
rect 2302 2443 2309 2446
rect 2274 2403 2277 2416
rect 2306 2396 2309 2443
rect 2302 2393 2309 2396
rect 2178 2333 2189 2336
rect 2178 2273 2181 2326
rect 2186 2316 2189 2333
rect 2186 2313 2193 2316
rect 2190 2236 2193 2313
rect 2202 2303 2205 2316
rect 2226 2293 2229 2336
rect 2234 2333 2237 2346
rect 2242 2343 2249 2346
rect 2242 2243 2245 2343
rect 2258 2333 2261 2356
rect 2266 2333 2269 2346
rect 2258 2306 2261 2326
rect 2254 2303 2261 2306
rect 2146 2233 2153 2236
rect 2186 2233 2193 2236
rect 2146 2183 2149 2233
rect 2134 2173 2141 2176
rect 2106 1906 2109 2116
rect 2098 1903 2109 1906
rect 2082 1893 2109 1896
rect 2082 1883 2101 1886
rect 2058 1733 2069 1736
rect 2074 1733 2077 1816
rect 2082 1803 2085 1883
rect 2042 1723 2053 1726
rect 2034 1713 2045 1716
rect 2010 1653 2013 1706
rect 2034 1626 2037 1656
rect 2010 1623 2037 1626
rect 2010 1603 2013 1623
rect 2002 1433 2005 1586
rect 2018 1573 2021 1616
rect 2026 1593 2029 1616
rect 2034 1603 2037 1623
rect 2026 1523 2029 1556
rect 2026 1506 2029 1516
rect 1990 1103 1997 1106
rect 1978 983 1981 1006
rect 1990 976 1993 1103
rect 1978 973 1993 976
rect 2002 973 2005 1426
rect 2010 1213 2013 1496
rect 2018 1376 2021 1506
rect 2026 1503 2037 1506
rect 2034 1413 2037 1436
rect 2026 1383 2029 1406
rect 2018 1373 2029 1376
rect 2018 1223 2021 1336
rect 1978 923 1981 973
rect 1954 823 1989 826
rect 1930 803 1941 806
rect 1914 793 1921 796
rect 1898 743 1901 776
rect 1906 733 1909 766
rect 1918 736 1921 793
rect 1918 733 1925 736
rect 1890 713 1901 716
rect 1898 646 1901 713
rect 1890 643 1901 646
rect 1890 596 1893 643
rect 1898 613 1901 626
rect 1906 603 1909 626
rect 1890 593 1897 596
rect 1858 523 1885 526
rect 1850 483 1853 506
rect 1858 453 1861 523
rect 1850 443 1869 446
rect 1850 423 1853 443
rect 1866 426 1869 443
rect 1842 413 1853 416
rect 1858 413 1861 426
rect 1866 423 1877 426
rect 1882 423 1885 516
rect 1894 506 1897 593
rect 1914 536 1917 726
rect 1922 696 1925 733
rect 1946 726 1949 816
rect 1994 806 1997 966
rect 2010 963 2013 1206
rect 2018 1023 2021 1136
rect 2026 1016 2029 1373
rect 2042 1343 2045 1713
rect 2050 1663 2053 1723
rect 2058 1653 2061 1726
rect 2066 1653 2069 1733
rect 2082 1646 2085 1766
rect 2090 1733 2093 1816
rect 2098 1803 2101 1866
rect 2106 1736 2109 1893
rect 2114 1856 2117 2136
rect 2122 1883 2125 2076
rect 2130 1933 2133 2136
rect 2138 2073 2141 2173
rect 2146 2026 2149 2116
rect 2154 2076 2157 2206
rect 2162 2193 2165 2216
rect 2170 2186 2173 2206
rect 2178 2203 2181 2226
rect 2170 2183 2181 2186
rect 2170 2166 2173 2183
rect 2162 2163 2173 2166
rect 2162 2123 2165 2163
rect 2186 2156 2189 2233
rect 2170 2153 2189 2156
rect 2154 2073 2165 2076
rect 2154 2033 2157 2056
rect 2138 2023 2149 2026
rect 2138 1913 2141 2023
rect 2154 2016 2157 2026
rect 2162 2023 2165 2073
rect 2146 2013 2157 2016
rect 2170 2013 2173 2153
rect 2194 2146 2197 2216
rect 2234 2203 2237 2226
rect 2242 2213 2245 2236
rect 2254 2216 2257 2303
rect 2250 2213 2257 2216
rect 2186 2143 2197 2146
rect 2178 2103 2181 2126
rect 2186 2073 2189 2143
rect 2194 2083 2197 2126
rect 2114 1853 2125 1856
rect 2098 1733 2109 1736
rect 2098 1723 2101 1733
rect 2050 1643 2101 1646
rect 2050 1613 2053 1643
rect 2050 1593 2053 1606
rect 2058 1543 2061 1616
rect 2066 1603 2069 1626
rect 2074 1583 2077 1636
rect 2082 1576 2085 1636
rect 2066 1573 2085 1576
rect 2050 1473 2053 1516
rect 2058 1503 2061 1536
rect 2050 1403 2053 1446
rect 2058 1386 2061 1496
rect 2066 1486 2069 1573
rect 2082 1516 2085 1536
rect 2074 1513 2085 1516
rect 2074 1493 2077 1513
rect 2066 1483 2077 1486
rect 2066 1423 2069 1446
rect 2074 1416 2077 1483
rect 2054 1383 2061 1386
rect 2066 1413 2077 1416
rect 2082 1413 2085 1506
rect 2090 1476 2093 1576
rect 2098 1536 2101 1643
rect 2106 1593 2109 1726
rect 2114 1716 2117 1846
rect 2122 1763 2125 1853
rect 2130 1756 2133 1846
rect 2138 1773 2141 1816
rect 2146 1813 2149 2013
rect 2154 2003 2173 2006
rect 2154 1813 2157 2003
rect 2178 1996 2181 2026
rect 2194 1996 2197 2026
rect 2162 1993 2181 1996
rect 2186 1993 2197 1996
rect 2202 1996 2205 2166
rect 2210 2123 2213 2136
rect 2226 2123 2229 2136
rect 2202 1993 2213 1996
rect 2146 1763 2149 1806
rect 2122 1723 2125 1756
rect 2130 1753 2149 1756
rect 2162 1753 2165 1993
rect 2170 1923 2181 1926
rect 2186 1923 2189 1993
rect 2194 1933 2197 1986
rect 2202 1923 2205 1946
rect 2170 1903 2173 1923
rect 2170 1813 2173 1886
rect 2170 1753 2173 1806
rect 2178 1803 2181 1896
rect 2130 1726 2133 1736
rect 2130 1723 2141 1726
rect 2114 1713 2125 1716
rect 2098 1533 2109 1536
rect 2098 1493 2101 1526
rect 2090 1473 2097 1476
rect 2034 1263 2037 1336
rect 2054 1326 2057 1383
rect 2042 1306 2045 1326
rect 2054 1323 2061 1326
rect 2042 1303 2049 1306
rect 2046 1256 2049 1303
rect 2042 1253 2049 1256
rect 2034 1113 2037 1206
rect 2042 1166 2045 1253
rect 2042 1163 2053 1166
rect 2022 1013 2029 1016
rect 2034 1013 2037 1106
rect 2042 1093 2045 1156
rect 2050 1123 2053 1163
rect 2058 1123 2061 1323
rect 2066 1233 2069 1413
rect 2082 1366 2085 1406
rect 2074 1363 2085 1366
rect 2066 1163 2069 1226
rect 2066 1093 2069 1106
rect 2074 1076 2077 1363
rect 2082 1246 2085 1356
rect 2094 1346 2097 1473
rect 2106 1403 2109 1533
rect 2090 1343 2097 1346
rect 2090 1323 2093 1343
rect 2106 1333 2109 1356
rect 2114 1276 2117 1686
rect 2122 1613 2125 1713
rect 2130 1663 2133 1716
rect 2138 1653 2141 1723
rect 2146 1713 2149 1753
rect 2154 1693 2157 1736
rect 2130 1583 2133 1616
rect 2138 1603 2141 1616
rect 2130 1566 2133 1576
rect 2146 1573 2149 1606
rect 2130 1563 2149 1566
rect 2122 1486 2125 1526
rect 2130 1493 2133 1536
rect 2146 1533 2149 1563
rect 2154 1526 2157 1606
rect 2138 1523 2157 1526
rect 2154 1486 2157 1516
rect 2122 1483 2157 1486
rect 2122 1413 2125 1426
rect 2130 1403 2133 1426
rect 2122 1363 2125 1396
rect 2138 1356 2141 1466
rect 2146 1383 2149 1436
rect 2122 1353 2141 1356
rect 2122 1323 2125 1353
rect 2154 1343 2157 1426
rect 2130 1313 2133 1336
rect 2138 1283 2141 1326
rect 2146 1293 2149 1336
rect 2114 1273 2149 1276
rect 2082 1243 2101 1246
rect 2082 1226 2085 1243
rect 2082 1223 2089 1226
rect 2086 1156 2089 1223
rect 2098 1213 2101 1243
rect 2098 1196 2101 1206
rect 2106 1203 2109 1256
rect 2114 1213 2133 1216
rect 2122 1196 2125 1206
rect 2130 1203 2133 1213
rect 2098 1193 2125 1196
rect 2086 1153 2117 1156
rect 2022 956 2025 1013
rect 2018 953 2025 956
rect 2002 813 2005 936
rect 2010 893 2013 936
rect 1986 803 1997 806
rect 1942 723 1949 726
rect 1922 693 1933 696
rect 1930 616 1933 693
rect 1942 656 1945 723
rect 1954 683 1957 726
rect 1986 706 1989 803
rect 2002 723 2005 796
rect 1942 653 1949 656
rect 1946 636 1949 653
rect 1962 646 1965 706
rect 1986 703 1997 706
rect 1994 666 1997 703
rect 1986 663 1997 666
rect 1962 643 1973 646
rect 1946 633 1965 636
rect 1922 613 1933 616
rect 1922 593 1925 613
rect 1930 583 1933 596
rect 1890 503 1897 506
rect 1906 533 1917 536
rect 1890 473 1893 503
rect 1874 413 1877 423
rect 1890 413 1893 466
rect 1842 333 1845 346
rect 1850 326 1853 413
rect 1866 376 1869 406
rect 1898 383 1901 486
rect 1866 373 1893 376
rect 1818 243 1829 246
rect 1842 323 1853 326
rect 1842 243 1845 323
rect 1786 196 1789 216
rect 1762 193 1789 196
rect 1794 193 1797 206
rect 1818 176 1821 243
rect 1842 213 1853 216
rect 1866 213 1869 306
rect 1818 173 1829 176
rect 1850 173 1853 213
rect 1810 143 1813 156
rect 1682 103 1685 123
rect 1722 63 1725 123
rect 1762 116 1765 136
rect 1826 133 1829 173
rect 1730 113 1765 116
rect 1770 103 1773 126
rect 1834 113 1837 136
rect 1842 123 1845 166
rect 1858 136 1861 206
rect 1874 203 1877 226
rect 1882 203 1885 246
rect 1890 213 1893 373
rect 1906 333 1909 533
rect 1914 493 1917 526
rect 1922 486 1925 576
rect 1938 533 1941 596
rect 1930 513 1933 526
rect 1946 523 1949 566
rect 1914 483 1925 486
rect 1914 193 1917 483
rect 1922 386 1925 406
rect 1930 403 1933 416
rect 1922 383 1933 386
rect 1930 316 1933 383
rect 1946 323 1949 436
rect 1954 403 1957 616
rect 1962 613 1965 633
rect 1970 603 1973 643
rect 1986 616 1989 663
rect 2002 623 2005 716
rect 2010 646 2013 806
rect 2018 796 2021 953
rect 2042 943 2045 1076
rect 2070 1073 2077 1076
rect 2050 1003 2053 1016
rect 2058 983 2061 1066
rect 2070 996 2073 1073
rect 2082 1013 2085 1126
rect 2098 1123 2101 1136
rect 2098 1063 2101 1116
rect 2106 1103 2109 1146
rect 2114 1036 2117 1153
rect 2122 1103 2125 1166
rect 2114 1033 2121 1036
rect 2130 1033 2133 1126
rect 2138 1123 2141 1206
rect 2070 993 2077 996
rect 2026 813 2029 936
rect 2042 863 2045 936
rect 2034 806 2037 846
rect 2050 813 2053 966
rect 2058 923 2061 976
rect 2074 973 2077 993
rect 2058 896 2061 916
rect 2066 913 2069 946
rect 2058 893 2065 896
rect 2062 826 2065 893
rect 2058 823 2065 826
rect 2026 803 2037 806
rect 2042 803 2053 806
rect 2058 803 2061 823
rect 2018 793 2029 796
rect 2018 716 2021 746
rect 2026 733 2029 793
rect 2034 723 2037 756
rect 2042 733 2053 736
rect 2042 716 2045 726
rect 2018 713 2045 716
rect 2010 643 2029 646
rect 2026 626 2029 643
rect 2050 626 2053 733
rect 2066 703 2069 736
rect 2026 623 2033 626
rect 2050 623 2061 626
rect 1986 613 1997 616
rect 1994 573 1997 613
rect 2002 533 2005 546
rect 1962 433 1965 526
rect 1986 523 1997 526
rect 1970 513 1981 516
rect 1954 316 1957 336
rect 1962 323 1965 426
rect 1970 403 1973 506
rect 1978 486 1981 513
rect 1986 503 1989 523
rect 1978 483 1985 486
rect 1982 396 1985 483
rect 2010 426 2013 526
rect 2002 423 2013 426
rect 1978 393 1985 396
rect 1970 323 1973 336
rect 1978 333 1981 393
rect 1994 316 1997 416
rect 1930 313 1949 316
rect 1954 313 1997 316
rect 1946 306 1949 313
rect 1938 213 1941 306
rect 1946 303 1957 306
rect 1954 286 1957 303
rect 1954 283 1965 286
rect 1962 236 1965 283
rect 2002 273 2005 423
rect 2018 416 2021 606
rect 2030 556 2033 623
rect 2010 413 2021 416
rect 2026 553 2033 556
rect 2010 386 2013 413
rect 2026 403 2029 553
rect 2034 506 2037 536
rect 2042 523 2045 606
rect 2050 603 2053 616
rect 2034 503 2041 506
rect 2038 446 2041 503
rect 2050 483 2053 526
rect 2058 503 2061 623
rect 2066 583 2069 606
rect 2066 533 2069 576
rect 2074 486 2077 966
rect 2082 943 2085 1006
rect 2082 856 2085 936
rect 2090 913 2093 926
rect 2098 866 2101 1016
rect 2106 1013 2109 1026
rect 2106 933 2109 976
rect 2118 966 2121 1033
rect 2138 1023 2141 1036
rect 2130 973 2133 1016
rect 2114 963 2121 966
rect 2098 863 2105 866
rect 2082 853 2093 856
rect 2082 556 2085 816
rect 2090 813 2093 853
rect 2102 806 2105 863
rect 2098 803 2105 806
rect 2090 713 2093 736
rect 2090 623 2093 696
rect 2082 553 2093 556
rect 2082 523 2085 546
rect 2074 483 2081 486
rect 2038 443 2053 446
rect 2034 386 2037 436
rect 2010 383 2021 386
rect 2018 296 2021 383
rect 2010 293 2021 296
rect 2030 383 2037 386
rect 2030 296 2033 383
rect 2030 293 2037 296
rect 1954 233 1965 236
rect 1930 193 1933 206
rect 1946 203 1949 226
rect 1954 213 1957 233
rect 1954 166 1957 206
rect 2002 203 2005 216
rect 1914 163 1957 166
rect 1850 133 1861 136
rect 1874 116 1877 126
rect 1882 123 1885 136
rect 1914 133 1917 163
rect 1938 133 1941 156
rect 1890 116 1893 126
rect 1946 123 1949 136
rect 1954 133 1957 163
rect 1874 113 1893 116
rect 1962 113 1965 136
rect 1994 133 1997 146
rect 2010 133 2013 293
rect 2034 276 2037 293
rect 2042 283 2045 416
rect 2050 413 2053 443
rect 2066 423 2069 476
rect 2078 416 2081 483
rect 2074 413 2081 416
rect 2050 383 2053 406
rect 2058 316 2061 336
rect 2074 326 2077 413
rect 2074 323 2081 326
rect 2054 313 2061 316
rect 2018 193 2021 276
rect 2034 273 2045 276
rect 2026 203 2029 216
rect 2042 203 2045 273
rect 2054 246 2057 313
rect 2066 273 2069 316
rect 2078 266 2081 323
rect 2090 313 2093 553
rect 2098 286 2101 803
rect 2114 746 2117 963
rect 2122 823 2125 946
rect 2138 913 2141 936
rect 2146 923 2149 1273
rect 2154 1196 2157 1326
rect 2162 1203 2165 1716
rect 2170 1523 2173 1746
rect 2178 1586 2181 1756
rect 2186 1683 2189 1866
rect 2186 1593 2189 1626
rect 2178 1583 2189 1586
rect 2170 1423 2173 1446
rect 2154 1193 2165 1196
rect 2154 1053 2157 1166
rect 2162 1036 2165 1193
rect 2170 1093 2173 1346
rect 2178 1146 2181 1536
rect 2186 1506 2189 1583
rect 2194 1516 2197 1816
rect 2202 1813 2205 1856
rect 2202 1773 2205 1806
rect 2202 1633 2205 1696
rect 2210 1623 2213 1993
rect 2218 1863 2221 2056
rect 2226 1986 2229 2096
rect 2234 2013 2237 2136
rect 2242 2133 2245 2166
rect 2250 2116 2253 2213
rect 2258 2183 2261 2206
rect 2246 2113 2253 2116
rect 2246 2046 2249 2113
rect 2246 2043 2253 2046
rect 2250 2023 2253 2043
rect 2258 2033 2261 2126
rect 2266 2093 2269 2316
rect 2274 2213 2277 2276
rect 2274 2083 2277 2206
rect 2282 2133 2285 2206
rect 2290 2163 2293 2376
rect 2302 2346 2305 2393
rect 2302 2343 2309 2346
rect 2306 2323 2309 2343
rect 2282 2093 2285 2126
rect 2242 2013 2253 2016
rect 2258 2003 2261 2016
rect 2266 2013 2269 2076
rect 2274 2003 2277 2026
rect 2282 2013 2285 2036
rect 2226 1983 2269 1986
rect 2218 1793 2221 1816
rect 2218 1723 2221 1766
rect 2226 1716 2229 1966
rect 2234 1903 2237 1936
rect 2242 1933 2261 1936
rect 2234 1763 2237 1806
rect 2242 1753 2245 1933
rect 2250 1893 2253 1926
rect 2258 1913 2261 1933
rect 2266 1896 2269 1983
rect 2274 1923 2277 1986
rect 2274 1903 2277 1916
rect 2262 1893 2269 1896
rect 2262 1826 2265 1893
rect 2274 1836 2277 1896
rect 2282 1863 2285 1936
rect 2290 1903 2293 2136
rect 2298 2106 2301 2246
rect 2306 2193 2309 2226
rect 2314 2213 2317 2386
rect 2322 2333 2325 2416
rect 2354 2413 2357 2453
rect 2330 2333 2333 2346
rect 2362 2326 2365 2573
rect 2386 2526 2389 2566
rect 2402 2533 2413 2536
rect 2386 2523 2413 2526
rect 2426 2493 2429 2646
rect 2442 2613 2445 2656
rect 2434 2533 2437 2586
rect 2450 2566 2453 2616
rect 2442 2563 2453 2566
rect 2442 2523 2445 2563
rect 2378 2403 2381 2416
rect 2402 2366 2405 2416
rect 2394 2363 2405 2366
rect 2394 2333 2397 2363
rect 2362 2323 2381 2326
rect 2322 2296 2325 2316
rect 2322 2293 2333 2296
rect 2330 2236 2333 2293
rect 2326 2233 2333 2236
rect 2306 2123 2309 2156
rect 2298 2103 2305 2106
rect 2314 2103 2317 2206
rect 2326 2156 2329 2233
rect 2338 2183 2341 2216
rect 2346 2206 2349 2246
rect 2354 2213 2357 2236
rect 2346 2203 2357 2206
rect 2362 2203 2365 2226
rect 2370 2203 2373 2216
rect 2322 2153 2329 2156
rect 2302 2036 2305 2103
rect 2298 2033 2305 2036
rect 2298 1903 2301 2033
rect 2306 1993 2309 2016
rect 2306 1923 2309 1966
rect 2314 1896 2317 2006
rect 2290 1893 2317 1896
rect 2274 1833 2285 1836
rect 2262 1823 2269 1826
rect 2234 1733 2237 1746
rect 2250 1736 2253 1806
rect 2242 1733 2253 1736
rect 2218 1613 2221 1716
rect 2226 1713 2233 1716
rect 2230 1636 2233 1713
rect 2242 1703 2245 1726
rect 2258 1723 2261 1806
rect 2226 1633 2233 1636
rect 2202 1526 2205 1536
rect 2210 1533 2213 1586
rect 2202 1523 2213 1526
rect 2194 1513 2205 1516
rect 2186 1503 2197 1506
rect 2186 1413 2189 1436
rect 2186 1306 2189 1406
rect 2194 1363 2197 1503
rect 2202 1476 2205 1513
rect 2210 1493 2213 1516
rect 2202 1473 2209 1476
rect 2206 1356 2209 1473
rect 2218 1403 2221 1576
rect 2202 1353 2209 1356
rect 2202 1323 2205 1353
rect 2218 1336 2221 1346
rect 2210 1333 2221 1336
rect 2210 1313 2213 1333
rect 2218 1306 2221 1326
rect 2186 1303 2221 1306
rect 2186 1293 2197 1296
rect 2186 1153 2189 1293
rect 2194 1233 2205 1236
rect 2194 1163 2197 1206
rect 2202 1153 2205 1233
rect 2210 1156 2213 1236
rect 2218 1223 2221 1256
rect 2218 1163 2221 1216
rect 2226 1213 2229 1633
rect 2234 1523 2237 1616
rect 2242 1583 2245 1606
rect 2258 1603 2261 1636
rect 2234 1423 2237 1446
rect 2234 1383 2237 1416
rect 2234 1323 2237 1366
rect 2234 1226 2237 1256
rect 2242 1233 2245 1576
rect 2258 1533 2261 1596
rect 2250 1493 2253 1526
rect 2266 1456 2269 1823
rect 2274 1793 2277 1816
rect 2274 1633 2277 1756
rect 2274 1613 2277 1626
rect 2274 1523 2277 1546
rect 2266 1453 2277 1456
rect 2250 1253 2253 1426
rect 2258 1403 2261 1416
rect 2258 1333 2261 1356
rect 2266 1343 2269 1446
rect 2274 1326 2277 1453
rect 2282 1396 2285 1833
rect 2290 1813 2293 1893
rect 2290 1573 2293 1736
rect 2290 1443 2293 1536
rect 2290 1403 2293 1436
rect 2298 1403 2301 1886
rect 2306 1813 2309 1886
rect 2322 1816 2325 2153
rect 2330 2123 2333 2136
rect 2338 2123 2341 2136
rect 2346 2123 2349 2176
rect 2354 2116 2357 2203
rect 2362 2133 2373 2136
rect 2346 2113 2357 2116
rect 2330 1923 2333 1996
rect 2338 1983 2341 2016
rect 2346 2013 2349 2113
rect 2362 2096 2365 2126
rect 2378 2123 2381 2323
rect 2386 2293 2389 2316
rect 2402 2243 2405 2336
rect 2386 2106 2389 2126
rect 2358 2093 2365 2096
rect 2382 2103 2389 2106
rect 2358 2026 2361 2093
rect 2358 2023 2365 2026
rect 2346 2003 2357 2006
rect 2338 1906 2341 1936
rect 2346 1923 2349 2003
rect 2354 1923 2357 1986
rect 2362 1956 2365 2023
rect 2370 2013 2373 2076
rect 2382 2036 2385 2103
rect 2382 2033 2389 2036
rect 2394 2033 2397 2136
rect 2410 2116 2413 2206
rect 2426 2166 2429 2286
rect 2434 2266 2437 2326
rect 2450 2323 2453 2446
rect 2458 2413 2461 2606
rect 2466 2546 2469 2616
rect 2466 2543 2477 2546
rect 2466 2513 2469 2536
rect 2474 2523 2477 2543
rect 2482 2506 2485 2616
rect 2474 2503 2485 2506
rect 2490 2503 2493 2896
rect 2506 2846 2509 2913
rect 2498 2843 2509 2846
rect 2538 2906 2541 2926
rect 2546 2923 2557 2926
rect 2554 2913 2557 2923
rect 2562 2913 2565 2936
rect 2570 2933 2581 2936
rect 2570 2906 2573 2926
rect 2538 2903 2573 2906
rect 2498 2796 2501 2843
rect 2506 2813 2509 2826
rect 2498 2793 2505 2796
rect 2502 2706 2505 2793
rect 2514 2723 2517 2806
rect 2530 2793 2533 2836
rect 2538 2796 2541 2903
rect 2578 2843 2581 2933
rect 2610 2856 2613 3023
rect 2658 3006 2661 3023
rect 2666 3013 2669 3026
rect 2674 3013 2677 3123
rect 2690 3023 2693 3116
rect 2698 3106 2701 3126
rect 2698 3103 2705 3106
rect 2702 3036 2705 3103
rect 2698 3033 2705 3036
rect 2650 3003 2661 3006
rect 2650 2993 2653 3003
rect 2690 2996 2693 3006
rect 2658 2993 2693 2996
rect 2634 2923 2637 2946
rect 2674 2936 2677 2956
rect 2674 2933 2681 2936
rect 2678 2886 2681 2933
rect 2690 2913 2693 2926
rect 2674 2883 2681 2886
rect 2674 2856 2677 2883
rect 2602 2853 2613 2856
rect 2670 2853 2677 2856
rect 2554 2813 2573 2816
rect 2538 2793 2549 2796
rect 2554 2733 2557 2813
rect 2586 2776 2589 2806
rect 2602 2803 2605 2853
rect 2650 2813 2653 2826
rect 2670 2806 2673 2853
rect 2670 2803 2677 2806
rect 2674 2783 2677 2803
rect 2586 2773 2605 2776
rect 2562 2753 2581 2756
rect 2502 2703 2509 2706
rect 2506 2606 2509 2703
rect 2498 2603 2509 2606
rect 2530 2603 2533 2726
rect 2546 2653 2549 2726
rect 2562 2723 2565 2753
rect 2578 2733 2581 2753
rect 2578 2613 2581 2726
rect 2602 2723 2605 2773
rect 2658 2686 2661 2726
rect 2634 2683 2661 2686
rect 2634 2636 2637 2683
rect 2498 2586 2501 2603
rect 2498 2583 2525 2586
rect 2474 2403 2477 2416
rect 2498 2396 2501 2583
rect 2506 2516 2509 2526
rect 2522 2523 2525 2583
rect 2530 2533 2533 2586
rect 2610 2546 2613 2616
rect 2594 2543 2613 2546
rect 2594 2533 2597 2543
rect 2506 2513 2557 2516
rect 2490 2393 2501 2396
rect 2474 2316 2477 2336
rect 2490 2326 2493 2393
rect 2506 2333 2509 2416
rect 2554 2413 2557 2513
rect 2594 2453 2597 2526
rect 2602 2523 2605 2536
rect 2618 2533 2621 2636
rect 2630 2633 2637 2636
rect 2630 2586 2633 2633
rect 2650 2603 2653 2616
rect 2682 2596 2685 2846
rect 2690 2733 2693 2816
rect 2698 2783 2701 3033
rect 2706 2833 2709 3016
rect 2714 3003 2717 3163
rect 2722 3133 2725 3156
rect 2738 3133 2741 3163
rect 2754 3133 2757 3173
rect 2770 3153 2773 3216
rect 2778 3203 2781 3226
rect 2794 3213 2813 3216
rect 2826 3213 2829 3236
rect 2850 3233 2853 3246
rect 2866 3216 2869 3256
rect 2810 3206 2813 3213
rect 2762 3123 2765 3146
rect 2786 3133 2789 3166
rect 2802 3136 2805 3206
rect 2810 3203 2821 3206
rect 2842 3203 2845 3216
rect 2858 3213 2869 3216
rect 2818 3183 2821 3196
rect 2826 3193 2837 3196
rect 2834 3163 2837 3193
rect 2858 3166 2861 3213
rect 2874 3173 2877 3226
rect 2858 3163 2869 3166
rect 2866 3146 2869 3163
rect 2882 3146 2885 3216
rect 2906 3203 2909 3236
rect 2914 3223 2949 3226
rect 2986 3223 2989 3256
rect 2994 3243 3029 3246
rect 2994 3216 2997 3243
rect 2914 3146 2917 3216
rect 2970 3213 2997 3216
rect 3018 3213 3021 3236
rect 3026 3213 3029 3243
rect 3042 3213 3061 3216
rect 2954 3193 2957 3206
rect 2962 3153 2965 3206
rect 2866 3143 2873 3146
rect 2882 3143 2965 3146
rect 2802 3133 2813 3136
rect 2714 2933 2717 2946
rect 2714 2826 2717 2926
rect 2722 2906 2725 3056
rect 2770 3013 2773 3026
rect 2738 2933 2741 2976
rect 2762 2923 2765 3006
rect 2778 3003 2781 3126
rect 2810 3123 2813 3133
rect 2842 3096 2845 3136
rect 2834 3093 2845 3096
rect 2834 3036 2837 3093
rect 2834 3033 2845 3036
rect 2786 2923 2789 3016
rect 2826 3006 2829 3016
rect 2810 3003 2829 3006
rect 2826 2993 2837 2996
rect 2826 2953 2829 2986
rect 2818 2923 2821 2946
rect 2722 2903 2741 2906
rect 2826 2903 2829 2916
rect 2834 2903 2837 2993
rect 2706 2823 2717 2826
rect 2706 2753 2709 2823
rect 2714 2746 2717 2816
rect 2722 2803 2725 2826
rect 2730 2813 2733 2846
rect 2706 2743 2717 2746
rect 2722 2743 2725 2786
rect 2738 2783 2741 2903
rect 2842 2836 2845 3033
rect 2850 3003 2853 3056
rect 2858 3023 2861 3126
rect 2870 3086 2873 3143
rect 2882 3103 2885 3136
rect 2890 3123 2893 3136
rect 2898 3113 2901 3143
rect 2906 3113 2909 3126
rect 2870 3083 2877 3086
rect 2874 3036 2877 3083
rect 2938 3053 2941 3136
rect 2962 3123 2965 3143
rect 2970 3133 2973 3146
rect 2978 3133 2981 3186
rect 2986 3173 2989 3206
rect 2994 3133 2997 3206
rect 3042 3203 3045 3213
rect 3034 3133 3037 3146
rect 2962 3046 2965 3116
rect 3034 3103 3037 3116
rect 3042 3096 3045 3196
rect 3050 3163 3053 3206
rect 3058 3183 3061 3213
rect 3106 3156 3109 3326
rect 3258 3253 3301 3256
rect 3106 3153 3117 3156
rect 3082 3143 3109 3146
rect 3050 3133 3069 3136
rect 3050 3123 3053 3133
rect 2866 3033 2877 3036
rect 2866 2966 2869 3033
rect 2898 3023 2901 3046
rect 2946 3043 2965 3046
rect 2946 3023 2949 3043
rect 2858 2963 2869 2966
rect 2850 2923 2853 2936
rect 2858 2846 2861 2963
rect 2866 2913 2869 2956
rect 2858 2843 2869 2846
rect 2842 2833 2861 2836
rect 2746 2753 2749 2806
rect 2754 2756 2757 2816
rect 2762 2803 2765 2826
rect 2770 2766 2773 2816
rect 2778 2783 2781 2806
rect 2818 2803 2821 2816
rect 2842 2813 2845 2826
rect 2858 2786 2861 2833
rect 2850 2783 2861 2786
rect 2770 2763 2785 2766
rect 2754 2753 2773 2756
rect 2770 2743 2773 2753
rect 2698 2733 2717 2736
rect 2698 2613 2701 2733
rect 2722 2723 2725 2736
rect 2730 2723 2733 2736
rect 2770 2713 2773 2726
rect 2782 2716 2785 2763
rect 2818 2756 2821 2766
rect 2794 2753 2821 2756
rect 2794 2723 2797 2753
rect 2802 2743 2813 2746
rect 2782 2713 2789 2716
rect 2786 2646 2789 2713
rect 2786 2643 2793 2646
rect 2678 2593 2685 2596
rect 2630 2583 2637 2586
rect 2570 2403 2573 2416
rect 2514 2333 2517 2346
rect 2490 2323 2517 2326
rect 2450 2303 2453 2316
rect 2474 2313 2509 2316
rect 2434 2263 2445 2266
rect 2442 2213 2445 2263
rect 2498 2246 2501 2266
rect 2450 2166 2453 2246
rect 2498 2243 2505 2246
rect 2474 2223 2477 2236
rect 2458 2203 2469 2206
rect 2426 2163 2445 2166
rect 2450 2163 2461 2166
rect 2426 2123 2429 2136
rect 2410 2113 2421 2116
rect 2378 2003 2381 2016
rect 2362 1953 2373 1956
rect 2334 1903 2341 1906
rect 2334 1836 2337 1903
rect 2346 1853 2349 1906
rect 2334 1833 2341 1836
rect 2314 1813 2325 1816
rect 2306 1623 2309 1796
rect 2314 1776 2317 1813
rect 2322 1783 2325 1806
rect 2314 1773 2325 1776
rect 2314 1603 2317 1766
rect 2306 1533 2309 1576
rect 2306 1493 2309 1526
rect 2306 1396 2309 1446
rect 2282 1393 2293 1396
rect 2282 1343 2285 1386
rect 2258 1323 2277 1326
rect 2258 1233 2261 1323
rect 2234 1223 2245 1226
rect 2242 1213 2245 1223
rect 2266 1213 2269 1316
rect 2282 1266 2285 1336
rect 2274 1263 2285 1266
rect 2210 1153 2221 1156
rect 2178 1143 2213 1146
rect 2178 1103 2181 1126
rect 2158 1033 2165 1036
rect 2158 906 2161 1033
rect 2154 903 2161 906
rect 2114 743 2125 746
rect 2106 683 2109 726
rect 2106 596 2109 646
rect 2114 603 2117 706
rect 2122 663 2125 743
rect 2122 623 2125 636
rect 2106 593 2125 596
rect 2106 513 2109 526
rect 2106 396 2109 426
rect 2114 403 2117 536
rect 2122 526 2125 593
rect 2130 543 2133 866
rect 2154 836 2157 903
rect 2170 863 2173 1056
rect 2186 1033 2189 1106
rect 2194 1103 2197 1116
rect 2202 1106 2205 1136
rect 2210 1123 2213 1143
rect 2202 1103 2209 1106
rect 2178 1023 2189 1026
rect 2194 1023 2197 1096
rect 2206 1026 2209 1103
rect 2206 1023 2213 1026
rect 2194 953 2197 1016
rect 2202 963 2205 1016
rect 2210 936 2213 1023
rect 2218 1013 2221 1153
rect 2218 983 2221 1006
rect 2178 923 2181 936
rect 2194 933 2213 936
rect 2202 916 2205 926
rect 2178 913 2205 916
rect 2210 913 2213 933
rect 2138 823 2141 836
rect 2154 833 2165 836
rect 2146 813 2157 816
rect 2138 746 2141 766
rect 2138 743 2145 746
rect 2142 636 2145 743
rect 2154 733 2157 813
rect 2162 763 2165 833
rect 2170 813 2173 836
rect 2178 803 2189 806
rect 2162 723 2173 726
rect 2154 683 2157 716
rect 2178 693 2181 726
rect 2138 633 2145 636
rect 2138 573 2141 633
rect 2162 623 2165 636
rect 2146 613 2181 616
rect 2186 613 2189 736
rect 2194 733 2197 896
rect 2210 876 2213 896
rect 2206 873 2213 876
rect 2218 873 2221 926
rect 2206 746 2209 873
rect 2206 743 2213 746
rect 2218 743 2221 826
rect 2146 536 2149 606
rect 2178 596 2181 613
rect 2178 593 2189 596
rect 2142 533 2149 536
rect 2162 533 2173 536
rect 2178 533 2181 593
rect 2186 533 2189 586
rect 2122 523 2129 526
rect 2126 446 2129 523
rect 2142 486 2145 533
rect 2154 513 2157 526
rect 2178 523 2189 526
rect 2122 443 2129 446
rect 2138 483 2145 486
rect 2122 423 2125 443
rect 2106 393 2117 396
rect 2106 353 2109 376
rect 2106 333 2109 346
rect 2114 313 2117 393
rect 2122 353 2125 416
rect 2138 406 2141 483
rect 2130 403 2141 406
rect 2122 323 2125 346
rect 2130 323 2133 386
rect 2138 336 2141 403
rect 2146 373 2149 476
rect 2154 403 2157 436
rect 2138 333 2149 336
rect 2162 333 2165 356
rect 2130 313 2141 316
rect 2074 263 2081 266
rect 2090 283 2101 286
rect 2054 243 2061 246
rect 2058 223 2061 243
rect 2050 213 2061 216
rect 2050 173 2053 213
rect 2074 203 2077 263
rect 2090 226 2093 283
rect 2090 223 2101 226
rect 2090 143 2093 206
rect 2098 196 2101 223
rect 2106 213 2109 276
rect 2122 213 2125 246
rect 2146 233 2149 333
rect 2154 213 2157 326
rect 2178 286 2181 523
rect 2186 503 2189 516
rect 2186 413 2189 436
rect 2194 383 2197 666
rect 2202 523 2205 726
rect 2210 663 2213 743
rect 2210 613 2213 626
rect 2218 593 2221 606
rect 2226 576 2229 1206
rect 2234 1133 2237 1206
rect 2242 1116 2245 1156
rect 2238 1113 2245 1116
rect 2238 1046 2241 1113
rect 2250 1103 2253 1206
rect 2258 1163 2261 1206
rect 2274 1156 2277 1263
rect 2266 1153 2277 1156
rect 2238 1043 2245 1046
rect 2234 1013 2237 1026
rect 2242 1006 2245 1043
rect 2250 1013 2253 1056
rect 2234 1003 2245 1006
rect 2234 953 2237 1003
rect 2234 846 2237 946
rect 2242 913 2245 976
rect 2234 843 2245 846
rect 2242 833 2245 843
rect 2222 573 2229 576
rect 2210 503 2213 526
rect 2222 476 2225 573
rect 2234 483 2237 816
rect 2242 716 2245 816
rect 2250 806 2253 1006
rect 2258 953 2261 1136
rect 2266 1023 2269 1153
rect 2266 963 2269 1006
rect 2258 893 2261 946
rect 2266 933 2269 946
rect 2274 926 2277 1146
rect 2282 1073 2285 1256
rect 2282 933 2285 1006
rect 2290 973 2293 1393
rect 2298 1393 2309 1396
rect 2298 1123 2301 1393
rect 2306 1333 2309 1346
rect 2306 1313 2309 1326
rect 2306 1253 2309 1296
rect 2306 1203 2309 1216
rect 2314 1156 2317 1566
rect 2322 1163 2325 1773
rect 2330 1753 2333 1816
rect 2338 1813 2341 1833
rect 2346 1756 2349 1826
rect 2338 1753 2349 1756
rect 2330 1653 2333 1726
rect 2338 1703 2341 1753
rect 2354 1746 2357 1866
rect 2362 1753 2365 1946
rect 2370 1813 2373 1953
rect 2386 1936 2389 2033
rect 2394 2013 2397 2026
rect 2402 2003 2405 2046
rect 2394 1983 2397 1996
rect 2386 1933 2405 1936
rect 2386 1923 2397 1926
rect 2378 1833 2381 1906
rect 2386 1846 2389 1923
rect 2394 1903 2397 1916
rect 2402 1906 2405 1933
rect 2410 1913 2413 2106
rect 2418 2096 2421 2113
rect 2418 2093 2425 2096
rect 2422 2036 2425 2093
rect 2418 2033 2425 2036
rect 2402 1903 2413 1906
rect 2386 1843 2397 1846
rect 2394 1823 2397 1843
rect 2378 1793 2381 1806
rect 2346 1743 2357 1746
rect 2346 1713 2349 1743
rect 2346 1633 2349 1686
rect 2330 1496 2333 1616
rect 2338 1533 2341 1586
rect 2346 1533 2349 1606
rect 2338 1496 2341 1526
rect 2330 1493 2341 1496
rect 2346 1493 2349 1516
rect 2330 1423 2333 1436
rect 2338 1406 2341 1466
rect 2346 1413 2349 1426
rect 2330 1323 2333 1406
rect 2338 1403 2349 1406
rect 2338 1316 2341 1366
rect 2346 1323 2349 1403
rect 2338 1313 2349 1316
rect 2354 1246 2357 1736
rect 2362 1723 2373 1726
rect 2378 1723 2381 1736
rect 2386 1733 2389 1816
rect 2394 1773 2397 1816
rect 2402 1803 2405 1866
rect 2362 1603 2365 1716
rect 2370 1663 2373 1723
rect 2370 1623 2373 1636
rect 2362 1423 2365 1536
rect 2370 1413 2373 1516
rect 2370 1386 2373 1406
rect 2362 1383 2373 1386
rect 2362 1353 2365 1383
rect 2362 1263 2365 1336
rect 2370 1256 2373 1376
rect 2330 1243 2357 1246
rect 2362 1253 2373 1256
rect 2306 1153 2317 1156
rect 2306 1143 2309 1153
rect 2322 1136 2325 1156
rect 2298 1103 2301 1116
rect 2306 1083 2309 1136
rect 2318 1133 2325 1136
rect 2318 1036 2321 1133
rect 2318 1033 2325 1036
rect 2298 983 2301 1006
rect 2314 983 2317 1016
rect 2322 976 2325 1033
rect 2330 1013 2333 1243
rect 2338 1203 2341 1236
rect 2346 1213 2357 1216
rect 2362 1213 2365 1253
rect 2346 1183 2349 1206
rect 2338 1146 2341 1166
rect 2338 1143 2345 1146
rect 2342 1056 2345 1143
rect 2338 1053 2345 1056
rect 2338 1003 2341 1053
rect 2346 996 2349 1036
rect 2314 973 2325 976
rect 2338 993 2349 996
rect 2290 926 2293 956
rect 2266 923 2277 926
rect 2282 923 2293 926
rect 2250 803 2257 806
rect 2254 746 2257 803
rect 2254 743 2261 746
rect 2250 723 2253 736
rect 2258 733 2261 743
rect 2242 713 2253 716
rect 2242 593 2245 666
rect 2222 473 2229 476
rect 2162 213 2165 226
rect 2098 193 2105 196
rect 2102 136 2105 193
rect 2058 133 2077 136
rect 2098 133 2105 136
rect 2034 103 2037 116
rect 2074 113 2077 126
rect 2098 53 2101 133
rect 2114 123 2117 206
rect 2146 123 2149 166
rect 2138 93 2141 116
rect 2154 113 2157 126
rect 2170 86 2173 286
rect 2178 283 2189 286
rect 2186 213 2189 283
rect 2202 203 2205 416
rect 2210 353 2213 416
rect 2226 346 2229 473
rect 2242 403 2245 536
rect 2250 513 2253 713
rect 2266 636 2269 923
rect 2274 823 2277 916
rect 2298 913 2301 946
rect 2306 856 2309 936
rect 2282 853 2309 856
rect 2282 733 2285 853
rect 2314 846 2317 973
rect 2322 933 2325 946
rect 2322 913 2325 926
rect 2330 893 2333 966
rect 2290 843 2317 846
rect 2290 726 2293 843
rect 2330 823 2333 866
rect 2282 723 2293 726
rect 2282 636 2285 723
rect 2298 676 2301 806
rect 2306 783 2309 816
rect 2330 763 2333 806
rect 2338 793 2341 993
rect 2346 823 2349 936
rect 2354 913 2357 1213
rect 2362 1033 2365 1196
rect 2370 1133 2373 1236
rect 2378 1143 2381 1656
rect 2386 1603 2389 1726
rect 2394 1626 2397 1756
rect 2402 1733 2405 1746
rect 2410 1723 2413 1903
rect 2418 1876 2421 2033
rect 2426 1983 2429 2016
rect 2434 2013 2437 2136
rect 2442 2113 2445 2163
rect 2450 2103 2453 2156
rect 2442 2013 2445 2096
rect 2434 1973 2437 2006
rect 2450 1956 2453 2036
rect 2426 1953 2453 1956
rect 2426 1893 2429 1953
rect 2442 1927 2445 1946
rect 2442 1924 2452 1927
rect 2418 1873 2429 1876
rect 2418 1803 2421 1856
rect 2426 1793 2429 1873
rect 2434 1803 2437 1916
rect 2442 1873 2445 1924
rect 2458 1916 2461 2163
rect 2466 2123 2469 2203
rect 2474 2116 2477 2216
rect 2482 2193 2485 2206
rect 2482 2123 2485 2176
rect 2466 2113 2477 2116
rect 2466 1963 2469 2113
rect 2450 1913 2461 1916
rect 2466 1913 2469 1926
rect 2442 1753 2445 1856
rect 2434 1733 2445 1736
rect 2434 1713 2437 1726
rect 2418 1676 2421 1696
rect 2418 1673 2429 1676
rect 2402 1633 2413 1636
rect 2394 1623 2405 1626
rect 2386 1363 2389 1536
rect 2394 1456 2397 1616
rect 2402 1466 2405 1623
rect 2418 1616 2421 1636
rect 2426 1623 2429 1673
rect 2410 1613 2421 1616
rect 2410 1523 2413 1613
rect 2418 1583 2421 1596
rect 2418 1513 2421 1536
rect 2426 1523 2429 1606
rect 2434 1593 2437 1626
rect 2442 1583 2445 1676
rect 2402 1463 2413 1466
rect 2394 1453 2405 1456
rect 2386 1323 2389 1346
rect 2386 1123 2389 1286
rect 2362 906 2365 1016
rect 2370 1013 2373 1066
rect 2394 1036 2397 1446
rect 2402 1403 2405 1453
rect 2410 1443 2413 1463
rect 2410 1373 2413 1416
rect 2418 1406 2421 1476
rect 2434 1443 2437 1506
rect 2442 1493 2445 1516
rect 2418 1403 2429 1406
rect 2410 1333 2413 1346
rect 2426 1333 2429 1403
rect 2434 1333 2437 1386
rect 2442 1363 2445 1456
rect 2402 1316 2405 1326
rect 2418 1323 2429 1326
rect 2402 1313 2421 1316
rect 2402 1303 2413 1306
rect 2418 1303 2421 1313
rect 2402 1113 2405 1266
rect 2378 1033 2397 1036
rect 2370 973 2373 1006
rect 2370 923 2373 966
rect 2358 903 2365 906
rect 2358 836 2361 903
rect 2354 833 2361 836
rect 2306 743 2333 746
rect 2306 733 2309 743
rect 2314 683 2317 736
rect 2330 733 2333 743
rect 2298 673 2317 676
rect 2258 633 2269 636
rect 2274 633 2285 636
rect 2258 503 2261 633
rect 2266 583 2269 616
rect 2274 613 2277 633
rect 2298 623 2301 646
rect 2290 613 2301 616
rect 2290 606 2293 613
rect 2274 603 2293 606
rect 2298 593 2301 606
rect 2306 603 2309 626
rect 2266 543 2285 546
rect 2266 496 2269 543
rect 2274 513 2277 526
rect 2266 493 2273 496
rect 2250 393 2253 406
rect 2258 386 2261 476
rect 2270 396 2273 493
rect 2282 463 2285 536
rect 2290 523 2301 526
rect 2298 503 2301 523
rect 2282 413 2285 436
rect 2298 396 2301 416
rect 2306 413 2309 536
rect 2314 493 2317 673
rect 2270 393 2301 396
rect 2306 393 2309 406
rect 2218 343 2229 346
rect 2250 383 2261 386
rect 2218 303 2221 343
rect 2226 333 2245 336
rect 2250 333 2253 383
rect 2258 333 2261 356
rect 2242 326 2245 333
rect 2234 306 2237 326
rect 2242 323 2253 326
rect 2258 323 2285 326
rect 2242 313 2253 316
rect 2258 306 2261 323
rect 2298 306 2301 393
rect 2314 363 2317 416
rect 2322 333 2325 726
rect 2330 723 2341 726
rect 2346 723 2349 746
rect 2330 563 2333 723
rect 2354 716 2357 833
rect 2370 826 2373 916
rect 2378 906 2381 1033
rect 2386 933 2389 1016
rect 2402 1013 2405 1026
rect 2394 963 2397 1006
rect 2410 986 2413 1303
rect 2426 1293 2429 1323
rect 2442 1276 2445 1356
rect 2450 1313 2453 1896
rect 2458 1883 2461 1906
rect 2474 1856 2477 2106
rect 2490 2093 2493 2216
rect 2502 2176 2505 2243
rect 2498 2173 2505 2176
rect 2498 2116 2501 2173
rect 2514 2156 2517 2323
rect 2506 2153 2517 2156
rect 2506 2123 2509 2153
rect 2514 2123 2517 2136
rect 2498 2113 2509 2116
rect 2466 1853 2477 1856
rect 2458 1746 2461 1826
rect 2466 1823 2469 1836
rect 2466 1773 2469 1816
rect 2474 1783 2477 1836
rect 2458 1743 2469 1746
rect 2458 1713 2461 1736
rect 2466 1693 2469 1743
rect 2474 1713 2477 1726
rect 2458 1653 2469 1656
rect 2458 1586 2461 1653
rect 2466 1623 2477 1626
rect 2482 1623 2485 2026
rect 2490 2013 2493 2076
rect 2490 1916 2493 2006
rect 2498 1923 2501 2086
rect 2506 1963 2509 2113
rect 2522 2106 2525 2136
rect 2518 2103 2525 2106
rect 2518 2036 2521 2103
rect 2518 2033 2525 2036
rect 2490 1913 2509 1916
rect 2490 1813 2493 1913
rect 2514 1906 2517 2016
rect 2502 1903 2517 1906
rect 2502 1836 2505 1903
rect 2498 1833 2505 1836
rect 2498 1813 2501 1833
rect 2514 1806 2517 1896
rect 2498 1793 2501 1806
rect 2506 1803 2517 1806
rect 2466 1613 2469 1623
rect 2490 1616 2493 1756
rect 2498 1716 2501 1776
rect 2506 1743 2509 1803
rect 2522 1743 2525 2033
rect 2530 1993 2533 2256
rect 2554 2213 2557 2326
rect 2594 2316 2597 2336
rect 2602 2333 2605 2376
rect 2610 2326 2613 2526
rect 2626 2513 2629 2536
rect 2634 2523 2637 2583
rect 2678 2546 2681 2593
rect 2678 2543 2685 2546
rect 2682 2526 2685 2543
rect 2690 2533 2693 2586
rect 2738 2533 2741 2616
rect 2762 2603 2765 2616
rect 2790 2596 2793 2643
rect 2802 2613 2805 2736
rect 2810 2716 2813 2743
rect 2818 2723 2821 2753
rect 2826 2733 2829 2776
rect 2826 2716 2829 2726
rect 2810 2713 2829 2716
rect 2850 2676 2853 2783
rect 2866 2683 2869 2843
rect 2898 2823 2901 2936
rect 2922 2923 2925 3006
rect 2930 2903 2933 3006
rect 2946 2993 2949 3016
rect 2962 3013 2965 3043
rect 3034 3093 3045 3096
rect 3034 3023 3037 3093
rect 3042 3023 3069 3026
rect 3042 3013 3045 3023
rect 3082 3016 3085 3143
rect 3090 3113 3093 3136
rect 3098 3116 3101 3126
rect 3106 3123 3109 3143
rect 3114 3126 3117 3153
rect 3130 3133 3133 3216
rect 3186 3176 3189 3216
rect 3258 3213 3261 3253
rect 3178 3173 3189 3176
rect 3178 3133 3181 3173
rect 3114 3123 3133 3126
rect 3098 3113 3125 3116
rect 3130 3066 3133 3123
rect 3178 3116 3181 3126
rect 3186 3123 3189 3136
rect 3194 3116 3197 3126
rect 3178 3113 3197 3116
rect 2954 3003 2973 3006
rect 2970 2983 2973 3003
rect 3034 2993 3037 3006
rect 3050 3003 3053 3016
rect 3066 3013 3085 3016
rect 3114 3063 3133 3066
rect 3018 2933 3021 2956
rect 3026 2943 3029 2966
rect 3034 2933 3037 2946
rect 2898 2773 2901 2816
rect 2914 2803 2917 2896
rect 2978 2893 2981 2926
rect 3002 2923 3053 2926
rect 3058 2906 3061 2996
rect 3050 2903 3061 2906
rect 3050 2836 3053 2903
rect 3034 2833 3053 2836
rect 2922 2813 2925 2826
rect 2962 2823 2981 2826
rect 2930 2813 2941 2816
rect 2962 2813 2965 2823
rect 2890 2696 2893 2736
rect 2930 2723 2933 2813
rect 2946 2763 2949 2806
rect 2970 2733 2973 2816
rect 2978 2813 2981 2823
rect 2994 2803 2997 2826
rect 3034 2803 3037 2833
rect 3042 2813 3045 2826
rect 3058 2766 3061 2816
rect 3066 2793 3069 3013
rect 3074 2923 3077 3006
rect 3098 2976 3101 3006
rect 3114 3003 3117 3063
rect 3138 2976 3141 3016
rect 3194 2993 3197 3016
rect 3098 2973 3141 2976
rect 3082 2913 3085 2926
rect 3090 2826 3093 2966
rect 3122 2913 3125 2926
rect 3130 2896 3133 2936
rect 3154 2923 3157 2946
rect 3162 2933 3165 2986
rect 3170 2923 3173 2946
rect 3146 2913 3157 2916
rect 3130 2893 3149 2896
rect 3146 2846 3149 2893
rect 3194 2866 3197 2976
rect 3202 2933 3205 3006
rect 3194 2863 3201 2866
rect 3146 2843 3189 2846
rect 3090 2823 3101 2826
rect 3146 2823 3149 2843
rect 3154 2833 3181 2836
rect 3050 2763 3061 2766
rect 2882 2693 2893 2696
rect 2850 2673 2861 2676
rect 2858 2616 2861 2673
rect 2882 2636 2885 2693
rect 2882 2633 2893 2636
rect 2786 2593 2793 2596
rect 2786 2576 2789 2593
rect 2762 2573 2797 2576
rect 2754 2533 2757 2546
rect 2666 2513 2669 2526
rect 2682 2523 2709 2526
rect 2618 2376 2621 2416
rect 2650 2413 2653 2456
rect 2674 2403 2677 2416
rect 2698 2386 2701 2406
rect 2694 2383 2701 2386
rect 2618 2373 2629 2376
rect 2626 2333 2629 2373
rect 2674 2333 2677 2356
rect 2682 2333 2685 2376
rect 2610 2323 2637 2326
rect 2570 2303 2573 2316
rect 2594 2313 2629 2316
rect 2562 2223 2581 2226
rect 2562 2206 2565 2216
rect 2546 2203 2565 2206
rect 2570 2203 2573 2216
rect 2546 2126 2549 2136
rect 2538 2123 2549 2126
rect 2530 1863 2533 1906
rect 2538 1856 2541 2123
rect 2546 1913 2549 2116
rect 2554 2103 2557 2136
rect 2562 2123 2565 2176
rect 2578 2116 2581 2223
rect 2586 2203 2589 2226
rect 2594 2203 2597 2216
rect 2570 2113 2581 2116
rect 2554 2013 2565 2016
rect 2570 2013 2573 2113
rect 2554 1983 2557 2013
rect 2554 1923 2557 1976
rect 2562 1936 2565 2006
rect 2562 1933 2573 1936
rect 2578 1933 2581 2056
rect 2586 1996 2589 2046
rect 2594 2013 2597 2146
rect 2602 2106 2605 2136
rect 2610 2123 2613 2146
rect 2618 2133 2621 2216
rect 2634 2213 2637 2323
rect 2642 2313 2645 2326
rect 2694 2316 2697 2383
rect 2690 2313 2697 2316
rect 2666 2223 2669 2246
rect 2690 2236 2693 2313
rect 2690 2233 2701 2236
rect 2658 2213 2669 2216
rect 2642 2153 2645 2206
rect 2602 2103 2609 2106
rect 2606 2026 2609 2103
rect 2602 2023 2609 2026
rect 2602 2003 2605 2023
rect 2618 2013 2621 2086
rect 2626 2053 2629 2126
rect 2634 2103 2637 2136
rect 2586 1993 2605 1996
rect 2570 1926 2573 1933
rect 2562 1916 2565 1926
rect 2570 1923 2581 1926
rect 2554 1913 2565 1916
rect 2538 1853 2549 1856
rect 2530 1803 2533 1816
rect 2506 1723 2525 1726
rect 2498 1713 2513 1716
rect 2474 1613 2493 1616
rect 2498 1613 2501 1706
rect 2458 1583 2469 1586
rect 2458 1413 2461 1576
rect 2466 1413 2469 1583
rect 2458 1343 2461 1396
rect 2466 1336 2469 1406
rect 2458 1333 2469 1336
rect 2426 1273 2445 1276
rect 2418 1213 2421 1236
rect 2426 1203 2429 1273
rect 2434 1193 2437 1266
rect 2418 1103 2421 1136
rect 2426 1076 2429 1096
rect 2422 1073 2429 1076
rect 2422 996 2425 1073
rect 2434 1063 2437 1136
rect 2422 993 2429 996
rect 2406 983 2413 986
rect 2406 936 2409 983
rect 2406 933 2413 936
rect 2394 916 2397 926
rect 2394 913 2405 916
rect 2378 903 2389 906
rect 2386 846 2389 903
rect 2386 843 2397 846
rect 2370 823 2377 826
rect 2342 713 2357 716
rect 2342 656 2345 713
rect 2338 653 2345 656
rect 2330 326 2333 546
rect 2234 303 2261 306
rect 2290 303 2301 306
rect 2314 323 2333 326
rect 2218 206 2221 226
rect 2218 203 2229 206
rect 2178 113 2181 146
rect 2186 113 2189 126
rect 2234 123 2237 256
rect 2290 236 2293 303
rect 2290 233 2301 236
rect 2186 86 2189 106
rect 2170 83 2189 86
rect 2242 83 2245 216
rect 2250 166 2253 206
rect 2258 193 2261 216
rect 2298 213 2301 233
rect 2314 213 2317 323
rect 2322 313 2333 316
rect 2330 213 2333 313
rect 2338 206 2341 653
rect 2346 573 2349 636
rect 2354 566 2357 706
rect 2346 563 2357 566
rect 2346 433 2349 563
rect 2362 533 2365 816
rect 2374 756 2377 823
rect 2370 753 2377 756
rect 2370 643 2373 753
rect 2378 626 2381 736
rect 2386 733 2389 826
rect 2386 633 2389 646
rect 2370 616 2373 626
rect 2378 623 2389 626
rect 2370 613 2377 616
rect 2386 613 2389 623
rect 2354 523 2365 526
rect 2362 516 2365 523
rect 2374 516 2377 613
rect 2386 533 2389 566
rect 2362 513 2377 516
rect 2370 423 2381 426
rect 2386 423 2389 486
rect 2394 416 2397 843
rect 2402 806 2405 913
rect 2410 906 2413 933
rect 2418 923 2421 976
rect 2426 933 2429 993
rect 2434 943 2437 1026
rect 2410 903 2421 906
rect 2418 836 2421 903
rect 2410 833 2421 836
rect 2434 833 2437 936
rect 2410 813 2413 833
rect 2442 826 2445 1256
rect 2450 1106 2453 1236
rect 2458 1203 2461 1333
rect 2474 1256 2477 1613
rect 2482 1526 2485 1606
rect 2490 1593 2493 1606
rect 2490 1533 2493 1576
rect 2482 1523 2493 1526
rect 2498 1523 2501 1606
rect 2510 1596 2513 1713
rect 2522 1603 2525 1716
rect 2510 1593 2517 1596
rect 2506 1533 2509 1576
rect 2482 1333 2485 1516
rect 2482 1313 2485 1326
rect 2466 1253 2477 1256
rect 2482 1236 2485 1256
rect 2478 1233 2485 1236
rect 2466 1203 2469 1226
rect 2478 1166 2481 1233
rect 2490 1213 2493 1523
rect 2506 1516 2509 1526
rect 2514 1523 2517 1593
rect 2522 1546 2525 1586
rect 2530 1553 2533 1736
rect 2522 1543 2533 1546
rect 2506 1513 2517 1516
rect 2498 1416 2501 1446
rect 2498 1413 2509 1416
rect 2498 1393 2509 1396
rect 2498 1383 2501 1393
rect 2514 1386 2517 1513
rect 2506 1383 2517 1386
rect 2458 1123 2461 1146
rect 2466 1133 2469 1166
rect 2478 1163 2485 1166
rect 2474 1133 2477 1146
rect 2482 1126 2485 1163
rect 2490 1143 2493 1206
rect 2450 1103 2457 1106
rect 2454 1036 2457 1103
rect 2434 823 2445 826
rect 2450 1033 2457 1036
rect 2402 803 2413 806
rect 2426 796 2429 816
rect 2410 793 2429 796
rect 2402 723 2405 766
rect 2402 563 2405 626
rect 2402 533 2405 556
rect 2354 413 2397 416
rect 2346 213 2349 386
rect 2250 163 2261 166
rect 2258 133 2261 163
rect 2282 123 2285 206
rect 2298 123 2301 206
rect 2322 203 2341 206
rect 2306 116 2309 136
rect 2346 123 2349 206
rect 2274 113 2309 116
rect 2354 113 2357 413
rect 2402 406 2405 526
rect 2410 503 2413 756
rect 2418 733 2421 746
rect 2418 683 2421 726
rect 2426 706 2429 766
rect 2434 723 2437 823
rect 2450 803 2453 1033
rect 2458 996 2461 1016
rect 2466 1003 2469 1126
rect 2474 1013 2477 1126
rect 2482 1123 2489 1126
rect 2486 1036 2489 1123
rect 2482 1033 2489 1036
rect 2474 996 2477 1006
rect 2458 993 2477 996
rect 2458 893 2461 916
rect 2466 863 2469 936
rect 2474 846 2477 946
rect 2482 906 2485 1033
rect 2490 983 2493 1016
rect 2490 923 2493 946
rect 2498 933 2501 1316
rect 2506 1106 2509 1383
rect 2514 1283 2517 1356
rect 2514 1223 2517 1256
rect 2514 1123 2517 1206
rect 2522 1203 2525 1526
rect 2522 1143 2525 1196
rect 2506 1103 2517 1106
rect 2514 1026 2517 1103
rect 2506 1023 2517 1026
rect 2482 903 2489 906
rect 2486 846 2489 903
rect 2470 843 2477 846
rect 2482 843 2489 846
rect 2458 796 2461 836
rect 2450 793 2461 796
rect 2426 703 2437 706
rect 2450 703 2453 793
rect 2418 633 2421 646
rect 2434 636 2437 703
rect 2426 633 2437 636
rect 2418 573 2421 626
rect 2426 566 2429 633
rect 2458 623 2461 786
rect 2470 766 2473 843
rect 2470 763 2477 766
rect 2474 743 2477 763
rect 2466 723 2477 726
rect 2418 563 2429 566
rect 2362 403 2405 406
rect 2410 403 2413 466
rect 2418 443 2421 563
rect 2442 533 2445 616
rect 2466 613 2469 723
rect 2426 513 2429 526
rect 2458 523 2461 576
rect 2362 296 2365 403
rect 2386 343 2421 346
rect 2386 333 2389 343
rect 2394 316 2397 326
rect 2370 313 2397 316
rect 2362 293 2373 296
rect 2370 196 2373 293
rect 2362 193 2373 196
rect 2362 173 2365 193
rect 2370 116 2373 136
rect 2378 123 2381 136
rect 2386 133 2389 266
rect 2410 253 2413 336
rect 2402 223 2405 236
rect 2410 233 2413 246
rect 2402 173 2405 216
rect 2418 156 2421 343
rect 2426 263 2429 416
rect 2426 223 2429 236
rect 2418 153 2429 156
rect 2386 123 2397 126
rect 2402 116 2405 136
rect 2426 123 2429 153
rect 2434 133 2437 506
rect 2442 493 2445 516
rect 2442 403 2445 456
rect 2442 233 2445 376
rect 2450 333 2453 516
rect 2458 423 2461 486
rect 2466 416 2469 536
rect 2458 413 2469 416
rect 2458 336 2461 413
rect 2474 383 2477 626
rect 2482 576 2485 843
rect 2498 826 2501 926
rect 2490 823 2501 826
rect 2490 783 2493 823
rect 2498 803 2501 816
rect 2490 663 2493 746
rect 2498 723 2501 756
rect 2506 636 2509 1023
rect 2514 1003 2525 1006
rect 2514 923 2517 1003
rect 2522 933 2525 946
rect 2514 816 2517 856
rect 2514 813 2525 816
rect 2514 716 2517 806
rect 2522 733 2525 813
rect 2530 763 2533 1543
rect 2538 1403 2541 1836
rect 2546 1713 2549 1853
rect 2562 1833 2565 1906
rect 2570 1883 2573 1916
rect 2578 1873 2581 1923
rect 2578 1803 2581 1826
rect 2562 1756 2565 1776
rect 2578 1763 2581 1796
rect 2546 1416 2549 1706
rect 2554 1613 2557 1756
rect 2562 1753 2581 1756
rect 2562 1696 2565 1726
rect 2578 1713 2581 1753
rect 2562 1693 2581 1696
rect 2562 1623 2565 1656
rect 2562 1546 2565 1606
rect 2570 1553 2573 1646
rect 2586 1616 2589 1966
rect 2594 1883 2597 1986
rect 2594 1753 2597 1816
rect 2594 1703 2597 1726
rect 2582 1613 2589 1616
rect 2582 1556 2585 1613
rect 2594 1593 2597 1606
rect 2582 1553 2589 1556
rect 2554 1543 2565 1546
rect 2554 1426 2557 1543
rect 2562 1533 2581 1536
rect 2562 1493 2565 1533
rect 2578 1483 2581 1516
rect 2586 1513 2589 1553
rect 2594 1523 2597 1576
rect 2602 1506 2605 1993
rect 2610 1983 2613 2006
rect 2610 1893 2613 1936
rect 2626 1876 2629 1976
rect 2610 1813 2613 1876
rect 2626 1873 2637 1876
rect 2610 1793 2613 1806
rect 2618 1803 2621 1826
rect 2610 1693 2613 1716
rect 2610 1533 2613 1686
rect 2618 1663 2621 1796
rect 2626 1596 2629 1866
rect 2622 1593 2629 1596
rect 2622 1506 2625 1593
rect 2634 1573 2637 1873
rect 2642 1826 2645 2136
rect 2650 2023 2653 2186
rect 2650 2003 2653 2016
rect 2658 2013 2661 2213
rect 2666 2136 2669 2206
rect 2674 2196 2677 2206
rect 2690 2196 2693 2216
rect 2674 2193 2693 2196
rect 2698 2186 2701 2233
rect 2706 2213 2709 2523
rect 2714 2316 2717 2436
rect 2738 2433 2741 2526
rect 2762 2523 2765 2573
rect 2770 2533 2773 2566
rect 2722 2333 2725 2416
rect 2754 2413 2757 2516
rect 2794 2446 2797 2573
rect 2842 2546 2845 2616
rect 2858 2613 2865 2616
rect 2850 2593 2853 2606
rect 2826 2543 2845 2546
rect 2826 2533 2829 2543
rect 2826 2473 2829 2526
rect 2834 2493 2837 2536
rect 2850 2533 2853 2566
rect 2862 2546 2865 2613
rect 2858 2543 2865 2546
rect 2858 2526 2861 2543
rect 2842 2523 2861 2526
rect 2874 2523 2877 2606
rect 2882 2563 2885 2616
rect 2890 2613 2893 2633
rect 2898 2556 2901 2686
rect 2906 2603 2909 2636
rect 2922 2613 2925 2696
rect 2970 2693 2973 2726
rect 2890 2553 2901 2556
rect 2794 2443 2805 2446
rect 2842 2443 2845 2523
rect 2890 2506 2893 2553
rect 2906 2533 2909 2576
rect 2946 2546 2949 2566
rect 2942 2543 2949 2546
rect 2890 2503 2909 2506
rect 2770 2403 2773 2416
rect 2802 2396 2805 2443
rect 2842 2416 2845 2436
rect 2906 2426 2909 2503
rect 2930 2456 2933 2526
rect 2942 2476 2945 2543
rect 2942 2473 2949 2476
rect 2930 2453 2937 2456
rect 2898 2423 2909 2426
rect 2714 2313 2721 2316
rect 2718 2196 2721 2313
rect 2690 2183 2701 2186
rect 2714 2193 2721 2196
rect 2666 2133 2681 2136
rect 2666 2053 2669 2126
rect 2678 2066 2681 2133
rect 2690 2083 2693 2183
rect 2714 2176 2717 2193
rect 2698 2173 2717 2176
rect 2678 2063 2685 2066
rect 2682 2023 2685 2063
rect 2698 2023 2701 2173
rect 2706 2123 2709 2136
rect 2714 2026 2717 2136
rect 2722 2123 2725 2146
rect 2706 2023 2717 2026
rect 2706 2006 2709 2023
rect 2666 1973 2669 2006
rect 2682 2003 2709 2006
rect 2666 1943 2677 1946
rect 2666 1933 2669 1943
rect 2650 1913 2653 1926
rect 2666 1913 2669 1926
rect 2674 1906 2677 1936
rect 2658 1903 2677 1906
rect 2682 1853 2685 2003
rect 2642 1823 2677 1826
rect 2598 1503 2605 1506
rect 2618 1503 2625 1506
rect 2598 1446 2601 1503
rect 2618 1486 2621 1503
rect 2610 1483 2621 1486
rect 2598 1443 2605 1446
rect 2554 1423 2597 1426
rect 2546 1413 2565 1416
rect 2562 1383 2565 1413
rect 2570 1373 2573 1416
rect 2594 1413 2597 1423
rect 2538 1303 2541 1366
rect 2594 1356 2597 1396
rect 2546 1353 2597 1356
rect 2546 1333 2549 1353
rect 2562 1333 2565 1346
rect 2602 1336 2605 1443
rect 2610 1346 2613 1483
rect 2618 1403 2621 1456
rect 2626 1353 2629 1416
rect 2610 1343 2621 1346
rect 2546 1246 2549 1326
rect 2554 1293 2557 1326
rect 2546 1243 2557 1246
rect 2570 1243 2573 1336
rect 2594 1333 2605 1336
rect 2578 1303 2581 1326
rect 2594 1266 2597 1333
rect 2610 1273 2613 1336
rect 2618 1323 2621 1343
rect 2626 1323 2629 1346
rect 2594 1263 2605 1266
rect 2538 1213 2541 1236
rect 2538 1093 2541 1206
rect 2554 1176 2557 1243
rect 2546 1173 2557 1176
rect 2538 1003 2541 1016
rect 2538 923 2541 976
rect 2546 853 2549 1173
rect 2586 1163 2589 1206
rect 2554 1133 2557 1156
rect 2570 1123 2589 1126
rect 2562 1113 2581 1116
rect 2578 1096 2581 1113
rect 2574 1093 2581 1096
rect 2574 1036 2577 1093
rect 2574 1033 2581 1036
rect 2538 813 2541 846
rect 2546 806 2549 816
rect 2538 803 2549 806
rect 2554 783 2557 1026
rect 2562 893 2565 1016
rect 2578 1013 2581 1033
rect 2586 966 2589 1123
rect 2594 1103 2597 1116
rect 2594 1013 2597 1026
rect 2594 993 2597 1006
rect 2578 963 2589 966
rect 2578 936 2581 963
rect 2570 933 2581 936
rect 2586 933 2589 946
rect 2594 933 2597 976
rect 2562 756 2565 856
rect 2570 813 2573 826
rect 2578 796 2581 926
rect 2570 793 2581 796
rect 2570 763 2573 793
rect 2586 786 2589 856
rect 2594 813 2597 926
rect 2578 783 2589 786
rect 2578 756 2581 783
rect 2554 753 2565 756
rect 2570 753 2581 756
rect 2554 746 2557 753
rect 2530 743 2557 746
rect 2530 733 2533 743
rect 2546 733 2549 743
rect 2562 726 2565 746
rect 2514 713 2521 716
rect 2518 646 2521 713
rect 2530 703 2533 726
rect 2518 643 2525 646
rect 2490 623 2493 636
rect 2506 633 2517 636
rect 2498 583 2501 616
rect 2482 573 2509 576
rect 2458 333 2477 336
rect 2458 213 2461 326
rect 2482 323 2485 546
rect 2490 503 2493 516
rect 2490 413 2493 486
rect 2506 466 2509 573
rect 2514 483 2517 633
rect 2522 526 2525 643
rect 2530 533 2533 616
rect 2538 613 2541 626
rect 2538 596 2541 606
rect 2546 603 2549 726
rect 2558 723 2565 726
rect 2558 646 2561 723
rect 2570 653 2573 753
rect 2578 693 2581 726
rect 2586 723 2589 776
rect 2594 706 2597 736
rect 2590 703 2597 706
rect 2558 643 2565 646
rect 2562 626 2565 643
rect 2590 636 2593 703
rect 2602 643 2605 1263
rect 2618 1153 2621 1316
rect 2626 1213 2629 1296
rect 2626 1123 2629 1136
rect 2626 1066 2629 1086
rect 2622 1063 2629 1066
rect 2610 923 2613 1016
rect 2622 986 2625 1063
rect 2634 996 2637 1556
rect 2642 1516 2645 1816
rect 2650 1793 2653 1806
rect 2658 1746 2661 1816
rect 2682 1803 2685 1826
rect 2690 1803 2693 1996
rect 2698 1913 2701 1926
rect 2698 1823 2701 1856
rect 2658 1743 2685 1746
rect 2658 1723 2661 1736
rect 2666 1713 2669 1736
rect 2674 1703 2677 1726
rect 2650 1643 2669 1646
rect 2650 1633 2653 1643
rect 2650 1613 2653 1626
rect 2658 1606 2661 1636
rect 2666 1623 2669 1643
rect 2658 1603 2677 1606
rect 2674 1546 2677 1596
rect 2682 1586 2685 1743
rect 2690 1723 2693 1796
rect 2698 1763 2701 1806
rect 2698 1703 2701 1726
rect 2690 1593 2693 1626
rect 2682 1583 2693 1586
rect 2674 1543 2685 1546
rect 2650 1533 2677 1536
rect 2682 1533 2685 1543
rect 2674 1526 2677 1533
rect 2642 1513 2649 1516
rect 2646 1446 2649 1513
rect 2642 1443 2649 1446
rect 2642 1253 2645 1443
rect 2650 1403 2653 1426
rect 2650 1373 2653 1396
rect 2658 1363 2661 1526
rect 2674 1523 2685 1526
rect 2690 1516 2693 1583
rect 2698 1533 2701 1696
rect 2706 1623 2709 1936
rect 2714 1933 2717 2016
rect 2722 2013 2725 2056
rect 2722 1916 2725 1976
rect 2718 1913 2725 1916
rect 2718 1846 2721 1913
rect 2730 1863 2733 2366
rect 2746 2326 2749 2396
rect 2794 2393 2805 2396
rect 2794 2353 2797 2393
rect 2742 2323 2749 2326
rect 2742 2226 2745 2323
rect 2754 2273 2757 2316
rect 2762 2256 2765 2336
rect 2786 2326 2789 2336
rect 2802 2333 2805 2376
rect 2818 2353 2821 2416
rect 2842 2413 2853 2416
rect 2866 2403 2869 2416
rect 2898 2366 2901 2423
rect 2914 2376 2917 2416
rect 2914 2373 2925 2376
rect 2898 2363 2909 2366
rect 2858 2333 2861 2356
rect 2866 2333 2869 2346
rect 2770 2306 2773 2326
rect 2786 2323 2797 2326
rect 2834 2323 2901 2326
rect 2770 2303 2777 2306
rect 2786 2303 2789 2316
rect 2754 2253 2765 2256
rect 2742 2223 2749 2226
rect 2738 2193 2741 2206
rect 2738 2113 2741 2126
rect 2738 2023 2741 2066
rect 2738 2003 2741 2016
rect 2718 1843 2725 1846
rect 2674 1466 2677 1516
rect 2690 1513 2697 1516
rect 2666 1463 2677 1466
rect 2666 1413 2669 1463
rect 2674 1403 2677 1416
rect 2682 1373 2685 1496
rect 2694 1426 2697 1513
rect 2690 1423 2697 1426
rect 2650 1343 2685 1346
rect 2650 1206 2653 1216
rect 2642 1203 2653 1206
rect 2658 1193 2661 1336
rect 2666 1233 2677 1236
rect 2666 1213 2669 1233
rect 2682 1226 2685 1343
rect 2690 1323 2693 1423
rect 2682 1223 2693 1226
rect 2666 1166 2669 1206
rect 2650 1163 2669 1166
rect 2650 1126 2653 1163
rect 2642 1123 2653 1126
rect 2658 1123 2661 1156
rect 2666 1133 2677 1136
rect 2642 1083 2645 1123
rect 2666 1106 2669 1126
rect 2642 1013 2645 1076
rect 2650 1003 2653 1106
rect 2662 1103 2669 1106
rect 2662 1036 2665 1103
rect 2662 1033 2669 1036
rect 2674 1033 2677 1133
rect 2682 1113 2685 1216
rect 2690 1133 2693 1223
rect 2698 1203 2701 1406
rect 2706 1103 2709 1606
rect 2714 1533 2717 1826
rect 2722 1803 2725 1843
rect 2730 1813 2733 1826
rect 2738 1803 2741 1936
rect 2746 1903 2749 2223
rect 2754 2166 2757 2253
rect 2762 2203 2765 2246
rect 2774 2216 2777 2303
rect 2794 2273 2797 2323
rect 2874 2296 2877 2316
rect 2898 2306 2901 2323
rect 2866 2293 2877 2296
rect 2866 2236 2869 2293
rect 2866 2233 2877 2236
rect 2786 2223 2805 2226
rect 2774 2213 2789 2216
rect 2786 2203 2789 2213
rect 2754 2163 2773 2166
rect 2794 2163 2797 2216
rect 2802 2173 2805 2223
rect 2810 2183 2813 2226
rect 2874 2216 2877 2233
rect 2882 2223 2885 2306
rect 2894 2303 2901 2306
rect 2894 2226 2897 2303
rect 2894 2223 2901 2226
rect 2906 2223 2909 2363
rect 2922 2333 2925 2373
rect 2934 2356 2937 2453
rect 2946 2413 2949 2473
rect 2954 2433 2957 2616
rect 2986 2613 2989 2756
rect 3002 2656 3005 2736
rect 3050 2723 3053 2763
rect 3074 2753 3077 2806
rect 3074 2726 3077 2746
rect 3082 2733 3085 2816
rect 3070 2723 3077 2726
rect 2998 2653 3005 2656
rect 2998 2596 3001 2653
rect 3058 2616 3061 2686
rect 3070 2636 3073 2723
rect 3070 2633 3077 2636
rect 3034 2603 3037 2616
rect 3058 2613 3065 2616
rect 2998 2593 3005 2596
rect 3002 2573 3005 2593
rect 3034 2523 3037 2596
rect 3034 2503 3037 2516
rect 3050 2513 3053 2606
rect 3062 2566 3065 2613
rect 3058 2563 3065 2566
rect 3058 2543 3061 2563
rect 3066 2533 3069 2546
rect 3074 2526 3077 2633
rect 3082 2606 3085 2726
rect 3098 2656 3101 2823
rect 3130 2813 3149 2816
rect 3122 2686 3125 2806
rect 3146 2763 3149 2806
rect 3154 2736 3157 2833
rect 3154 2733 3165 2736
rect 3170 2726 3173 2826
rect 3090 2653 3101 2656
rect 3114 2683 3125 2686
rect 3130 2723 3173 2726
rect 3090 2633 3093 2653
rect 3090 2613 3093 2626
rect 3114 2616 3117 2683
rect 3130 2623 3133 2723
rect 3146 2633 3149 2706
rect 3154 2633 3157 2716
rect 3186 2713 3189 2843
rect 3198 2756 3201 2863
rect 3198 2753 3205 2756
rect 3194 2683 3197 2736
rect 3202 2726 3205 2753
rect 3210 2743 3213 3206
rect 3290 3136 3293 3216
rect 3298 3213 3301 3253
rect 3362 3223 3397 3226
rect 3306 3193 3309 3206
rect 3322 3146 3325 3206
rect 3330 3163 3333 3216
rect 3354 3193 3357 3206
rect 3362 3183 3365 3216
rect 3370 3173 3373 3206
rect 3394 3203 3397 3223
rect 3402 3166 3405 3206
rect 3354 3163 3405 3166
rect 3322 3143 3333 3146
rect 3226 3096 3229 3136
rect 3274 3133 3293 3136
rect 3234 3113 3237 3126
rect 3226 3093 3237 3096
rect 3234 3026 3237 3093
rect 3274 3033 3277 3133
rect 3282 3106 3285 3126
rect 3306 3106 3309 3136
rect 3282 3103 3309 3106
rect 3306 3026 3309 3103
rect 3226 3023 3237 3026
rect 3218 2973 3221 3016
rect 3226 3003 3229 3023
rect 3266 3016 3269 3026
rect 3306 3023 3313 3026
rect 3266 3013 3285 3016
rect 3290 3013 3301 3016
rect 3242 2933 3245 2956
rect 3258 2943 3261 3006
rect 3266 2986 3269 3013
rect 3274 3003 3285 3006
rect 3266 2983 3277 2986
rect 3226 2783 3229 2816
rect 3202 2723 3209 2726
rect 3206 2676 3209 2723
rect 3202 2673 3209 2676
rect 3082 2603 3093 2606
rect 3066 2523 3077 2526
rect 2970 2403 2973 2416
rect 2930 2353 2937 2356
rect 2930 2323 2933 2353
rect 2938 2323 2941 2336
rect 2954 2333 2957 2376
rect 2770 2156 2773 2163
rect 2754 2043 2757 2136
rect 2762 2026 2765 2156
rect 2770 2153 2797 2156
rect 2770 2133 2773 2146
rect 2794 2133 2797 2153
rect 2810 2126 2813 2146
rect 2826 2133 2845 2136
rect 2770 2053 2773 2126
rect 2810 2123 2821 2126
rect 2778 2046 2781 2116
rect 2758 2023 2765 2026
rect 2770 2043 2781 2046
rect 2786 2113 2797 2116
rect 2758 1896 2761 2023
rect 2770 1906 2773 2043
rect 2786 2013 2789 2113
rect 2802 2013 2805 2046
rect 2810 2006 2813 2056
rect 2778 2003 2797 2006
rect 2802 2003 2813 2006
rect 2778 1923 2781 2003
rect 2802 1933 2805 2003
rect 2794 1906 2797 1926
rect 2770 1903 2781 1906
rect 2746 1893 2761 1896
rect 2746 1796 2749 1893
rect 2722 1603 2725 1756
rect 2722 1543 2725 1596
rect 2730 1526 2733 1796
rect 2738 1793 2749 1796
rect 2738 1733 2741 1793
rect 2754 1786 2757 1826
rect 2762 1793 2765 1866
rect 2778 1846 2781 1903
rect 2770 1843 2781 1846
rect 2790 1903 2797 1906
rect 2746 1783 2757 1786
rect 2738 1533 2741 1716
rect 2746 1666 2749 1783
rect 2754 1683 2757 1766
rect 2770 1746 2773 1843
rect 2790 1826 2793 1903
rect 2778 1823 2793 1826
rect 2778 1813 2781 1823
rect 2802 1816 2805 1926
rect 2794 1813 2805 1816
rect 2810 1813 2813 1926
rect 2762 1743 2773 1746
rect 2762 1673 2765 1743
rect 2746 1663 2765 1666
rect 2762 1623 2765 1663
rect 2746 1613 2757 1616
rect 2714 1473 2717 1526
rect 2730 1523 2741 1526
rect 2722 1513 2733 1516
rect 2722 1416 2725 1513
rect 2738 1506 2741 1523
rect 2714 1413 2725 1416
rect 2730 1503 2741 1506
rect 2722 1393 2725 1406
rect 2714 1203 2717 1376
rect 2722 1196 2725 1366
rect 2718 1193 2725 1196
rect 2718 1096 2721 1193
rect 2714 1093 2721 1096
rect 2690 1056 2693 1076
rect 2690 1053 2697 1056
rect 2634 993 2641 996
rect 2622 983 2629 986
rect 2610 736 2613 916
rect 2618 913 2621 966
rect 2626 923 2629 983
rect 2638 916 2641 993
rect 2658 973 2661 1016
rect 2666 993 2669 1033
rect 2658 933 2661 966
rect 2634 913 2641 916
rect 2650 913 2653 926
rect 2618 813 2621 896
rect 2626 823 2629 836
rect 2610 733 2621 736
rect 2626 726 2629 816
rect 2618 723 2629 726
rect 2562 623 2573 626
rect 2554 596 2557 616
rect 2538 593 2557 596
rect 2562 566 2565 606
rect 2522 523 2533 526
rect 2530 503 2533 523
rect 2546 506 2549 566
rect 2554 563 2565 566
rect 2554 523 2557 563
rect 2570 523 2573 623
rect 2578 596 2581 636
rect 2590 633 2597 636
rect 2594 613 2597 633
rect 2618 613 2621 723
rect 2634 706 2637 913
rect 2666 863 2669 926
rect 2642 813 2645 826
rect 2674 816 2677 1026
rect 2682 1023 2685 1036
rect 2682 853 2685 1016
rect 2694 956 2697 1053
rect 2690 953 2697 956
rect 2706 953 2709 1016
rect 2714 996 2717 1093
rect 2722 1006 2725 1026
rect 2730 1013 2733 1503
rect 2746 1466 2749 1556
rect 2754 1526 2757 1536
rect 2762 1533 2765 1606
rect 2770 1603 2773 1736
rect 2770 1533 2773 1556
rect 2754 1523 2765 1526
rect 2738 1463 2749 1466
rect 2738 1353 2741 1463
rect 2738 1323 2741 1346
rect 2746 1333 2749 1426
rect 2738 1196 2741 1256
rect 2746 1203 2749 1306
rect 2738 1193 2749 1196
rect 2738 1123 2741 1146
rect 2738 1013 2741 1116
rect 2722 1003 2733 1006
rect 2714 993 2741 996
rect 2666 813 2677 816
rect 2666 793 2669 813
rect 2690 806 2693 953
rect 2698 933 2717 936
rect 2722 933 2725 986
rect 2698 876 2701 933
rect 2714 926 2717 933
rect 2706 896 2709 926
rect 2714 923 2725 926
rect 2714 913 2725 916
rect 2730 896 2733 976
rect 2738 923 2741 993
rect 2746 966 2749 1193
rect 2754 1136 2757 1516
rect 2762 1493 2765 1523
rect 2770 1506 2773 1526
rect 2778 1523 2781 1806
rect 2786 1763 2789 1806
rect 2770 1503 2777 1506
rect 2762 1403 2765 1466
rect 2774 1416 2777 1503
rect 2774 1413 2781 1416
rect 2778 1396 2781 1413
rect 2762 1343 2765 1396
rect 2774 1393 2781 1396
rect 2762 1313 2765 1336
rect 2774 1306 2777 1393
rect 2786 1376 2789 1756
rect 2794 1686 2797 1806
rect 2802 1703 2805 1726
rect 2810 1693 2813 1806
rect 2818 1733 2821 2123
rect 2826 2106 2829 2126
rect 2842 2123 2845 2133
rect 2850 2106 2853 2216
rect 2826 2103 2837 2106
rect 2834 2026 2837 2103
rect 2846 2103 2853 2106
rect 2846 2036 2849 2103
rect 2846 2033 2853 2036
rect 2826 2023 2837 2026
rect 2826 2003 2829 2023
rect 2850 2013 2853 2033
rect 2826 1923 2829 1956
rect 2834 1933 2837 2006
rect 2842 1916 2845 2006
rect 2858 1966 2861 2206
rect 2866 2193 2869 2216
rect 2874 2213 2885 2216
rect 2882 2203 2885 2213
rect 2866 2113 2869 2186
rect 2890 2156 2893 2206
rect 2874 2153 2893 2156
rect 2874 2143 2877 2153
rect 2866 2023 2869 2076
rect 2866 1983 2869 2006
rect 2850 1923 2853 1966
rect 2858 1963 2865 1966
rect 2838 1913 2845 1916
rect 2826 1763 2829 1906
rect 2838 1826 2841 1913
rect 2838 1823 2845 1826
rect 2850 1823 2853 1916
rect 2862 1836 2865 1963
rect 2858 1833 2865 1836
rect 2834 1793 2837 1806
rect 2826 1733 2829 1756
rect 2826 1713 2829 1726
rect 2834 1703 2837 1726
rect 2794 1683 2829 1686
rect 2818 1656 2821 1676
rect 2814 1653 2821 1656
rect 2802 1623 2805 1636
rect 2794 1453 2797 1616
rect 2814 1546 2817 1653
rect 2814 1543 2821 1546
rect 2794 1383 2797 1406
rect 2786 1373 2797 1376
rect 2770 1303 2777 1306
rect 2762 1213 2765 1236
rect 2762 1153 2765 1196
rect 2770 1173 2773 1303
rect 2754 1133 2761 1136
rect 2758 1006 2761 1133
rect 2754 1003 2761 1006
rect 2754 983 2757 1003
rect 2746 963 2757 966
rect 2754 916 2757 963
rect 2706 893 2717 896
rect 2698 873 2705 876
rect 2702 816 2705 873
rect 2674 803 2693 806
rect 2698 813 2705 816
rect 2698 796 2701 813
rect 2690 793 2701 796
rect 2630 703 2637 706
rect 2630 646 2633 703
rect 2630 643 2637 646
rect 2634 626 2637 643
rect 2642 633 2645 786
rect 2634 623 2645 626
rect 2626 613 2637 616
rect 2642 596 2645 623
rect 2650 613 2653 756
rect 2690 746 2693 793
rect 2674 743 2693 746
rect 2658 723 2661 736
rect 2658 683 2661 716
rect 2666 666 2669 726
rect 2674 693 2677 743
rect 2714 736 2717 893
rect 2726 893 2733 896
rect 2726 766 2729 893
rect 2726 763 2733 766
rect 2682 703 2685 726
rect 2662 663 2669 666
rect 2662 606 2665 663
rect 2578 593 2585 596
rect 2582 516 2585 593
rect 2634 593 2645 596
rect 2578 513 2585 516
rect 2546 503 2557 506
rect 2506 463 2525 466
rect 2498 383 2501 406
rect 2474 193 2477 226
rect 2482 186 2485 316
rect 2498 293 2501 316
rect 2506 233 2509 456
rect 2522 446 2525 463
rect 2514 413 2517 446
rect 2522 443 2529 446
rect 2514 323 2517 406
rect 2526 316 2529 443
rect 2538 413 2541 496
rect 2554 436 2557 503
rect 2546 433 2557 436
rect 2546 406 2549 433
rect 2578 416 2581 513
rect 2522 313 2529 316
rect 2538 403 2549 406
rect 2554 413 2581 416
rect 2594 413 2597 536
rect 2602 523 2605 546
rect 2634 536 2637 593
rect 2602 513 2613 516
rect 2602 493 2605 513
rect 2618 506 2621 536
rect 2634 533 2645 536
rect 2642 513 2645 533
rect 2650 523 2653 606
rect 2658 603 2665 606
rect 2658 563 2661 603
rect 2658 523 2661 536
rect 2666 516 2669 596
rect 2658 513 2669 516
rect 2674 513 2677 646
rect 2690 603 2693 736
rect 2706 733 2717 736
rect 2722 733 2725 746
rect 2682 533 2685 556
rect 2610 503 2621 506
rect 2610 426 2613 503
rect 2666 486 2669 506
rect 2690 486 2693 586
rect 2698 526 2701 726
rect 2706 686 2709 733
rect 2714 693 2717 726
rect 2722 686 2725 726
rect 2706 683 2725 686
rect 2706 543 2709 596
rect 2714 583 2717 616
rect 2730 606 2733 763
rect 2738 703 2741 916
rect 2746 913 2757 916
rect 2746 893 2749 913
rect 2770 883 2773 1146
rect 2778 1113 2781 1216
rect 2786 1096 2789 1326
rect 2794 1306 2797 1373
rect 2802 1326 2805 1536
rect 2810 1353 2813 1526
rect 2818 1363 2821 1543
rect 2826 1343 2829 1683
rect 2834 1533 2837 1636
rect 2842 1596 2845 1823
rect 2850 1773 2853 1816
rect 2850 1633 2853 1766
rect 2858 1733 2861 1833
rect 2866 1713 2869 1816
rect 2874 1786 2877 2126
rect 2882 2106 2885 2136
rect 2890 2123 2893 2146
rect 2882 2103 2889 2106
rect 2886 2036 2889 2103
rect 2882 2033 2889 2036
rect 2882 1946 2885 2033
rect 2890 2003 2893 2016
rect 2898 2013 2901 2223
rect 2914 2183 2917 2216
rect 2922 2206 2925 2316
rect 2930 2223 2933 2306
rect 2922 2203 2933 2206
rect 2938 2196 2941 2246
rect 2978 2206 2981 2246
rect 2994 2226 2997 2446
rect 3042 2416 3045 2476
rect 3010 2333 3013 2416
rect 3042 2413 3053 2416
rect 3066 2336 3069 2523
rect 3090 2413 3093 2526
rect 3098 2503 3101 2616
rect 3114 2613 3141 2616
rect 3130 2593 3133 2613
rect 3170 2606 3173 2646
rect 3138 2603 3165 2606
rect 3170 2603 3181 2606
rect 3138 2516 3141 2603
rect 3178 2546 3181 2603
rect 3186 2583 3189 2626
rect 3202 2603 3205 2673
rect 3218 2613 3221 2736
rect 3234 2706 3237 2836
rect 3242 2823 3245 2926
rect 3274 2886 3277 2983
rect 3290 2923 3293 3013
rect 3310 2966 3313 3023
rect 3310 2963 3317 2966
rect 3250 2883 3277 2886
rect 3250 2803 3253 2883
rect 3290 2766 3293 2826
rect 3290 2763 3301 2766
rect 3266 2716 3269 2736
rect 3282 2726 3285 2736
rect 3258 2713 3269 2716
rect 3274 2723 3285 2726
rect 3234 2703 3245 2706
rect 3242 2646 3245 2703
rect 3234 2643 3245 2646
rect 3258 2646 3261 2713
rect 3258 2643 3269 2646
rect 3234 2613 3237 2643
rect 3266 2626 3269 2643
rect 3242 2623 3269 2626
rect 3210 2586 3213 2606
rect 3226 2593 3229 2606
rect 3242 2603 3245 2623
rect 3250 2586 3253 2596
rect 3210 2583 3253 2586
rect 3162 2533 3165 2546
rect 3178 2543 3205 2546
rect 3130 2513 3141 2516
rect 3146 2523 3165 2526
rect 3178 2523 3181 2543
rect 3186 2533 3197 2536
rect 3130 2466 3133 2513
rect 3130 2463 3137 2466
rect 3090 2336 3093 2406
rect 3034 2316 3037 2336
rect 3050 2333 3069 2336
rect 3026 2313 3037 2316
rect 3042 2313 3045 2326
rect 3026 2246 3029 2313
rect 3026 2243 3037 2246
rect 2994 2223 3013 2226
rect 2986 2213 3005 2216
rect 2930 2193 2941 2196
rect 2906 2133 2909 2176
rect 2906 2033 2909 2116
rect 2914 2083 2917 2126
rect 2930 2086 2933 2193
rect 2946 2113 2949 2206
rect 2978 2203 2989 2206
rect 2994 2203 2997 2213
rect 2926 2083 2933 2086
rect 2926 2026 2929 2083
rect 2914 1966 2917 2026
rect 2926 2023 2933 2026
rect 2906 1963 2917 1966
rect 2882 1943 2917 1946
rect 2882 1813 2885 1846
rect 2890 1813 2893 1936
rect 2914 1933 2917 1943
rect 2914 1913 2917 1926
rect 2874 1783 2885 1786
rect 2874 1706 2877 1776
rect 2882 1763 2885 1783
rect 2890 1743 2893 1806
rect 2898 1803 2901 1856
rect 2906 1733 2909 1756
rect 2922 1753 2925 2006
rect 2930 1933 2933 2023
rect 2938 1923 2941 2076
rect 2954 2036 2957 2136
rect 2946 2033 2957 2036
rect 2946 1986 2949 2033
rect 2962 2026 2965 2136
rect 2978 2133 2981 2146
rect 2970 2093 2973 2126
rect 2986 2123 2989 2203
rect 3002 2193 3005 2206
rect 3010 2153 3013 2223
rect 2954 2023 2965 2026
rect 2954 2003 2957 2023
rect 2946 1983 2953 1986
rect 2950 1916 2953 1983
rect 2962 1943 2965 2016
rect 2978 2003 2981 2056
rect 2986 2003 2989 2116
rect 2994 1993 2997 2136
rect 3002 1983 3005 2076
rect 3002 1936 3005 1956
rect 2970 1933 3005 1936
rect 3010 1933 3013 2136
rect 3018 2063 3021 2226
rect 3026 2173 3029 2206
rect 3018 2013 3021 2056
rect 3018 1963 3021 2006
rect 2946 1913 2953 1916
rect 2930 1793 2933 1806
rect 2922 1726 2925 1746
rect 2930 1733 2933 1766
rect 2866 1703 2877 1706
rect 2866 1623 2869 1703
rect 2850 1603 2853 1616
rect 2874 1603 2877 1626
rect 2842 1593 2877 1596
rect 2850 1546 2853 1566
rect 2850 1543 2861 1546
rect 2850 1523 2853 1536
rect 2834 1503 2837 1516
rect 2834 1403 2837 1416
rect 2842 1383 2845 1456
rect 2850 1376 2853 1476
rect 2842 1373 2853 1376
rect 2834 1336 2837 1366
rect 2826 1333 2837 1336
rect 2842 1326 2845 1373
rect 2802 1323 2813 1326
rect 2794 1303 2801 1306
rect 2798 1146 2801 1303
rect 2782 1093 2789 1096
rect 2794 1143 2801 1146
rect 2782 1006 2785 1093
rect 2794 1073 2797 1143
rect 2794 1033 2797 1066
rect 2802 1033 2805 1126
rect 2810 1123 2813 1323
rect 2818 1293 2821 1326
rect 2834 1323 2845 1326
rect 2834 1216 2837 1323
rect 2850 1306 2853 1336
rect 2846 1303 2853 1306
rect 2846 1236 2849 1303
rect 2846 1233 2853 1236
rect 2818 1203 2821 1216
rect 2826 1213 2837 1216
rect 2826 1183 2829 1213
rect 2842 1206 2845 1216
rect 2834 1203 2845 1206
rect 2850 1203 2853 1233
rect 2794 1016 2797 1026
rect 2794 1013 2805 1016
rect 2782 1003 2789 1006
rect 2786 953 2789 1003
rect 2802 923 2805 1013
rect 2810 916 2813 1106
rect 2818 1023 2821 1176
rect 2834 1153 2837 1203
rect 2842 1123 2845 1196
rect 2802 913 2813 916
rect 2818 913 2821 956
rect 2826 943 2829 1116
rect 2834 1103 2845 1106
rect 2850 1103 2853 1116
rect 2834 1023 2837 1103
rect 2842 1013 2845 1036
rect 2858 1016 2861 1543
rect 2866 1523 2869 1556
rect 2866 1403 2869 1446
rect 2866 1336 2869 1346
rect 2874 1343 2877 1593
rect 2882 1523 2885 1726
rect 2906 1723 2917 1726
rect 2922 1723 2933 1726
rect 2906 1716 2909 1723
rect 2890 1713 2909 1716
rect 2890 1593 2893 1616
rect 2898 1543 2901 1616
rect 2906 1583 2909 1606
rect 2922 1533 2925 1626
rect 2930 1533 2933 1556
rect 2938 1533 2941 1816
rect 2946 1796 2949 1913
rect 2962 1806 2965 1926
rect 2978 1923 2989 1926
rect 3026 1916 3029 2156
rect 3034 2046 3037 2243
rect 3042 2193 3045 2226
rect 3042 2113 3045 2126
rect 3042 2066 3045 2106
rect 3050 2073 3053 2333
rect 3058 2233 3061 2326
rect 3074 2323 3077 2336
rect 3090 2333 3097 2336
rect 3074 2303 3077 2316
rect 3082 2313 3085 2326
rect 3058 2133 3061 2226
rect 3066 2183 3069 2206
rect 3074 2203 3077 2216
rect 3058 2103 3061 2116
rect 3042 2063 3053 2066
rect 3034 2043 3041 2046
rect 3038 1966 3041 2043
rect 3050 2023 3053 2063
rect 3050 2003 3053 2016
rect 3058 2003 3061 2066
rect 3066 2003 3069 2146
rect 3074 2086 3077 2196
rect 3082 2103 3085 2286
rect 3094 2156 3097 2333
rect 3106 2316 3109 2376
rect 3134 2366 3137 2463
rect 3146 2386 3149 2523
rect 3186 2516 3189 2533
rect 3162 2513 3189 2516
rect 3202 2456 3205 2543
rect 3210 2476 3213 2583
rect 3250 2566 3253 2583
rect 3226 2563 3245 2566
rect 3250 2563 3269 2566
rect 3226 2506 3229 2563
rect 3242 2533 3245 2563
rect 3226 2503 3237 2506
rect 3210 2473 3221 2476
rect 3154 2453 3197 2456
rect 3202 2453 3209 2456
rect 3154 2413 3157 2453
rect 3170 2403 3173 2436
rect 3194 2413 3197 2453
rect 3206 2406 3209 2453
rect 3202 2403 3209 2406
rect 3146 2383 3165 2386
rect 3134 2363 3141 2366
rect 3138 2343 3141 2363
rect 3162 2323 3165 2383
rect 3106 2313 3117 2316
rect 3114 2256 3117 2313
rect 3170 2296 3173 2316
rect 3106 2253 3117 2256
rect 3162 2293 3173 2296
rect 3106 2186 3109 2253
rect 3162 2236 3165 2293
rect 3114 2216 3117 2236
rect 3162 2233 3173 2236
rect 3122 2223 3133 2226
rect 3114 2213 3125 2216
rect 3130 2213 3141 2216
rect 3122 2203 3125 2213
rect 3138 2203 3149 2206
rect 3106 2183 3125 2186
rect 3090 2153 3097 2156
rect 3074 2083 3081 2086
rect 3034 1963 3041 1966
rect 3034 1943 3037 1963
rect 3034 1923 3045 1926
rect 2970 1913 2997 1916
rect 3018 1913 3029 1916
rect 2970 1896 2973 1913
rect 2970 1893 2981 1896
rect 2978 1836 2981 1893
rect 2970 1833 2981 1836
rect 3018 1836 3021 1913
rect 3018 1833 3029 1836
rect 2970 1813 2973 1833
rect 2962 1803 2973 1806
rect 2946 1793 2965 1796
rect 2946 1693 2949 1726
rect 2954 1636 2957 1786
rect 2962 1716 2965 1793
rect 2970 1783 2973 1803
rect 3002 1783 3005 1816
rect 3026 1813 3029 1833
rect 3034 1806 3037 1916
rect 3042 1823 3045 1923
rect 3010 1793 3013 1806
rect 2970 1733 2973 1746
rect 2986 1733 2989 1766
rect 2994 1733 2997 1756
rect 2978 1723 2989 1726
rect 3002 1723 3005 1736
rect 2962 1713 2973 1716
rect 2970 1656 2973 1713
rect 2986 1703 2989 1723
rect 3010 1706 3013 1726
rect 3002 1703 3013 1706
rect 2970 1653 2981 1656
rect 2950 1633 2957 1636
rect 2950 1576 2953 1633
rect 2962 1583 2965 1626
rect 2970 1623 2973 1636
rect 2978 1616 2981 1653
rect 2986 1623 2989 1696
rect 3002 1646 3005 1703
rect 3002 1643 3013 1646
rect 3010 1623 3013 1643
rect 2970 1613 2997 1616
rect 2970 1603 2973 1613
rect 2950 1573 2957 1576
rect 2898 1496 2901 1516
rect 2894 1493 2901 1496
rect 2882 1413 2885 1466
rect 2894 1426 2897 1493
rect 2894 1423 2901 1426
rect 2890 1386 2893 1406
rect 2886 1383 2893 1386
rect 2866 1333 2877 1336
rect 2866 1293 2869 1326
rect 2874 1276 2877 1333
rect 2886 1296 2889 1383
rect 2898 1306 2901 1423
rect 2906 1403 2909 1526
rect 2954 1516 2957 1573
rect 2986 1546 2989 1606
rect 2994 1596 2997 1613
rect 2994 1593 3013 1596
rect 2986 1543 2997 1546
rect 2922 1503 2925 1516
rect 2946 1513 2957 1516
rect 2946 1426 2949 1513
rect 2962 1433 2965 1526
rect 2978 1503 2981 1516
rect 2946 1423 2957 1426
rect 2962 1423 2973 1426
rect 2906 1363 2909 1396
rect 2922 1373 2925 1406
rect 2938 1386 2941 1406
rect 2906 1333 2909 1356
rect 2914 1323 2917 1336
rect 2922 1306 2925 1366
rect 2930 1333 2933 1386
rect 2938 1383 2945 1386
rect 2898 1303 2909 1306
rect 2886 1293 2893 1296
rect 2866 1273 2877 1276
rect 2866 1193 2869 1273
rect 2874 1193 2877 1266
rect 2890 1236 2893 1293
rect 2886 1233 2893 1236
rect 2886 1156 2889 1233
rect 2866 1023 2869 1156
rect 2886 1153 2893 1156
rect 2898 1153 2901 1216
rect 2906 1176 2909 1303
rect 2918 1303 2925 1306
rect 2918 1226 2921 1303
rect 2930 1243 2933 1326
rect 2942 1236 2945 1383
rect 2938 1233 2945 1236
rect 2918 1223 2925 1226
rect 2922 1203 2925 1223
rect 2930 1203 2933 1226
rect 2914 1193 2933 1196
rect 2930 1176 2933 1193
rect 2906 1173 2917 1176
rect 2890 1113 2893 1153
rect 2898 1113 2901 1146
rect 2914 1106 2917 1173
rect 2874 1023 2877 1106
rect 2882 1073 2885 1106
rect 2906 1103 2917 1106
rect 2926 1173 2933 1176
rect 2850 936 2853 1016
rect 2858 1013 2869 1016
rect 2866 956 2869 1013
rect 2866 953 2877 956
rect 2850 933 2861 936
rect 2850 913 2853 926
rect 2858 906 2861 933
rect 2874 913 2877 953
rect 2882 906 2885 1036
rect 2810 903 2829 906
rect 2858 903 2885 906
rect 2826 893 2829 903
rect 2890 896 2893 1036
rect 2898 913 2901 1016
rect 2906 913 2909 1103
rect 2926 1096 2929 1173
rect 2926 1093 2933 1096
rect 2914 1073 2925 1076
rect 2922 1033 2925 1073
rect 2930 1016 2933 1093
rect 2938 1053 2941 1233
rect 2946 1123 2949 1216
rect 2954 1076 2957 1423
rect 2978 1393 2981 1436
rect 2986 1403 2989 1536
rect 2994 1463 2997 1543
rect 2994 1423 2997 1446
rect 3002 1413 3005 1576
rect 3010 1523 3013 1593
rect 3010 1453 3013 1516
rect 2986 1343 2989 1356
rect 2978 1316 2981 1336
rect 2986 1323 2989 1336
rect 2974 1313 2981 1316
rect 2962 1213 2965 1296
rect 2974 1236 2977 1313
rect 2974 1233 2981 1236
rect 2970 1173 2973 1206
rect 2978 1183 2981 1233
rect 2986 1166 2989 1316
rect 2962 1163 2989 1166
rect 2962 1123 2965 1163
rect 2994 1156 2997 1256
rect 3010 1216 3013 1436
rect 3018 1373 3021 1806
rect 3026 1803 3037 1806
rect 3026 1613 3029 1803
rect 3034 1613 3037 1786
rect 3042 1743 3045 1806
rect 3042 1723 3045 1736
rect 3050 1716 3053 1986
rect 3058 1933 3061 1966
rect 3066 1933 3069 1956
rect 3078 1946 3081 2083
rect 3074 1943 3081 1946
rect 3058 1896 3061 1916
rect 3058 1893 3065 1896
rect 3062 1816 3065 1893
rect 3058 1813 3065 1816
rect 3074 1813 3077 1943
rect 3090 1936 3093 2153
rect 3098 2113 3101 2136
rect 3098 1986 3101 2106
rect 3106 2093 3109 2176
rect 3122 2063 3125 2183
rect 3170 2156 3173 2233
rect 3154 2153 3173 2156
rect 3138 2116 3141 2136
rect 3134 2113 3141 2116
rect 3134 2046 3137 2113
rect 3146 2076 3149 2126
rect 3154 2096 3157 2153
rect 3162 2143 3173 2146
rect 3162 2113 3165 2136
rect 3178 2133 3181 2146
rect 3154 2093 3165 2096
rect 3146 2073 3153 2076
rect 3134 2043 3141 2046
rect 3106 2023 3133 2026
rect 3106 2003 3109 2023
rect 3114 1986 3117 2016
rect 3130 2013 3133 2023
rect 3122 1993 3125 2006
rect 3098 1983 3117 1986
rect 3090 1933 3097 1936
rect 3082 1823 3085 1926
rect 3094 1846 3097 1933
rect 3106 1913 3109 1983
rect 3114 1943 3117 1976
rect 3130 1933 3133 2006
rect 3138 1993 3141 2043
rect 3150 2006 3153 2073
rect 3146 2003 3153 2006
rect 3138 1933 3141 1956
rect 3146 1916 3149 2003
rect 3162 1986 3165 2093
rect 3162 1983 3173 1986
rect 3154 1926 3157 1966
rect 3162 1933 3165 1976
rect 3170 1956 3173 1983
rect 3178 1963 3181 2126
rect 3186 2113 3189 2326
rect 3202 2313 3205 2403
rect 3218 2333 3221 2473
rect 3234 2433 3237 2503
rect 3266 2413 3269 2563
rect 3274 2466 3277 2723
rect 3290 2716 3293 2726
rect 3298 2723 3301 2763
rect 3306 2723 3309 2956
rect 3314 2903 3317 2963
rect 3330 2816 3333 3143
rect 3354 3123 3357 3163
rect 3394 3133 3397 3163
rect 3402 3146 3405 3156
rect 3402 3143 3429 3146
rect 3386 3086 3389 3126
rect 3418 3106 3421 3126
rect 3346 3083 3389 3086
rect 3410 3103 3421 3106
rect 3346 3003 3349 3083
rect 3354 3013 3357 3026
rect 3346 2933 3349 2956
rect 3370 2923 3373 3016
rect 3410 2976 3413 3103
rect 3410 2973 3421 2976
rect 3314 2716 3317 2816
rect 3282 2646 3285 2716
rect 3290 2713 3317 2716
rect 3322 2813 3333 2816
rect 3322 2656 3325 2813
rect 3330 2776 3333 2806
rect 3346 2793 3349 2906
rect 3378 2826 3381 2946
rect 3418 2943 3421 2973
rect 3426 2826 3429 3143
rect 3434 3123 3437 3176
rect 3378 2823 3389 2826
rect 3370 2776 3373 2816
rect 3386 2776 3389 2823
rect 3330 2773 3373 2776
rect 3378 2773 3389 2776
rect 3418 2823 3429 2826
rect 3338 2723 3341 2736
rect 3314 2653 3325 2656
rect 3282 2643 3301 2646
rect 3298 2613 3301 2643
rect 3282 2486 3285 2586
rect 3314 2546 3317 2653
rect 3314 2543 3325 2546
rect 3290 2493 3293 2526
rect 3322 2523 3325 2543
rect 3282 2483 3293 2486
rect 3274 2463 3281 2466
rect 3278 2406 3281 2463
rect 3290 2436 3293 2483
rect 3290 2433 3325 2436
rect 3290 2413 3293 2433
rect 3330 2426 3333 2646
rect 3338 2603 3341 2616
rect 3346 2613 3349 2656
rect 3362 2636 3365 2736
rect 3354 2633 3365 2636
rect 3346 2533 3349 2606
rect 3354 2603 3357 2633
rect 3362 2593 3365 2616
rect 3346 2433 3349 2526
rect 3370 2523 3373 2596
rect 3378 2563 3381 2773
rect 3418 2746 3421 2823
rect 3418 2743 3429 2746
rect 3386 2723 3389 2736
rect 3418 2713 3421 2726
rect 3426 2696 3429 2743
rect 3434 2733 3437 2816
rect 3418 2693 3429 2696
rect 3418 2616 3421 2693
rect 3434 2653 3437 2666
rect 3394 2613 3421 2616
rect 3394 2566 3397 2613
rect 3390 2563 3397 2566
rect 3410 2566 3413 2606
rect 3410 2563 3421 2566
rect 3390 2506 3393 2563
rect 3386 2503 3393 2506
rect 3386 2456 3389 2503
rect 3418 2496 3421 2563
rect 3410 2493 3421 2496
rect 3386 2453 3397 2456
rect 3394 2433 3397 2453
rect 3314 2423 3333 2426
rect 3314 2413 3317 2423
rect 3354 2406 3357 2426
rect 3274 2403 3281 2406
rect 3274 2383 3277 2403
rect 3298 2383 3301 2396
rect 3322 2346 3325 2406
rect 3266 2343 3325 2346
rect 3346 2403 3357 2406
rect 3362 2406 3365 2426
rect 3402 2413 3405 2436
rect 3362 2403 3373 2406
rect 3266 2333 3269 2343
rect 3346 2336 3349 2403
rect 3370 2356 3373 2403
rect 3322 2333 3349 2336
rect 3362 2353 3373 2356
rect 3362 2333 3365 2353
rect 3194 2123 3197 2136
rect 3194 1966 3197 2036
rect 3202 2003 3205 2226
rect 3250 2216 3253 2326
rect 3282 2323 3301 2326
rect 3322 2316 3325 2333
rect 3298 2313 3325 2316
rect 3234 2213 3245 2216
rect 3250 2213 3269 2216
rect 3210 2153 3213 2196
rect 3226 2156 3229 2206
rect 3234 2163 3237 2213
rect 3250 2156 3253 2196
rect 3226 2153 3237 2156
rect 3210 2123 3213 2136
rect 3210 2003 3213 2026
rect 3194 1963 3205 1966
rect 3170 1953 3197 1956
rect 3154 1923 3161 1926
rect 3090 1843 3097 1846
rect 3058 1733 3061 1813
rect 3066 1733 3069 1796
rect 3050 1713 3057 1716
rect 3042 1606 3045 1686
rect 3054 1646 3057 1713
rect 3074 1693 3077 1806
rect 3082 1733 3085 1746
rect 3026 1596 3029 1606
rect 3034 1603 3045 1606
rect 3050 1643 3057 1646
rect 3026 1593 3045 1596
rect 3026 1513 3029 1526
rect 3010 1213 3017 1216
rect 3002 1193 3005 1206
rect 2970 1153 2997 1156
rect 2970 1133 2973 1153
rect 3002 1146 3005 1186
rect 3014 1146 3017 1213
rect 2978 1093 2981 1146
rect 2994 1143 3005 1146
rect 3010 1143 3017 1146
rect 2994 1123 2997 1143
rect 2954 1073 2961 1076
rect 2914 1013 2933 1016
rect 2946 1013 2949 1066
rect 2958 1026 2961 1073
rect 2978 1026 2981 1036
rect 2954 1023 2961 1026
rect 2970 1023 2981 1026
rect 2986 1023 2989 1076
rect 2914 903 2917 1013
rect 2922 1003 2941 1006
rect 2866 893 2893 896
rect 2922 893 2925 1003
rect 2954 996 2957 1023
rect 2970 1006 2973 1023
rect 2994 1016 2997 1106
rect 3002 1023 3005 1136
rect 2962 1003 2973 1006
rect 2950 993 2957 996
rect 2930 913 2933 946
rect 2938 923 2941 936
rect 2754 776 2757 806
rect 2786 776 2789 786
rect 2754 773 2789 776
rect 2802 776 2805 816
rect 2834 813 2837 886
rect 2866 846 2869 893
rect 2950 876 2953 993
rect 2962 913 2965 956
rect 2978 923 2981 1016
rect 2986 1013 2997 1016
rect 2986 953 2989 1013
rect 3010 976 3013 1143
rect 3026 1133 3029 1466
rect 3034 1383 3037 1516
rect 3042 1513 3045 1593
rect 3042 1423 3045 1436
rect 3042 1333 3045 1416
rect 3034 1323 3045 1326
rect 3042 1303 3045 1316
rect 3042 1213 3045 1226
rect 3050 1196 3053 1643
rect 3058 1546 3061 1626
rect 3066 1553 3069 1676
rect 3074 1613 3077 1656
rect 3058 1543 3065 1546
rect 3062 1476 3065 1543
rect 3062 1473 3069 1476
rect 3058 1433 3061 1456
rect 3058 1403 3061 1426
rect 3058 1253 3061 1396
rect 3058 1213 3061 1226
rect 3066 1203 3069 1473
rect 3074 1426 3077 1526
rect 3082 1513 3085 1726
rect 3090 1613 3093 1843
rect 3098 1823 3109 1826
rect 3098 1803 3109 1806
rect 3090 1593 3093 1606
rect 3090 1513 3093 1586
rect 3098 1573 3101 1726
rect 3114 1723 3117 1916
rect 3138 1913 3149 1916
rect 3138 1836 3141 1913
rect 3138 1833 3149 1836
rect 3122 1733 3125 1816
rect 3130 1803 3133 1816
rect 3106 1546 3109 1696
rect 3130 1673 3133 1726
rect 3138 1713 3141 1726
rect 3146 1676 3149 1833
rect 3158 1786 3161 1923
rect 3170 1796 3173 1946
rect 3178 1933 3181 1946
rect 3178 1803 3181 1926
rect 3186 1913 3189 1926
rect 3186 1803 3189 1846
rect 3170 1793 3189 1796
rect 3158 1783 3165 1786
rect 3162 1746 3165 1783
rect 3162 1743 3169 1746
rect 3154 1683 3157 1736
rect 3166 1686 3169 1743
rect 3178 1696 3181 1766
rect 3186 1733 3189 1793
rect 3186 1703 3189 1716
rect 3178 1693 3189 1696
rect 3162 1683 3169 1686
rect 3138 1673 3149 1676
rect 3138 1653 3141 1673
rect 3162 1656 3165 1683
rect 3150 1653 3165 1656
rect 3122 1603 3125 1616
rect 3098 1543 3109 1546
rect 3098 1506 3101 1536
rect 3082 1503 3101 1506
rect 3074 1423 3081 1426
rect 3078 1346 3081 1423
rect 3074 1343 3081 1346
rect 3074 1203 3077 1343
rect 3082 1213 3085 1236
rect 3042 1193 3053 1196
rect 3042 1126 3045 1193
rect 3058 1133 3061 1166
rect 2994 973 3013 976
rect 3018 973 3021 1126
rect 3042 1123 3061 1126
rect 3026 1056 3029 1076
rect 3026 1053 3037 1056
rect 3034 976 3037 1053
rect 3058 1003 3061 1123
rect 3074 1113 3077 1126
rect 3090 1026 3093 1486
rect 3106 1396 3109 1543
rect 3138 1506 3141 1596
rect 3150 1566 3153 1653
rect 3170 1646 3173 1666
rect 3098 1393 3109 1396
rect 3130 1503 3141 1506
rect 3146 1563 3153 1566
rect 3162 1643 3173 1646
rect 3146 1503 3149 1563
rect 3098 1363 3101 1393
rect 3106 1236 3109 1386
rect 3102 1233 3109 1236
rect 3102 1166 3105 1233
rect 3114 1213 3117 1226
rect 3114 1173 3117 1196
rect 3102 1163 3109 1166
rect 3086 1023 3093 1026
rect 3026 973 3037 976
rect 2986 923 2989 936
rect 2858 843 2869 846
rect 2938 873 2953 876
rect 2818 803 2845 806
rect 2818 776 2821 803
rect 2802 773 2821 776
rect 2842 773 2845 803
rect 2726 603 2733 606
rect 2746 603 2749 716
rect 2726 546 2729 603
rect 2726 543 2733 546
rect 2698 523 2709 526
rect 2666 483 2693 486
rect 2618 433 2645 436
rect 2610 423 2621 426
rect 2538 313 2541 403
rect 2546 316 2549 336
rect 2554 333 2557 413
rect 2562 403 2605 406
rect 2562 323 2589 326
rect 2546 313 2553 316
rect 2522 236 2525 313
rect 2550 256 2553 313
rect 2550 253 2557 256
rect 2518 233 2525 236
rect 2518 216 2521 233
rect 2510 213 2521 216
rect 2482 183 2493 186
rect 2466 133 2469 146
rect 2370 113 2405 116
rect 2458 103 2461 126
rect 2474 123 2477 156
rect 2490 116 2493 183
rect 2510 156 2513 213
rect 2510 153 2525 156
rect 2514 123 2517 136
rect 2522 123 2525 153
rect 2482 113 2493 116
rect 2482 43 2485 113
rect 2530 103 2533 226
rect 2546 223 2549 236
rect 2554 223 2557 253
rect 2562 216 2565 323
rect 2538 213 2565 216
rect 2570 213 2573 316
rect 2578 303 2581 316
rect 2602 313 2605 403
rect 2610 326 2613 416
rect 2618 366 2621 423
rect 2626 383 2629 426
rect 2618 363 2629 366
rect 2610 323 2621 326
rect 2610 306 2613 316
rect 2586 303 2613 306
rect 2618 303 2621 323
rect 2626 306 2629 363
rect 2626 303 2637 306
rect 2586 236 2589 303
rect 2586 233 2597 236
rect 2538 196 2541 213
rect 2538 193 2549 196
rect 2546 126 2549 193
rect 2562 133 2565 206
rect 2578 156 2581 226
rect 2570 153 2581 156
rect 2546 123 2565 126
rect 2554 113 2557 123
rect 2562 96 2565 116
rect 2570 103 2573 153
rect 2594 126 2597 233
rect 2578 113 2581 126
rect 2586 123 2597 126
rect 2586 106 2589 123
rect 2610 113 2613 236
rect 2578 103 2589 106
rect 2578 96 2581 103
rect 2562 93 2581 96
rect 2618 96 2621 106
rect 2626 103 2629 296
rect 2634 233 2637 303
rect 2642 296 2645 433
rect 2650 413 2653 436
rect 2658 383 2661 406
rect 2674 393 2677 446
rect 2682 393 2685 406
rect 2690 353 2693 483
rect 2706 456 2709 523
rect 2702 453 2709 456
rect 2650 303 2653 326
rect 2666 313 2669 326
rect 2674 303 2677 316
rect 2642 293 2653 296
rect 2634 113 2637 136
rect 2650 133 2653 293
rect 2690 286 2693 306
rect 2686 283 2693 286
rect 2658 206 2661 226
rect 2658 203 2669 206
rect 2674 203 2677 216
rect 2686 206 2689 283
rect 2702 276 2705 453
rect 2722 446 2725 526
rect 2730 473 2733 543
rect 2722 443 2729 446
rect 2738 443 2741 596
rect 2754 503 2757 773
rect 2762 683 2765 756
rect 2786 733 2789 773
rect 2858 746 2861 843
rect 2874 813 2877 836
rect 2858 743 2869 746
rect 2802 626 2805 646
rect 2794 623 2805 626
rect 2762 593 2765 616
rect 2770 583 2773 606
rect 2794 566 2797 623
rect 2794 563 2805 566
rect 2770 543 2797 546
rect 2698 273 2705 276
rect 2698 213 2701 273
rect 2714 256 2717 436
rect 2726 326 2729 443
rect 2770 413 2773 543
rect 2778 523 2781 536
rect 2794 533 2797 543
rect 2786 516 2789 526
rect 2802 523 2805 563
rect 2810 533 2813 616
rect 2818 516 2821 526
rect 2786 513 2821 516
rect 2826 516 2829 726
rect 2866 723 2869 743
rect 2874 636 2877 806
rect 2898 756 2901 826
rect 2938 766 2941 873
rect 2994 846 2997 973
rect 3002 873 3005 926
rect 3010 906 3013 966
rect 3026 923 3029 973
rect 3058 956 3061 986
rect 3086 976 3089 1023
rect 3098 993 3101 1016
rect 3106 983 3109 1163
rect 3122 1113 3125 1216
rect 3130 1163 3133 1503
rect 3130 1143 3133 1156
rect 3138 1093 3141 1446
rect 3162 1416 3165 1643
rect 3170 1613 3173 1626
rect 3186 1563 3189 1693
rect 3194 1636 3197 1953
rect 3202 1843 3205 1963
rect 3202 1813 3205 1836
rect 3210 1743 3213 1936
rect 3218 1786 3221 2116
rect 3226 2086 3229 2146
rect 3234 2103 3237 2153
rect 3242 2153 3253 2156
rect 3242 2123 3245 2153
rect 3226 2083 3233 2086
rect 3230 2016 3233 2083
rect 3226 2013 3233 2016
rect 3226 1993 3229 2013
rect 3226 1913 3229 1936
rect 3234 1913 3237 1996
rect 3226 1813 3237 1816
rect 3226 1793 3229 1806
rect 3218 1783 3229 1786
rect 3202 1653 3205 1726
rect 3194 1633 3201 1636
rect 3198 1526 3201 1633
rect 3146 1323 3149 1416
rect 3154 1413 3165 1416
rect 3186 1413 3189 1526
rect 3194 1523 3201 1526
rect 3194 1483 3197 1523
rect 3202 1466 3205 1506
rect 3210 1476 3213 1706
rect 3218 1593 3221 1776
rect 3226 1743 3229 1783
rect 3242 1773 3245 2066
rect 3250 2033 3253 2126
rect 3258 2106 3261 2206
rect 3266 2143 3269 2213
rect 3282 2203 3285 2216
rect 3330 2213 3333 2316
rect 3362 2313 3365 2326
rect 3386 2313 3389 2326
rect 3394 2313 3397 2326
rect 3410 2296 3413 2493
rect 3426 2453 3429 2476
rect 3426 2323 3429 2426
rect 3402 2293 3413 2296
rect 3402 2226 3405 2293
rect 3402 2223 3413 2226
rect 3266 2123 3269 2136
rect 3282 2116 3285 2146
rect 3298 2123 3301 2206
rect 3314 2193 3317 2206
rect 3338 2183 3341 2196
rect 3338 2146 3341 2156
rect 3306 2143 3341 2146
rect 3346 2143 3349 2206
rect 3362 2156 3365 2216
rect 3354 2153 3365 2156
rect 3306 2116 3309 2136
rect 3282 2113 3309 2116
rect 3258 2103 3269 2106
rect 3266 2046 3269 2103
rect 3258 2043 3269 2046
rect 3258 2023 3261 2043
rect 3250 1943 3253 2006
rect 3258 1953 3261 2016
rect 3266 2003 3269 2016
rect 3282 2013 3285 2106
rect 3258 1906 3261 1946
rect 3282 1933 3285 1946
rect 3290 1926 3293 2026
rect 3298 1936 3301 2016
rect 3306 1943 3309 1976
rect 3298 1933 3309 1936
rect 3282 1923 3301 1926
rect 3298 1913 3301 1923
rect 3258 1903 3269 1906
rect 3266 1826 3269 1903
rect 3258 1823 3269 1826
rect 3258 1763 3261 1823
rect 3306 1813 3309 1933
rect 3322 1876 3325 2126
rect 3330 2123 3333 2136
rect 3338 2123 3341 2143
rect 3346 1893 3349 2136
rect 3354 2083 3357 2153
rect 3362 2143 3373 2146
rect 3362 2116 3365 2136
rect 3378 2133 3381 2206
rect 3394 2133 3397 2206
rect 3402 2133 3405 2206
rect 3410 2196 3413 2223
rect 3426 2213 3429 2316
rect 3410 2193 3421 2196
rect 3418 2146 3421 2193
rect 3410 2143 3421 2146
rect 3362 2113 3373 2116
rect 3370 2036 3373 2113
rect 3394 2093 3397 2126
rect 3402 2113 3405 2126
rect 3410 2123 3413 2143
rect 3434 2096 3437 2566
rect 3418 2093 3437 2096
rect 3362 2033 3373 2036
rect 3354 1903 3357 1926
rect 3322 1873 3341 1876
rect 3282 1803 3301 1806
rect 3226 1713 3229 1736
rect 3234 1626 3237 1736
rect 3258 1636 3261 1756
rect 3282 1733 3285 1803
rect 3274 1703 3277 1726
rect 3226 1623 3237 1626
rect 3242 1633 3261 1636
rect 3290 1636 3293 1796
rect 3330 1756 3333 1816
rect 3322 1753 3333 1756
rect 3298 1723 3309 1726
rect 3290 1633 3317 1636
rect 3226 1516 3229 1623
rect 3234 1536 3237 1616
rect 3242 1553 3245 1633
rect 3250 1546 3253 1616
rect 3258 1603 3261 1626
rect 3266 1623 3309 1626
rect 3266 1613 3269 1623
rect 3250 1543 3261 1546
rect 3234 1533 3253 1536
rect 3258 1516 3261 1543
rect 3226 1513 3237 1516
rect 3210 1473 3217 1476
rect 3198 1463 3205 1466
rect 3198 1416 3201 1463
rect 3214 1426 3217 1473
rect 3234 1466 3237 1513
rect 3226 1463 3237 1466
rect 3250 1513 3261 1516
rect 3226 1443 3229 1463
rect 3250 1446 3253 1513
rect 3250 1443 3261 1446
rect 3214 1423 3221 1426
rect 3198 1413 3205 1416
rect 3154 1383 3157 1413
rect 3162 1393 3165 1406
rect 3186 1376 3189 1406
rect 3178 1356 3181 1376
rect 3186 1373 3197 1376
rect 3174 1353 3181 1356
rect 3138 1013 3141 1076
rect 3122 976 3125 996
rect 3086 973 3093 976
rect 3122 973 3129 976
rect 3042 953 3061 956
rect 3090 953 3093 973
rect 3010 903 3021 906
rect 2994 843 3005 846
rect 2938 763 2957 766
rect 2890 753 2901 756
rect 2890 733 2893 753
rect 2938 676 2941 726
rect 2946 713 2949 736
rect 2938 673 2949 676
rect 2874 633 2885 636
rect 2882 586 2885 633
rect 2874 583 2885 586
rect 2898 613 2933 616
rect 2866 533 2869 546
rect 2874 516 2877 583
rect 2826 513 2837 516
rect 2810 456 2813 506
rect 2810 453 2817 456
rect 2746 393 2749 406
rect 2710 253 2717 256
rect 2722 323 2729 326
rect 2686 203 2693 206
rect 2642 96 2645 126
rect 2690 113 2693 203
rect 2710 186 2713 253
rect 2722 193 2725 323
rect 2738 313 2741 386
rect 2814 376 2817 453
rect 2834 436 2837 513
rect 2866 513 2877 516
rect 2866 456 2869 513
rect 2866 453 2877 456
rect 2826 433 2837 436
rect 2874 433 2877 453
rect 2826 413 2829 433
rect 2890 426 2893 536
rect 2898 513 2901 613
rect 2914 596 2917 606
rect 2922 603 2933 606
rect 2938 603 2941 616
rect 2946 613 2949 673
rect 2946 596 2949 606
rect 2914 593 2949 596
rect 2906 516 2909 586
rect 2922 533 2925 546
rect 2954 536 2957 763
rect 2962 746 2965 826
rect 2978 783 2981 806
rect 3002 803 3005 843
rect 3018 836 3021 903
rect 3042 856 3045 953
rect 3058 933 3061 953
rect 3042 853 3049 856
rect 3010 833 3021 836
rect 3010 786 3013 833
rect 3010 783 3021 786
rect 2962 743 3005 746
rect 2962 696 2965 736
rect 2970 713 2973 726
rect 2986 706 2989 726
rect 2982 703 2989 706
rect 2962 693 2973 696
rect 2970 626 2973 693
rect 2962 623 2973 626
rect 2962 603 2965 623
rect 2982 606 2985 703
rect 2994 613 2997 736
rect 3002 723 3005 743
rect 3010 706 3013 776
rect 3006 703 3013 706
rect 2978 603 2985 606
rect 3006 606 3009 703
rect 3006 603 3013 606
rect 2962 583 2965 596
rect 2978 586 2981 603
rect 2978 583 2989 586
rect 3010 583 3013 603
rect 2938 533 2957 536
rect 2906 513 2917 516
rect 2914 436 2917 513
rect 2938 463 2941 533
rect 2946 486 2949 526
rect 2962 523 2973 526
rect 2962 486 2965 523
rect 2946 483 2965 486
rect 2978 446 2981 536
rect 2986 513 2989 583
rect 2994 523 2997 536
rect 3010 456 3013 536
rect 3018 513 3021 783
rect 3026 776 3029 816
rect 3046 806 3049 853
rect 3058 813 3061 916
rect 3106 846 3109 926
rect 3126 856 3129 973
rect 3138 893 3141 926
rect 3146 913 3149 1236
rect 3154 1216 3157 1346
rect 3174 1306 3177 1353
rect 3186 1313 3189 1326
rect 3174 1303 3181 1306
rect 3162 1223 3165 1236
rect 3154 1213 3165 1216
rect 3170 1213 3173 1226
rect 3154 1103 3157 1126
rect 3162 1123 3165 1213
rect 3178 1143 3181 1303
rect 3186 1213 3189 1226
rect 3194 1193 3197 1373
rect 3202 1323 3205 1413
rect 3218 1346 3221 1423
rect 3250 1413 3253 1426
rect 3234 1383 3237 1396
rect 3210 1343 3221 1346
rect 3202 1213 3205 1226
rect 3170 1113 3173 1136
rect 3186 1133 3189 1156
rect 3194 1106 3197 1126
rect 3202 1113 3205 1186
rect 3186 1103 3197 1106
rect 3186 1036 3189 1103
rect 3170 1013 3173 1036
rect 3178 1033 3189 1036
rect 3170 933 3173 996
rect 3178 906 3181 1033
rect 3202 1026 3205 1096
rect 3210 1033 3213 1343
rect 3218 1223 3221 1236
rect 3234 1216 3237 1356
rect 3242 1333 3245 1406
rect 3250 1233 3253 1406
rect 3258 1403 3261 1443
rect 3258 1383 3261 1396
rect 3266 1373 3269 1606
rect 3274 1563 3277 1606
rect 3282 1593 3285 1606
rect 3266 1333 3269 1346
rect 3266 1313 3269 1326
rect 3274 1226 3277 1556
rect 3282 1353 3285 1546
rect 3290 1536 3293 1616
rect 3298 1593 3301 1606
rect 3306 1543 3309 1623
rect 3314 1553 3317 1633
rect 3322 1603 3325 1753
rect 3338 1663 3341 1873
rect 3346 1803 3349 1886
rect 3362 1733 3365 2033
rect 3418 1956 3421 2093
rect 3418 1953 3437 1956
rect 3402 1913 3405 1926
rect 3410 1923 3429 1926
rect 3434 1906 3437 1953
rect 3362 1656 3365 1726
rect 3330 1653 3365 1656
rect 3330 1596 3333 1653
rect 3346 1603 3349 1616
rect 3322 1593 3333 1596
rect 3322 1543 3325 1593
rect 3290 1533 3317 1536
rect 3290 1503 3293 1526
rect 3306 1426 3309 1526
rect 3298 1423 3309 1426
rect 3290 1403 3293 1416
rect 3290 1336 3293 1396
rect 3314 1383 3317 1533
rect 3322 1413 3325 1526
rect 3322 1393 3325 1406
rect 3330 1366 3333 1586
rect 3322 1363 3333 1366
rect 3290 1333 3309 1336
rect 3298 1306 3301 1326
rect 3290 1303 3301 1306
rect 3290 1246 3293 1303
rect 3290 1243 3301 1246
rect 3274 1223 3281 1226
rect 3226 1213 3237 1216
rect 3226 1156 3229 1213
rect 3266 1183 3269 1216
rect 3278 1176 3281 1223
rect 3218 1153 3229 1156
rect 3274 1173 3281 1176
rect 3194 1013 3197 1026
rect 3202 1023 3209 1026
rect 3186 963 3189 1006
rect 3186 923 3189 956
rect 3194 906 3197 1006
rect 3206 966 3209 1023
rect 3218 976 3221 1153
rect 3274 1146 3277 1173
rect 3258 1143 3277 1146
rect 3226 1023 3229 1136
rect 3234 1086 3237 1116
rect 3242 1103 3245 1126
rect 3250 1113 3253 1136
rect 3258 1093 3261 1143
rect 3234 1083 3241 1086
rect 3238 1016 3241 1083
rect 3234 1013 3241 1016
rect 3218 973 3225 976
rect 3206 963 3213 966
rect 3210 943 3213 963
rect 3170 903 3181 906
rect 3190 903 3197 906
rect 3126 853 3133 856
rect 3106 843 3117 846
rect 3106 823 3109 836
rect 3114 826 3117 843
rect 3114 823 3121 826
rect 3042 803 3049 806
rect 3042 783 3045 803
rect 3066 776 3069 806
rect 3026 773 3069 776
rect 3026 756 3029 773
rect 3026 753 3033 756
rect 3030 656 3033 753
rect 3066 713 3069 726
rect 3090 703 3093 816
rect 3118 766 3121 823
rect 3114 763 3121 766
rect 3026 653 3033 656
rect 3026 546 3029 653
rect 3034 613 3037 636
rect 3098 633 3101 736
rect 3114 733 3117 763
rect 3130 746 3133 853
rect 3170 826 3173 903
rect 3190 836 3193 903
rect 3190 833 3197 836
rect 3146 806 3149 826
rect 3170 823 3181 826
rect 3122 743 3133 746
rect 3142 803 3149 806
rect 3122 693 3125 743
rect 3142 676 3145 803
rect 3154 686 3157 806
rect 3162 733 3165 796
rect 3178 733 3181 823
rect 3194 816 3197 833
rect 3202 823 3205 936
rect 3194 813 3205 816
rect 3186 803 3205 806
rect 3186 793 3189 803
rect 3170 713 3173 726
rect 3178 693 3181 726
rect 3202 703 3205 716
rect 3210 686 3213 936
rect 3222 846 3225 973
rect 3234 906 3237 1013
rect 3242 913 3245 926
rect 3250 923 3253 1046
rect 3258 993 3261 1006
rect 3258 906 3261 986
rect 3266 966 3269 1136
rect 3282 1133 3285 1156
rect 3290 1143 3293 1226
rect 3298 1216 3301 1243
rect 3306 1236 3309 1316
rect 3322 1256 3325 1363
rect 3338 1323 3341 1556
rect 3346 1516 3349 1546
rect 3362 1533 3365 1576
rect 3346 1513 3357 1516
rect 3354 1446 3357 1513
rect 3378 1503 3381 1886
rect 3410 1816 3413 1906
rect 3426 1903 3437 1906
rect 3426 1826 3429 1903
rect 3426 1823 3437 1826
rect 3394 1763 3397 1816
rect 3406 1813 3413 1816
rect 3406 1716 3409 1813
rect 3418 1723 3421 1806
rect 3434 1753 3437 1823
rect 3406 1713 3413 1716
rect 3394 1593 3397 1616
rect 3410 1566 3413 1713
rect 3406 1563 3413 1566
rect 3418 1566 3421 1616
rect 3426 1573 3429 1616
rect 3418 1563 3429 1566
rect 3346 1443 3357 1446
rect 3346 1403 3349 1443
rect 3394 1426 3397 1526
rect 3406 1446 3409 1563
rect 3406 1443 3413 1446
rect 3354 1393 3357 1406
rect 3346 1323 3349 1336
rect 3362 1333 3365 1426
rect 3378 1383 3381 1416
rect 3386 1403 3389 1426
rect 3394 1423 3405 1426
rect 3410 1423 3413 1443
rect 3394 1336 3397 1416
rect 3402 1403 3405 1423
rect 3402 1356 3405 1396
rect 3418 1383 3421 1526
rect 3426 1366 3429 1563
rect 3422 1363 3429 1366
rect 3402 1353 3413 1356
rect 3370 1286 3373 1336
rect 3386 1333 3397 1336
rect 3338 1283 3373 1286
rect 3338 1266 3341 1283
rect 3338 1263 3349 1266
rect 3322 1253 3333 1256
rect 3306 1233 3317 1236
rect 3330 1233 3333 1253
rect 3314 1226 3317 1233
rect 3314 1223 3333 1226
rect 3298 1213 3309 1216
rect 3298 1193 3301 1206
rect 3290 1133 3301 1136
rect 3274 1123 3285 1126
rect 3290 1113 3293 1126
rect 3298 1106 3301 1133
rect 3306 1123 3309 1213
rect 3322 1196 3325 1216
rect 3318 1193 3325 1196
rect 3318 1126 3321 1193
rect 3318 1123 3325 1126
rect 3298 1103 3305 1106
rect 3274 986 3277 1096
rect 3290 1013 3293 1096
rect 3302 1036 3305 1103
rect 3298 1033 3305 1036
rect 3298 1016 3301 1033
rect 3298 1013 3309 1016
rect 3282 1003 3309 1006
rect 3314 1003 3317 1106
rect 3322 1093 3325 1123
rect 3274 983 3285 986
rect 3266 963 3273 966
rect 3234 903 3245 906
rect 3154 683 3161 686
rect 3138 673 3145 676
rect 3138 626 3141 673
rect 3158 636 3161 683
rect 3206 683 3213 686
rect 3218 843 3225 846
rect 3154 633 3161 636
rect 3138 623 3149 626
rect 3042 603 3053 606
rect 3026 543 3037 546
rect 3002 453 3013 456
rect 2978 443 2985 446
rect 2906 433 2917 436
rect 2858 423 2893 426
rect 2858 406 2861 423
rect 2810 373 2817 376
rect 2730 223 2733 306
rect 2746 293 2749 336
rect 2754 303 2757 326
rect 2746 233 2773 236
rect 2746 213 2749 233
rect 2762 216 2765 226
rect 2754 213 2765 216
rect 2770 213 2773 233
rect 2710 183 2717 186
rect 2698 123 2701 136
rect 2618 93 2645 96
rect 2714 73 2717 183
rect 2738 106 2741 206
rect 2746 113 2749 136
rect 2754 123 2757 213
rect 2778 203 2781 356
rect 2810 333 2813 373
rect 2842 286 2845 406
rect 2854 403 2861 406
rect 2854 346 2857 403
rect 2866 396 2869 416
rect 2874 413 2885 416
rect 2890 403 2893 416
rect 2898 396 2901 426
rect 2906 416 2909 433
rect 2906 413 2917 416
rect 2866 393 2901 396
rect 2954 393 2957 406
rect 2982 396 2985 443
rect 2978 393 2985 396
rect 2854 343 2861 346
rect 2858 323 2861 343
rect 2930 333 2933 356
rect 2786 133 2789 286
rect 2810 283 2845 286
rect 2890 283 2893 326
rect 2978 323 2981 393
rect 2994 366 2997 416
rect 3002 413 3005 453
rect 3026 446 3029 536
rect 3034 503 3037 543
rect 3042 533 3045 546
rect 3058 523 3061 616
rect 3074 593 3077 616
rect 3074 506 3077 566
rect 3090 546 3093 616
rect 3098 603 3101 616
rect 3114 583 3117 616
rect 3146 603 3149 623
rect 3154 603 3157 633
rect 3186 623 3189 636
rect 3090 543 3101 546
rect 3090 516 3093 536
rect 3066 503 3077 506
rect 3086 513 3093 516
rect 3098 513 3101 543
rect 3106 523 3109 536
rect 3122 523 3125 536
rect 3018 443 3029 446
rect 3066 446 3069 503
rect 3066 443 3077 446
rect 3026 413 3037 416
rect 3066 403 3069 416
rect 3074 413 3077 443
rect 3086 426 3089 513
rect 3082 423 3089 426
rect 2994 363 3005 366
rect 3002 286 3005 363
rect 3050 333 3053 356
rect 2978 283 3005 286
rect 2810 203 2813 283
rect 2906 233 2933 236
rect 2858 203 2861 226
rect 2866 183 2869 206
rect 2890 203 2893 216
rect 2906 213 2909 233
rect 2922 216 2925 226
rect 2914 213 2925 216
rect 2930 213 2933 233
rect 2858 143 2893 146
rect 2858 133 2861 143
rect 2762 106 2765 116
rect 2810 113 2813 126
rect 2866 113 2869 136
rect 2874 123 2877 136
rect 2890 123 2893 143
rect 2906 123 2909 136
rect 2914 123 2917 213
rect 2922 193 2925 206
rect 2738 103 2765 106
rect 2922 93 2925 186
rect 2930 133 2933 206
rect 2978 203 2981 283
rect 3034 236 3037 326
rect 3082 323 3085 423
rect 3098 413 3101 506
rect 3130 483 3133 536
rect 3138 513 3141 526
rect 3114 393 3117 406
rect 3146 396 3149 416
rect 3142 393 3149 396
rect 3130 236 3133 326
rect 3142 316 3145 393
rect 3142 313 3149 316
rect 3154 313 3157 536
rect 3162 523 3165 616
rect 3186 593 3189 606
rect 3194 603 3197 616
rect 3206 576 3209 683
rect 3218 643 3221 843
rect 3226 806 3229 826
rect 3226 803 3233 806
rect 3230 676 3233 803
rect 3226 673 3233 676
rect 3226 653 3229 673
rect 3218 583 3221 626
rect 3194 573 3209 576
rect 3170 523 3173 536
rect 3194 436 3197 573
rect 3218 543 3221 556
rect 3226 543 3229 606
rect 3194 433 3213 436
rect 3162 413 3165 426
rect 3186 413 3197 416
rect 3210 396 3213 433
rect 3218 423 3221 536
rect 3234 523 3237 536
rect 3242 533 3245 903
rect 3254 903 3261 906
rect 3254 826 3257 903
rect 3270 896 3273 963
rect 3266 893 3273 896
rect 3254 823 3261 826
rect 3258 803 3261 823
rect 3258 783 3261 796
rect 3266 766 3269 893
rect 3262 763 3269 766
rect 3250 713 3253 736
rect 3262 706 3265 763
rect 3282 756 3285 983
rect 3298 813 3301 826
rect 3298 783 3301 806
rect 3258 703 3265 706
rect 3274 753 3285 756
rect 3258 623 3261 703
rect 3274 666 3277 753
rect 3282 703 3285 716
rect 3306 686 3309 1003
rect 3322 973 3325 996
rect 3314 913 3317 926
rect 3322 923 3325 936
rect 3322 803 3325 916
rect 3314 783 3317 796
rect 3298 683 3309 686
rect 3274 663 3285 666
rect 3258 526 3261 536
rect 3250 523 3261 526
rect 3250 516 3253 523
rect 3226 513 3253 516
rect 3266 513 3269 656
rect 3282 566 3285 663
rect 3298 613 3301 683
rect 3322 626 3325 726
rect 3330 696 3333 1216
rect 3346 1176 3349 1263
rect 3386 1233 3389 1326
rect 3338 1173 3349 1176
rect 3338 913 3341 1173
rect 3362 1133 3365 1226
rect 3386 1223 3397 1226
rect 3386 1206 3389 1223
rect 3378 1203 3389 1206
rect 3354 1043 3357 1126
rect 3362 1103 3365 1116
rect 3370 1113 3373 1126
rect 3378 1113 3381 1203
rect 3402 1126 3405 1336
rect 3410 1323 3413 1353
rect 3422 1306 3425 1363
rect 3418 1303 3425 1306
rect 3418 1136 3421 1303
rect 3418 1133 3425 1136
rect 3386 1113 3389 1126
rect 3394 1123 3405 1126
rect 3346 1013 3349 1026
rect 3354 993 3357 1006
rect 3362 983 3365 1036
rect 3378 1023 3381 1106
rect 3402 1096 3405 1116
rect 3394 1093 3405 1096
rect 3394 1016 3397 1093
rect 3378 1003 3381 1016
rect 3394 1013 3405 1016
rect 3346 913 3349 936
rect 3394 896 3397 996
rect 3386 893 3397 896
rect 3386 836 3389 893
rect 3338 813 3341 826
rect 3338 783 3341 806
rect 3354 733 3357 836
rect 3386 833 3397 836
rect 3402 833 3405 1013
rect 3410 1006 3413 1116
rect 3422 1056 3425 1133
rect 3422 1053 3429 1056
rect 3418 1013 3421 1036
rect 3410 1003 3417 1006
rect 3414 946 3417 1003
rect 3414 943 3421 946
rect 3410 903 3413 926
rect 3418 913 3421 943
rect 3394 816 3397 833
rect 3378 813 3389 816
rect 3394 813 3405 816
rect 3410 813 3413 826
rect 3378 793 3381 813
rect 3418 806 3421 816
rect 3410 803 3421 806
rect 3338 703 3341 726
rect 3362 716 3365 736
rect 3362 713 3373 716
rect 3330 693 3337 696
rect 3314 623 3325 626
rect 3274 563 3285 566
rect 3274 523 3277 563
rect 3298 546 3301 606
rect 3314 586 3317 606
rect 3282 543 3301 546
rect 3310 583 3317 586
rect 3258 413 3261 486
rect 3282 456 3285 543
rect 3274 453 3285 456
rect 3210 393 3221 396
rect 3234 393 3237 406
rect 3274 396 3277 453
rect 3274 393 3285 396
rect 3218 386 3221 393
rect 3218 383 3229 386
rect 3194 333 3197 356
rect 3146 296 3149 313
rect 3226 306 3229 383
rect 3282 376 3285 393
rect 3242 373 3285 376
rect 3242 323 3245 373
rect 3226 303 3237 306
rect 3146 293 3157 296
rect 3034 233 3045 236
rect 3026 203 3029 226
rect 3042 186 3045 233
rect 3066 203 3069 216
rect 3090 203 3093 236
rect 3098 233 3133 236
rect 2930 113 2933 126
rect 2954 106 2957 186
rect 3002 183 3045 186
rect 3098 183 3101 233
rect 3154 226 3157 293
rect 3146 223 3157 226
rect 3178 223 3181 236
rect 3146 203 3149 223
rect 3194 193 3197 236
rect 3202 206 3205 226
rect 3202 203 3213 206
rect 2978 113 2981 126
rect 2986 106 2989 126
rect 3002 123 3005 183
rect 3074 143 3109 146
rect 3074 133 3077 143
rect 2954 103 2989 106
rect 3090 93 3093 136
rect 3098 116 3101 126
rect 3106 123 3109 143
rect 3122 133 3125 146
rect 3098 113 3125 116
rect 3146 93 3149 136
rect 3218 133 3221 296
rect 3234 226 3237 303
rect 3274 236 3277 326
rect 3226 223 3237 226
rect 3250 233 3277 236
rect 3226 203 3229 223
rect 3250 216 3253 233
rect 3246 213 3253 216
rect 3246 156 3249 213
rect 3246 153 3253 156
rect 3250 136 3253 153
rect 3234 133 3253 136
rect 3186 123 3253 126
rect 3258 116 3261 216
rect 3298 213 3301 526
rect 3310 516 3313 583
rect 3322 563 3325 616
rect 3334 556 3337 693
rect 3346 613 3349 696
rect 3370 646 3373 713
rect 3402 706 3405 726
rect 3394 703 3405 706
rect 3394 656 3397 703
rect 3394 653 3405 656
rect 3362 643 3373 646
rect 3346 593 3349 606
rect 3334 553 3341 556
rect 3310 513 3317 516
rect 3322 513 3325 536
rect 3314 426 3317 513
rect 3330 503 3333 536
rect 3338 513 3341 553
rect 3362 546 3365 643
rect 3394 546 3397 616
rect 3402 603 3405 653
rect 3410 613 3413 626
rect 3346 543 3365 546
rect 3346 523 3349 543
rect 3362 533 3365 543
rect 3378 523 3381 546
rect 3394 543 3413 546
rect 3418 543 3421 726
rect 3378 503 3381 516
rect 3314 423 3325 426
rect 3306 413 3317 416
rect 3322 356 3325 423
rect 3386 413 3389 536
rect 3402 523 3405 536
rect 3410 516 3413 543
rect 3410 513 3421 516
rect 3418 413 3421 496
rect 3338 393 3341 406
rect 3314 353 3325 356
rect 3314 286 3317 353
rect 3338 333 3341 356
rect 3386 323 3389 406
rect 3426 393 3429 1053
rect 3434 563 3437 1506
rect 3434 403 3437 536
rect 3314 283 3349 286
rect 3322 213 3341 216
rect 3314 133 3317 206
rect 3322 193 3325 206
rect 3330 193 3333 206
rect 3346 203 3349 283
rect 3418 236 3421 326
rect 3370 233 3421 236
rect 3354 196 3357 216
rect 3346 193 3357 196
rect 3250 113 3261 116
rect 3250 93 3253 113
rect 3322 93 3325 136
rect 3346 133 3349 193
rect 3370 136 3373 233
rect 3354 133 3373 136
rect 3330 113 3333 126
rect 3370 93 3373 116
rect 3378 113 3381 126
rect 3426 123 3429 206
rect 3434 203 3437 216
rect 3446 37 3466 3303
rect 3470 13 3490 3327
<< metal3 >>
rect 1409 3332 1630 3337
rect 1409 3327 1414 3332
rect 505 3322 582 3327
rect 913 3322 966 3327
rect 1385 3322 1414 3327
rect 1625 3327 1630 3332
rect 1625 3322 1806 3327
rect 2361 3322 2590 3327
rect 2689 3322 3110 3327
rect 1425 3312 1454 3317
rect 1449 3307 1454 3312
rect 1529 3312 1622 3317
rect 1529 3307 1534 3312
rect 497 3302 726 3307
rect 1449 3302 1534 3307
rect 713 3292 1166 3297
rect 929 3272 1094 3277
rect 929 3267 934 3272
rect 537 3262 734 3267
rect 753 3262 886 3267
rect 905 3262 934 3267
rect 753 3257 758 3262
rect 673 3252 758 3257
rect 881 3257 886 3262
rect 953 3257 1046 3262
rect 881 3252 958 3257
rect 1041 3252 1070 3257
rect 1089 3247 1094 3272
rect 1961 3272 2118 3277
rect 1793 3262 1918 3267
rect 1793 3257 1798 3262
rect 1201 3252 1406 3257
rect 1769 3252 1798 3257
rect 1913 3257 1918 3262
rect 1961 3257 1966 3272
rect 2113 3257 2118 3272
rect 2665 3272 2846 3277
rect 2345 3262 2454 3267
rect 2473 3262 2582 3267
rect 2473 3257 2478 3262
rect 1913 3252 1966 3257
rect 2009 3252 2078 3257
rect 2113 3252 2166 3257
rect 2401 3252 2478 3257
rect 2577 3257 2582 3262
rect 2665 3257 2670 3272
rect 2577 3252 2606 3257
rect 2641 3252 2670 3257
rect 2841 3257 2846 3272
rect 2841 3252 2990 3257
rect 2009 3247 2014 3252
rect 921 3242 1078 3247
rect 1089 3242 1166 3247
rect 1185 3242 1302 3247
rect 1649 3242 1870 3247
rect 1937 3242 2014 3247
rect 2073 3247 2078 3252
rect 2073 3242 2102 3247
rect 2257 3242 2414 3247
rect 2457 3242 2854 3247
rect 681 3237 766 3242
rect 1937 3237 1942 3242
rect 561 3232 686 3237
rect 761 3232 910 3237
rect 929 3232 966 3237
rect 1081 3232 1310 3237
rect 1377 3232 1510 3237
rect 1561 3232 1942 3237
rect 1953 3232 2070 3237
rect 2297 3232 2470 3237
rect 2481 3232 2550 3237
rect 2609 3232 2662 3237
rect 2825 3232 2910 3237
rect 2977 3232 3022 3237
rect 489 3222 598 3227
rect 697 3222 806 3227
rect 817 3222 854 3227
rect 945 3222 1150 3227
rect 1249 3222 1582 3227
rect 1705 3222 2126 3227
rect 2177 3222 2454 3227
rect 2593 3222 2782 3227
rect 1169 3217 1254 3222
rect 1577 3217 1710 3222
rect 1121 3212 1174 3217
rect 1265 3212 1558 3217
rect 1729 3212 1766 3217
rect 1785 3212 1918 3217
rect 2033 3212 2326 3217
rect 2473 3212 2542 3217
rect 1729 3207 1734 3212
rect 2473 3207 2478 3212
rect 129 3202 206 3207
rect 633 3202 702 3207
rect 769 3202 942 3207
rect 1169 3202 1734 3207
rect 1745 3202 2030 3207
rect 2073 3202 2318 3207
rect 2433 3202 2478 3207
rect 2537 3207 2542 3212
rect 2977 3207 2982 3232
rect 2537 3202 2590 3207
rect 2673 3202 2846 3207
rect 2977 3202 2998 3207
rect 129 3197 134 3202
rect 81 3192 134 3197
rect 201 3197 206 3202
rect 1169 3197 1174 3202
rect 2673 3197 2678 3202
rect 201 3192 230 3197
rect 305 3192 414 3197
rect 449 3192 598 3197
rect 681 3192 710 3197
rect 993 3192 1174 3197
rect 1193 3192 1886 3197
rect 1921 3192 1966 3197
rect 2001 3192 2094 3197
rect 2169 3192 2278 3197
rect 2289 3192 2678 3197
rect 2953 3192 3046 3197
rect 3081 3192 3230 3197
rect 3305 3192 3358 3197
rect 865 3187 950 3192
rect 2001 3187 2006 3192
rect 3081 3187 3086 3192
rect 641 3182 718 3187
rect 753 3182 870 3187
rect 945 3182 1038 3187
rect 1105 3182 1382 3187
rect 1417 3182 1462 3187
rect 1473 3182 1598 3187
rect 1753 3182 1886 3187
rect 1881 3177 1886 3182
rect 1953 3182 2006 3187
rect 2017 3182 2270 3187
rect 2305 3182 2358 3187
rect 2369 3182 2510 3187
rect 2537 3182 2646 3187
rect 2673 3182 2822 3187
rect 2977 3182 3086 3187
rect 3225 3187 3230 3192
rect 3225 3182 3366 3187
rect 1953 3177 1958 3182
rect 145 3172 174 3177
rect 169 3167 174 3172
rect 233 3172 318 3177
rect 785 3172 854 3177
rect 865 3172 934 3177
rect 1025 3172 1702 3177
rect 1881 3172 1958 3177
rect 2081 3172 2438 3177
rect 2617 3172 2662 3177
rect 2873 3172 2990 3177
rect 3369 3172 3438 3177
rect 233 3167 238 3172
rect 2657 3167 2662 3172
rect 169 3162 238 3167
rect 481 3162 518 3167
rect 793 3162 894 3167
rect 1041 3162 1078 3167
rect 1169 3162 1462 3167
rect 1481 3162 1566 3167
rect 2001 3162 2094 3167
rect 2201 3162 2630 3167
rect 2657 3162 2686 3167
rect 2737 3162 2822 3167
rect 2833 3162 3214 3167
rect 1169 3157 1174 3162
rect 385 3152 438 3157
rect 505 3152 686 3157
rect 713 3152 958 3157
rect 1009 3152 1174 3157
rect 1193 3152 1430 3157
rect 1521 3152 1678 3157
rect 1889 3152 1974 3157
rect 2009 3152 2190 3157
rect 2297 3152 2366 3157
rect 2409 3152 2622 3157
rect 2721 3152 2774 3157
rect 1521 3147 1526 3152
rect 1889 3147 1894 3152
rect 417 3142 582 3147
rect 705 3142 774 3147
rect 833 3142 918 3147
rect 945 3142 982 3147
rect 1033 3142 1366 3147
rect 1417 3142 1526 3147
rect 1641 3142 1750 3147
rect 1865 3142 1894 3147
rect 1977 3142 2278 3147
rect 2329 3142 2374 3147
rect 2457 3142 2518 3147
rect 2737 3142 2766 3147
rect 2737 3137 2742 3142
rect 137 3132 270 3137
rect 361 3132 454 3137
rect 577 3132 718 3137
rect 833 3132 894 3137
rect 929 3132 1214 3137
rect 1313 3132 1486 3137
rect 1553 3132 1814 3137
rect 1841 3132 2030 3137
rect 2097 3132 2150 3137
rect 2201 3132 2390 3137
rect 2641 3132 2742 3137
rect 2817 3137 2822 3162
rect 3209 3157 3214 3162
rect 3305 3162 3350 3167
rect 3305 3157 3310 3162
rect 2945 3152 2966 3157
rect 3209 3152 3310 3157
rect 3345 3157 3350 3162
rect 3345 3152 3406 3157
rect 2817 3132 2894 3137
rect 713 3127 838 3132
rect 545 3122 694 3127
rect 1033 3122 1414 3127
rect 1545 3122 1646 3127
rect 1681 3122 1806 3127
rect 1937 3122 2270 3127
rect 2505 3122 2598 3127
rect 2609 3122 2694 3127
rect 73 3112 126 3117
rect 121 3107 126 3112
rect 201 3112 230 3117
rect 393 3112 470 3117
rect 489 3112 598 3117
rect 201 3107 206 3112
rect 265 3107 334 3112
rect 393 3107 398 3112
rect 121 3102 206 3107
rect 241 3102 270 3107
rect 329 3102 398 3107
rect 465 3107 470 3112
rect 689 3107 694 3122
rect 857 3117 1014 3122
rect 1433 3117 1526 3122
rect 2369 3117 2486 3122
rect 713 3112 862 3117
rect 1009 3112 1094 3117
rect 1305 3112 1438 3117
rect 1521 3112 1638 3117
rect 2065 3112 2286 3117
rect 2345 3112 2374 3117
rect 2481 3112 2566 3117
rect 1153 3107 1286 3112
rect 465 3102 550 3107
rect 561 3102 662 3107
rect 689 3102 782 3107
rect 873 3102 1110 3107
rect 1129 3102 1158 3107
rect 1281 3102 1326 3107
rect 1449 3102 1574 3107
rect 1769 3102 1894 3107
rect 2249 3102 2430 3107
rect 2489 3102 2582 3107
rect 2609 3102 2614 3122
rect 2945 3117 2950 3152
rect 2969 3142 3038 3147
rect 3105 3132 3190 3137
rect 2841 3112 2950 3117
rect 3193 3112 3238 3117
rect 2881 3102 3038 3107
rect 561 3097 566 3102
rect 777 3097 878 3102
rect 289 3092 318 3097
rect 537 3092 566 3097
rect 657 3092 758 3097
rect 897 3092 1062 3097
rect 1073 3092 1342 3097
rect 1553 3092 1870 3097
rect 1881 3092 2054 3097
rect 313 3087 318 3092
rect 409 3087 542 3092
rect 313 3082 414 3087
rect 569 3082 678 3087
rect 801 3082 878 3087
rect 985 3082 1214 3087
rect 1345 3082 1446 3087
rect 2457 3082 2510 3087
rect 801 3077 806 3082
rect 873 3077 966 3082
rect 1657 3077 1774 3082
rect 433 3072 630 3077
rect 777 3072 806 3077
rect 961 3072 1318 3077
rect 1329 3072 1358 3077
rect 1633 3072 1662 3077
rect 1769 3072 1870 3077
rect 1953 3072 2022 3077
rect 2417 3072 2478 3077
rect 625 3067 758 3072
rect 1313 3067 1318 3072
rect 1953 3067 1958 3072
rect 753 3062 1094 3067
rect 1113 3062 1142 3067
rect 1313 3062 1478 3067
rect 1569 3062 1782 3067
rect 1849 3062 1958 3067
rect 2745 3062 2830 3067
rect 2745 3057 2750 3062
rect 241 3052 350 3057
rect 585 3052 678 3057
rect 705 3052 798 3057
rect 1001 3052 1270 3057
rect 1617 3052 1726 3057
rect 1897 3052 2134 3057
rect 241 3047 246 3052
rect 217 3042 246 3047
rect 345 3047 350 3052
rect 1417 3047 1510 3052
rect 2129 3047 2134 3052
rect 2153 3052 2278 3057
rect 2553 3052 2750 3057
rect 2825 3057 2830 3062
rect 2825 3052 2942 3057
rect 2153 3047 2158 3052
rect 345 3042 406 3047
rect 625 3042 726 3047
rect 809 3042 1030 3047
rect 1049 3042 1206 3047
rect 1273 3042 1422 3047
rect 1505 3042 1534 3047
rect 1545 3042 1582 3047
rect 1625 3042 1846 3047
rect 2129 3042 2158 3047
rect 2273 3047 2278 3052
rect 2273 3042 2302 3047
rect 2689 3042 2718 3047
rect 2873 3042 2950 3047
rect 721 3037 814 3042
rect 2713 3037 2798 3042
rect 2873 3037 2878 3042
rect 153 3032 262 3037
rect 625 3032 702 3037
rect 1105 3032 1270 3037
rect 1433 3032 1542 3037
rect 1657 3032 1718 3037
rect 1881 3032 1950 3037
rect 1969 3032 2110 3037
rect 833 3027 990 3032
rect 1969 3027 1974 3032
rect 321 3022 430 3027
rect 449 3022 470 3027
rect 513 3022 574 3027
rect 665 3022 838 3027
rect 985 3022 1014 3027
rect 1097 3022 1254 3027
rect 1313 3022 1390 3027
rect 1409 3022 1630 3027
rect 1649 3022 1910 3027
rect 1929 3022 1974 3027
rect 2105 3027 2110 3032
rect 2321 3032 2398 3037
rect 2449 3032 2558 3037
rect 2793 3032 2878 3037
rect 3249 3032 3278 3037
rect 2321 3027 2326 3032
rect 2105 3022 2326 3027
rect 2393 3027 2398 3032
rect 2393 3022 2502 3027
rect 2665 3022 2774 3027
rect 1313 3017 1318 3022
rect 257 3012 310 3017
rect 537 3012 958 3017
rect 1241 3012 1318 3017
rect 1385 3017 1390 3022
rect 1385 3012 1422 3017
rect 1521 3012 1694 3017
rect 1833 3012 2142 3017
rect 2241 3012 2446 3017
rect 305 3007 310 3012
rect 377 3007 542 3012
rect 977 3007 1102 3012
rect 1689 3007 1838 3012
rect 3249 3007 3254 3032
rect 3265 3022 3358 3027
rect 305 3002 382 3007
rect 561 3002 982 3007
rect 1097 3002 1126 3007
rect 1137 3002 1222 3007
rect 1329 3002 1590 3007
rect 1969 3002 2046 3007
rect 2369 3002 2454 3007
rect 2465 3002 2566 3007
rect 3049 3002 3078 3007
rect 3097 3002 3174 3007
rect 3249 3002 3286 3007
rect 1137 2997 1142 3002
rect 2449 2997 2454 3002
rect 3097 2997 3102 3002
rect 137 2992 238 2997
rect 401 2992 454 2997
rect 521 2992 662 2997
rect 801 2992 870 2997
rect 889 2992 982 2997
rect 1041 2992 1142 2997
rect 1185 2992 1270 2997
rect 1281 2992 1310 2997
rect 1321 2992 1542 2997
rect 1625 2992 1718 2997
rect 1825 2992 1918 2997
rect 2001 2992 2070 2997
rect 2193 2992 2326 2997
rect 2449 2992 2830 2997
rect 2945 2992 3038 2997
rect 3057 2992 3102 2997
rect 3169 2997 3174 3002
rect 3169 2992 3198 2997
rect 449 2987 454 2992
rect 801 2987 806 2992
rect 1281 2987 1286 2992
rect 89 2982 438 2987
rect 449 2982 566 2987
rect 641 2982 806 2987
rect 857 2982 1150 2987
rect 1249 2982 1286 2987
rect 1537 2987 1542 2992
rect 1537 2982 1670 2987
rect 1681 2982 1886 2987
rect 1937 2982 1982 2987
rect 2225 2982 2342 2987
rect 2521 2982 2558 2987
rect 2969 2982 3166 2987
rect 1937 2977 1942 2982
rect 449 2972 606 2977
rect 985 2972 1526 2977
rect 105 2967 222 2972
rect 321 2967 398 2972
rect 1521 2967 1526 2972
rect 1625 2972 1670 2977
rect 1689 2972 1942 2977
rect 1953 2972 2526 2977
rect 2737 2972 3222 2977
rect 1625 2967 1630 2972
rect 81 2962 110 2967
rect 217 2962 326 2967
rect 393 2962 550 2967
rect 673 2962 806 2967
rect 865 2962 974 2967
rect 1065 2962 1094 2967
rect 1217 2962 1462 2967
rect 1521 2962 1630 2967
rect 1665 2967 1670 2972
rect 1665 2962 1830 2967
rect 1905 2962 2238 2967
rect 2281 2962 2358 2967
rect 3025 2962 3094 2967
rect 673 2957 678 2962
rect 865 2957 870 2962
rect 1089 2957 1222 2962
rect 2697 2957 2806 2962
rect 121 2952 206 2957
rect 337 2952 678 2957
rect 697 2952 870 2957
rect 889 2952 918 2957
rect 1241 2952 1270 2957
rect 1369 2952 1470 2957
rect 1665 2952 2486 2957
rect 2505 2952 2582 2957
rect 2673 2952 2702 2957
rect 2801 2952 2870 2957
rect 2929 2952 3022 2957
rect 3241 2952 3350 2957
rect 1265 2947 1374 2952
rect 3057 2947 3150 2952
rect 257 2942 398 2947
rect 481 2942 590 2947
rect 721 2942 926 2947
rect 945 2942 1094 2947
rect 1113 2942 1182 2947
rect 1393 2942 1574 2947
rect 1697 2942 1774 2947
rect 1801 2942 1910 2947
rect 2001 2942 2166 2947
rect 2233 2942 2302 2947
rect 2553 2942 2638 2947
rect 2713 2942 2822 2947
rect 3033 2942 3062 2947
rect 3145 2942 3286 2947
rect 945 2937 950 2942
rect 161 2932 406 2937
rect 417 2932 534 2937
rect 617 2932 670 2937
rect 833 2932 950 2937
rect 1089 2937 1094 2942
rect 1921 2937 2006 2942
rect 2161 2937 2166 2942
rect 3281 2937 3286 2942
rect 3353 2942 3422 2947
rect 3353 2937 3358 2942
rect 1089 2932 1510 2937
rect 1529 2932 1606 2937
rect 1705 2932 1926 2937
rect 2025 2932 2150 2937
rect 2161 2932 2206 2937
rect 2217 2932 2470 2937
rect 2849 2932 3134 2937
rect 3281 2932 3358 2937
rect 161 2917 166 2932
rect 289 2922 358 2927
rect 137 2912 166 2917
rect 401 2887 406 2932
rect 1505 2927 1510 2932
rect 497 2922 686 2927
rect 761 2922 862 2927
rect 961 2922 1182 2927
rect 1177 2917 1182 2922
rect 1297 2922 1326 2927
rect 1361 2922 1486 2927
rect 1505 2922 1526 2927
rect 1297 2917 1302 2922
rect 1521 2917 1526 2922
rect 1617 2922 2334 2927
rect 2545 2922 2790 2927
rect 2833 2922 2862 2927
rect 2977 2922 3110 2927
rect 3121 2922 3246 2927
rect 1617 2917 1622 2922
rect 2545 2917 2550 2922
rect 2857 2917 2982 2922
rect 3105 2917 3110 2922
rect 545 2912 750 2917
rect 785 2912 838 2917
rect 849 2912 886 2917
rect 905 2912 1006 2917
rect 1017 2912 1150 2917
rect 1177 2912 1302 2917
rect 1329 2912 1446 2917
rect 1465 2912 1494 2917
rect 1521 2912 1622 2917
rect 1729 2912 1782 2917
rect 1793 2912 1950 2917
rect 2017 2912 2094 2917
rect 2177 2912 2550 2917
rect 2561 2912 2590 2917
rect 833 2907 838 2912
rect 505 2902 566 2907
rect 641 2902 806 2907
rect 833 2902 878 2907
rect 1009 2902 1038 2907
rect 1129 2902 1158 2907
rect 1345 2902 1390 2907
rect 1033 2897 1134 2902
rect 1489 2897 1494 2912
rect 1729 2897 1734 2912
rect 2585 2907 2590 2912
rect 2665 2912 2694 2917
rect 3105 2912 3158 2917
rect 2665 2907 2670 2912
rect 1825 2902 1958 2907
rect 1993 2902 2030 2907
rect 2305 2902 2350 2907
rect 2489 2902 2518 2907
rect 2585 2902 2670 2907
rect 2801 2902 2934 2907
rect 3313 2902 3350 2907
rect 689 2892 742 2897
rect 865 2892 990 2897
rect 1489 2892 1734 2897
rect 1889 2892 1918 2897
rect 1913 2887 1918 2892
rect 2041 2892 2390 2897
rect 2041 2887 2046 2892
rect 2385 2887 2390 2892
rect 2465 2892 2494 2897
rect 2465 2887 2470 2892
rect 401 2882 686 2887
rect 681 2877 686 2882
rect 921 2882 950 2887
rect 1001 2882 1030 2887
rect 921 2877 926 2882
rect 681 2872 926 2877
rect 1025 2877 1030 2882
rect 1137 2882 1166 2887
rect 1753 2882 1814 2887
rect 1913 2882 2046 2887
rect 2265 2882 2366 2887
rect 2385 2882 2470 2887
rect 2513 2887 2518 2902
rect 2801 2897 2806 2902
rect 2705 2892 2806 2897
rect 2913 2892 2982 2897
rect 2705 2887 2710 2892
rect 2513 2882 2710 2887
rect 1137 2877 1142 2882
rect 1025 2872 1142 2877
rect 1809 2877 1814 2882
rect 1809 2872 1878 2877
rect 1873 2867 1878 2872
rect 2265 2867 2270 2882
rect 2289 2872 2342 2877
rect 265 2862 390 2867
rect 385 2857 390 2862
rect 529 2862 662 2867
rect 1873 2862 2270 2867
rect 529 2857 534 2862
rect 385 2852 534 2857
rect 553 2842 678 2847
rect 849 2842 918 2847
rect 929 2842 1014 2847
rect 2577 2842 2734 2847
rect 617 2832 670 2837
rect 745 2832 894 2837
rect 2417 2832 2454 2837
rect 2529 2832 2710 2837
rect 361 2822 454 2827
rect 465 2822 494 2827
rect 513 2822 870 2827
rect 1345 2822 1470 2827
rect 1641 2822 1766 2827
rect 2129 2822 2238 2827
rect 2401 2822 2510 2827
rect 2649 2822 2726 2827
rect 2761 2822 2846 2827
rect 2881 2822 2902 2827
rect 2921 2822 3046 2827
rect 1641 2817 1646 2822
rect 593 2812 790 2817
rect 969 2812 1126 2817
rect 1145 2812 1390 2817
rect 1497 2812 1566 2817
rect 1617 2812 1646 2817
rect 1761 2817 1766 2822
rect 2881 2817 2886 2822
rect 1761 2812 2182 2817
rect 2601 2812 2886 2817
rect 3185 2812 3254 2817
rect 969 2807 974 2812
rect 705 2802 846 2807
rect 945 2802 974 2807
rect 1121 2807 1126 2812
rect 1121 2802 1158 2807
rect 2401 2802 2582 2807
rect 1553 2797 1670 2802
rect 585 2792 638 2797
rect 657 2792 742 2797
rect 817 2792 886 2797
rect 1073 2792 1174 2797
rect 1233 2792 1558 2797
rect 1665 2792 1718 2797
rect 1737 2792 1814 2797
rect 1889 2792 1958 2797
rect 2033 2792 2118 2797
rect 2273 2792 2382 2797
rect 1233 2787 1238 2792
rect 1713 2787 1718 2792
rect 2273 2787 2278 2792
rect 425 2782 470 2787
rect 521 2782 630 2787
rect 753 2782 1014 2787
rect 1025 2782 1238 2787
rect 1337 2782 1414 2787
rect 1577 2782 1662 2787
rect 1713 2782 2278 2787
rect 2377 2787 2382 2792
rect 2401 2787 2406 2802
rect 2577 2797 2798 2802
rect 3105 2797 3246 2802
rect 2793 2792 3110 2797
rect 3241 2792 3350 2797
rect 2377 2782 2430 2787
rect 2449 2782 2678 2787
rect 2697 2782 2726 2787
rect 2737 2782 2782 2787
rect 3121 2782 3230 2787
rect 625 2777 758 2782
rect 1009 2777 1014 2782
rect 2449 2777 2454 2782
rect 121 2772 366 2777
rect 417 2772 454 2777
rect 553 2772 606 2777
rect 1009 2772 1110 2777
rect 1249 2772 1318 2777
rect 1105 2767 1254 2772
rect 1313 2767 1318 2772
rect 1433 2772 1590 2777
rect 1433 2767 1438 2772
rect 473 2762 782 2767
rect 1313 2762 1438 2767
rect 1585 2767 1590 2772
rect 1793 2772 1966 2777
rect 2289 2772 2366 2777
rect 2425 2772 2454 2777
rect 2473 2772 2502 2777
rect 2745 2772 2774 2777
rect 2825 2772 2902 2777
rect 2969 2772 3094 2777
rect 1793 2767 1798 2772
rect 1961 2767 2294 2772
rect 2361 2767 2430 2772
rect 2497 2767 2750 2772
rect 2969 2767 2974 2772
rect 1585 2762 1798 2767
rect 1817 2762 1942 2767
rect 2817 2762 2974 2767
rect 3089 2767 3094 2772
rect 3089 2762 3150 2767
rect 985 2757 1086 2762
rect 521 2752 574 2757
rect 865 2752 902 2757
rect 961 2752 990 2757
rect 1081 2752 1110 2757
rect 1225 2752 1294 2757
rect 1513 2752 1566 2757
rect 1849 2752 1926 2757
rect 1937 2752 2686 2757
rect 2705 2752 2750 2757
rect 2985 2752 3078 2757
rect 713 2747 822 2752
rect 1937 2747 1942 2752
rect 2681 2747 2686 2752
rect 2849 2747 2966 2752
rect 489 2742 518 2747
rect 513 2737 518 2742
rect 593 2742 718 2747
rect 817 2742 1134 2747
rect 1457 2742 1502 2747
rect 593 2737 598 2742
rect 1497 2737 1502 2742
rect 1577 2742 1942 2747
rect 1953 2742 1998 2747
rect 2265 2742 2310 2747
rect 2681 2742 2854 2747
rect 2961 2742 3214 2747
rect 1577 2737 1582 2742
rect 2137 2737 2238 2742
rect 2345 2737 2534 2742
rect 513 2732 598 2737
rect 697 2732 806 2737
rect 1497 2732 1582 2737
rect 1809 2732 2142 2737
rect 2233 2732 2254 2737
rect 2329 2732 2350 2737
rect 2529 2732 2758 2737
rect 2865 2732 3086 2737
rect 3169 2732 3366 2737
rect 3385 2732 3438 2737
rect 649 2722 758 2727
rect 777 2722 806 2727
rect 801 2717 806 2722
rect 937 2722 1070 2727
rect 1177 2722 1318 2727
rect 937 2717 942 2722
rect 1177 2717 1182 2722
rect 801 2712 942 2717
rect 1153 2712 1182 2717
rect 1313 2717 1318 2722
rect 1809 2717 1814 2732
rect 2249 2727 2334 2732
rect 2753 2727 2870 2732
rect 1833 2722 1942 2727
rect 2153 2722 2222 2727
rect 2353 2722 2566 2727
rect 2577 2722 2606 2727
rect 2601 2717 2606 2722
rect 2705 2722 2734 2727
rect 2889 2722 2918 2727
rect 2705 2717 2710 2722
rect 2913 2717 2918 2722
rect 3249 2722 3342 2727
rect 3249 2717 3254 2722
rect 1313 2712 1814 2717
rect 2097 2712 2462 2717
rect 2601 2712 2710 2717
rect 2745 2712 2774 2717
rect 2913 2712 3254 2717
rect 3273 2712 3302 2717
rect 2097 2707 2102 2712
rect 1129 2702 1158 2707
rect 1153 2697 1158 2702
rect 1793 2702 1846 2707
rect 1153 2692 1502 2697
rect 1497 2687 1502 2692
rect 1793 2687 1798 2702
rect 1497 2682 1798 2687
rect 1841 2687 1846 2702
rect 1953 2702 2102 2707
rect 2137 2702 2166 2707
rect 2273 2702 2302 2707
rect 1953 2687 1958 2702
rect 2161 2697 2278 2702
rect 2457 2697 2462 2712
rect 2745 2697 2750 2712
rect 3297 2707 3302 2712
rect 3393 2712 3422 2717
rect 3393 2707 3398 2712
rect 3297 2702 3398 2707
rect 2457 2692 2750 2697
rect 2921 2692 2974 2697
rect 1841 2682 1958 2687
rect 2201 2682 2438 2687
rect 2865 2682 2902 2687
rect 3057 2682 3198 2687
rect 841 2672 910 2677
rect 969 2672 1054 2677
rect 1281 2662 1478 2667
rect 1073 2652 1166 2657
rect 1073 2647 1078 2652
rect 721 2642 1078 2647
rect 1161 2647 1166 2652
rect 1281 2647 1286 2662
rect 1161 2642 1286 2647
rect 1473 2647 1478 2662
rect 1969 2662 2182 2667
rect 1785 2652 1854 2657
rect 1785 2647 1790 2652
rect 1473 2642 1790 2647
rect 1849 2647 1854 2652
rect 1969 2647 1974 2662
rect 2177 2657 2182 2662
rect 3393 2662 3438 2667
rect 3393 2657 3398 2662
rect 2177 2652 2406 2657
rect 2441 2652 2550 2657
rect 3193 2652 3262 2657
rect 3345 2652 3398 2657
rect 1849 2642 1974 2647
rect 2401 2647 2406 2652
rect 3193 2647 3198 2652
rect 2401 2642 2430 2647
rect 2641 2642 2886 2647
rect 3145 2642 3198 2647
rect 3257 2647 3262 2652
rect 3257 2642 3334 2647
rect 2241 2637 2318 2642
rect 2641 2637 2646 2642
rect 1297 2632 1462 2637
rect 1985 2632 2246 2637
rect 2313 2632 2646 2637
rect 2881 2637 2886 2642
rect 2881 2632 3158 2637
rect 417 2622 518 2627
rect 529 2622 630 2627
rect 1049 2622 1150 2627
rect 1433 2622 1478 2627
rect 1697 2622 1782 2627
rect 1801 2622 1838 2627
rect 1857 2622 1966 2627
rect 2257 2622 2310 2627
rect 3089 2622 3246 2627
rect 1337 2617 1414 2622
rect 1697 2617 1702 2622
rect 113 2612 326 2617
rect 353 2612 1118 2617
rect 1201 2612 1342 2617
rect 1409 2612 1702 2617
rect 1777 2617 1782 2622
rect 1857 2617 1862 2622
rect 1777 2612 1862 2617
rect 1961 2617 1966 2622
rect 1961 2612 2150 2617
rect 2393 2612 2470 2617
rect 2529 2612 2958 2617
rect 3081 2612 3342 2617
rect 2145 2607 2150 2612
rect 121 2602 342 2607
rect 1353 2602 1446 2607
rect 1457 2602 1486 2607
rect 1713 2602 1774 2607
rect 1825 2602 1998 2607
rect 2145 2602 2238 2607
rect 2385 2602 2462 2607
rect 2873 2602 3038 2607
rect 3201 2602 3414 2607
rect 361 2597 518 2602
rect 1073 2597 1198 2602
rect 2017 2597 2110 2602
rect 2233 2597 2238 2602
rect 2481 2597 2830 2602
rect 97 2592 214 2597
rect 321 2592 366 2597
rect 513 2592 542 2597
rect 897 2592 1078 2597
rect 1193 2592 1430 2597
rect 1449 2592 1670 2597
rect 1993 2592 2022 2597
rect 2105 2592 2134 2597
rect 2233 2592 2486 2597
rect 2825 2592 2854 2597
rect 3033 2592 3206 2597
rect 3225 2592 3366 2597
rect 209 2587 214 2592
rect 1425 2587 1430 2592
rect 2873 2587 3006 2592
rect 3201 2587 3206 2592
rect 209 2582 494 2587
rect 489 2577 494 2582
rect 553 2582 942 2587
rect 1089 2582 1214 2587
rect 1425 2582 2158 2587
rect 2265 2582 2350 2587
rect 2433 2582 2878 2587
rect 3001 2582 3030 2587
rect 553 2577 558 2582
rect 937 2577 1094 2582
rect 1233 2577 1326 2582
rect 3025 2577 3030 2582
rect 3161 2582 3190 2587
rect 3201 2582 3286 2587
rect 3161 2577 3166 2582
rect 345 2572 470 2577
rect 489 2572 558 2577
rect 1113 2572 1238 2577
rect 1321 2572 1414 2577
rect 1641 2572 3006 2577
rect 3025 2572 3166 2577
rect 1409 2567 1646 2572
rect 889 2562 958 2567
rect 393 2557 486 2562
rect 889 2557 894 2562
rect 305 2552 398 2557
rect 481 2552 726 2557
rect 865 2552 894 2557
rect 953 2557 958 2562
rect 1001 2562 1094 2567
rect 1241 2562 1310 2567
rect 1665 2562 1846 2567
rect 1913 2562 2086 2567
rect 2121 2562 2446 2567
rect 2481 2562 2510 2567
rect 2745 2562 2854 2567
rect 2881 2562 2950 2567
rect 3377 2562 3438 2567
rect 1001 2557 1006 2562
rect 953 2552 1006 2557
rect 1089 2557 1094 2562
rect 2505 2557 2750 2562
rect 1089 2552 2054 2557
rect 2049 2547 2158 2552
rect 2265 2547 2414 2552
rect 353 2542 550 2547
rect 545 2537 550 2542
rect 617 2542 742 2547
rect 857 2542 990 2547
rect 1017 2542 1086 2547
rect 1249 2542 1990 2547
rect 2153 2542 2270 2547
rect 2409 2542 2438 2547
rect 2497 2542 2758 2547
rect 3065 2542 3166 2547
rect 617 2537 622 2542
rect 545 2532 622 2537
rect 737 2527 742 2542
rect 1137 2537 1230 2542
rect 2497 2537 2502 2542
rect 889 2532 1142 2537
rect 1225 2532 1294 2537
rect 1385 2532 1542 2537
rect 1817 2532 2502 2537
rect 1289 2527 1390 2532
rect 1537 2527 1822 2532
rect 737 2522 926 2527
rect 1033 2522 1270 2527
rect 1409 2522 1518 2527
rect 1841 2522 1998 2527
rect 2089 2522 2166 2527
rect 2241 2522 2286 2527
rect 2473 2522 2606 2527
rect 3321 2522 3350 2527
rect 921 2517 926 2522
rect 2241 2517 2246 2522
rect 81 2512 182 2517
rect 465 2512 518 2517
rect 921 2512 1014 2517
rect 1161 2512 1318 2517
rect 1545 2512 1622 2517
rect 1721 2512 1926 2517
rect 1969 2512 2246 2517
rect 2289 2512 2630 2517
rect 2665 2512 2758 2517
rect 1009 2507 1014 2512
rect 1545 2507 1550 2512
rect 1009 2502 1078 2507
rect 1137 2502 1190 2507
rect 1265 2502 1550 2507
rect 1617 2507 1622 2512
rect 1617 2502 1758 2507
rect 1833 2502 1862 2507
rect 2097 2502 2198 2507
rect 2217 2502 2262 2507
rect 2401 2502 2478 2507
rect 2489 2502 2614 2507
rect 3033 2502 3102 2507
rect 1073 2497 1078 2502
rect 2097 2497 2102 2502
rect 2193 2497 2198 2502
rect 2401 2497 2406 2502
rect 625 2492 766 2497
rect 953 2492 1062 2497
rect 1073 2492 1254 2497
rect 1561 2492 1606 2497
rect 1769 2492 2102 2497
rect 2113 2492 2158 2497
rect 2193 2492 2406 2497
rect 2425 2492 2454 2497
rect 1249 2487 1566 2492
rect 1601 2487 1774 2492
rect 2449 2487 2454 2492
rect 2769 2492 2838 2497
rect 3289 2492 3430 2497
rect 2769 2487 2774 2492
rect 865 2482 950 2487
rect 2449 2482 2774 2487
rect 1105 2477 1206 2482
rect 377 2472 614 2477
rect 609 2467 614 2472
rect 689 2472 862 2477
rect 689 2467 694 2472
rect 609 2462 694 2467
rect 857 2467 862 2472
rect 1081 2472 1110 2477
rect 1201 2472 1230 2477
rect 1081 2467 1086 2472
rect 1225 2467 1230 2472
rect 1313 2472 1710 2477
rect 1921 2472 2014 2477
rect 2825 2472 3046 2477
rect 3425 2472 3430 2492
rect 1313 2467 1318 2472
rect 857 2462 1086 2467
rect 1105 2462 1206 2467
rect 1225 2462 1318 2467
rect 1729 2462 1902 2467
rect 1729 2457 1734 2462
rect 713 2452 838 2457
rect 1545 2452 1734 2457
rect 1897 2457 1902 2462
rect 2081 2462 2430 2467
rect 1897 2452 2014 2457
rect 2033 2452 2062 2457
rect 1545 2447 1550 2452
rect 2009 2447 2014 2452
rect 2081 2447 2086 2462
rect 2425 2447 2430 2462
rect 2593 2452 2654 2457
rect 1337 2442 1550 2447
rect 1753 2442 1878 2447
rect 2009 2442 2086 2447
rect 2105 2442 2406 2447
rect 2425 2442 2454 2447
rect 2473 2442 2574 2447
rect 2841 2442 2998 2447
rect 1753 2437 1758 2442
rect 241 2432 342 2437
rect 385 2432 430 2437
rect 609 2432 726 2437
rect 1561 2432 1758 2437
rect 1873 2437 1878 2442
rect 2105 2437 2110 2442
rect 1873 2432 2110 2437
rect 2401 2437 2406 2442
rect 2473 2437 2478 2442
rect 2569 2437 2694 2442
rect 2401 2432 2478 2437
rect 2689 2432 2718 2437
rect 2737 2432 2846 2437
rect 2953 2432 3238 2437
rect 3313 2432 3406 2437
rect 2129 2427 2382 2432
rect 449 2422 590 2427
rect 369 2417 454 2422
rect 585 2417 590 2422
rect 745 2422 1102 2427
rect 1145 2422 1246 2427
rect 1465 2422 1606 2427
rect 1753 2422 2134 2427
rect 2377 2422 2998 2427
rect 745 2417 750 2422
rect 345 2412 374 2417
rect 585 2412 750 2417
rect 1097 2417 1102 2422
rect 1097 2412 1126 2417
rect 1289 2412 1766 2417
rect 1777 2412 2974 2417
rect 913 2407 1054 2412
rect 2993 2407 2998 2422
rect 361 2402 414 2407
rect 777 2402 846 2407
rect 777 2397 782 2402
rect 313 2392 782 2397
rect 841 2397 846 2402
rect 889 2402 918 2407
rect 1049 2402 1078 2407
rect 889 2397 894 2402
rect 841 2392 894 2397
rect 1073 2397 1078 2402
rect 1185 2402 1702 2407
rect 1745 2402 1782 2407
rect 2137 2402 2702 2407
rect 2993 2402 3094 2407
rect 1185 2397 1190 2402
rect 1697 2397 1702 2402
rect 1777 2397 2142 2402
rect 1073 2392 1190 2397
rect 1209 2392 1366 2397
rect 1401 2392 1534 2397
rect 1577 2392 1686 2397
rect 1697 2392 1758 2397
rect 2161 2392 2342 2397
rect 2337 2387 2342 2392
rect 2425 2392 2606 2397
rect 2721 2392 2750 2397
rect 2425 2387 2430 2392
rect 2601 2387 2726 2392
rect 225 2382 294 2387
rect 721 2382 1054 2387
rect 1257 2382 1438 2387
rect 225 2377 230 2382
rect 89 2372 230 2377
rect 289 2377 294 2382
rect 1049 2377 1262 2382
rect 1433 2377 1438 2382
rect 1553 2382 1582 2387
rect 1689 2382 1814 2387
rect 1825 2382 1878 2387
rect 1897 2382 2134 2387
rect 2145 2382 2318 2387
rect 2337 2382 2430 2387
rect 3161 2382 3302 2387
rect 1553 2377 1558 2382
rect 1897 2377 1902 2382
rect 2129 2377 2134 2382
rect 2473 2377 2582 2382
rect 289 2372 1030 2377
rect 1433 2372 1558 2377
rect 1617 2372 1662 2377
rect 1281 2367 1390 2372
rect 1657 2367 1662 2372
rect 1873 2372 1902 2377
rect 2025 2372 2070 2377
rect 2129 2372 2294 2377
rect 2449 2372 2478 2377
rect 2577 2372 3110 2377
rect 1873 2367 1878 2372
rect 73 2362 102 2367
rect 809 2362 982 2367
rect 1081 2362 1286 2367
rect 1385 2362 1414 2367
rect 1657 2362 1878 2367
rect 1897 2362 1990 2367
rect 2081 2362 2734 2367
rect 97 2347 102 2362
rect 217 2357 582 2362
rect 689 2357 814 2362
rect 1985 2357 2086 2362
rect 217 2347 222 2357
rect 577 2352 694 2357
rect 833 2352 1038 2357
rect 1297 2352 1366 2357
rect 1497 2352 1598 2357
rect 2225 2352 2262 2357
rect 2465 2352 2542 2357
rect 2649 2352 2806 2357
rect 2817 2352 2862 2357
rect 1297 2347 1302 2352
rect 1385 2347 1470 2352
rect 2105 2347 2206 2352
rect 2353 2347 2470 2352
rect 2537 2347 2654 2352
rect 2801 2347 2806 2352
rect 97 2342 222 2347
rect 241 2342 294 2347
rect 321 2342 558 2347
rect 713 2342 870 2347
rect 881 2342 1070 2347
rect 1089 2342 1166 2347
rect 1257 2342 1302 2347
rect 1345 2342 1390 2347
rect 1465 2342 1638 2347
rect 1769 2342 2110 2347
rect 2201 2342 2358 2347
rect 2481 2342 2518 2347
rect 2801 2342 2870 2347
rect 881 2337 886 2342
rect 513 2332 606 2337
rect 761 2332 886 2337
rect 1041 2337 1046 2342
rect 2481 2337 2486 2342
rect 1041 2332 1454 2337
rect 1609 2332 1726 2337
rect 2121 2332 2486 2337
rect 2537 2332 2782 2337
rect 761 2327 766 2332
rect 945 2327 1022 2332
rect 1449 2327 1614 2332
rect 1953 2327 2102 2332
rect 2537 2327 2542 2332
rect 2777 2327 2918 2332
rect 257 2322 766 2327
rect 777 2322 950 2327
rect 1017 2322 1110 2327
rect 1153 2322 1294 2327
rect 1377 2322 1430 2327
rect 1753 2322 1958 2327
rect 2097 2322 2542 2327
rect 2913 2322 2942 2327
rect 3041 2322 3078 2327
rect 3385 2322 3430 2327
rect 1289 2317 1382 2322
rect 1425 2317 1430 2322
rect 529 2312 822 2317
rect 961 2312 1014 2317
rect 1425 2312 1638 2317
rect 1713 2312 1790 2317
rect 1969 2312 3174 2317
rect 3361 2312 3398 2317
rect 1097 2307 1270 2312
rect 1633 2307 1638 2312
rect 1785 2307 1974 2312
rect 273 2302 366 2307
rect 537 2302 814 2307
rect 841 2302 934 2307
rect 953 2302 1102 2307
rect 1265 2302 1294 2307
rect 1313 2302 1390 2307
rect 1633 2302 1766 2307
rect 1993 2302 2598 2307
rect 2761 2302 2958 2307
rect 841 2297 846 2302
rect 465 2292 566 2297
rect 617 2292 846 2297
rect 929 2297 934 2302
rect 1313 2297 1318 2302
rect 929 2292 966 2297
rect 1113 2292 1318 2297
rect 1385 2297 1390 2302
rect 2593 2297 2766 2302
rect 2953 2297 2958 2302
rect 3033 2302 3078 2307
rect 3033 2297 3038 2302
rect 1385 2292 1902 2297
rect 2033 2292 2134 2297
rect 2225 2292 2390 2297
rect 2953 2292 3038 2297
rect 985 2287 1094 2292
rect 673 2282 702 2287
rect 697 2277 702 2282
rect 785 2282 990 2287
rect 1089 2282 1374 2287
rect 2001 2282 2054 2287
rect 2137 2282 2822 2287
rect 785 2277 790 2282
rect 1641 2277 1982 2282
rect 2817 2277 2822 2282
rect 3057 2282 3086 2287
rect 3057 2277 3062 2282
rect 697 2272 790 2277
rect 809 2272 1102 2277
rect 1121 2272 1526 2277
rect 1617 2272 1646 2277
rect 1977 2272 2166 2277
rect 2177 2272 2278 2277
rect 2753 2272 2798 2277
rect 2817 2272 3062 2277
rect 833 2262 1214 2267
rect 1337 2262 1398 2267
rect 1209 2257 1342 2262
rect 1417 2257 1566 2262
rect 1617 2257 1622 2272
rect 2297 2267 2478 2272
rect 1641 2262 2302 2267
rect 2473 2262 2502 2267
rect 577 2252 678 2257
rect 705 2252 790 2257
rect 841 2252 1190 2257
rect 1361 2252 1422 2257
rect 1561 2252 1622 2257
rect 1689 2252 1814 2257
rect 1897 2252 1998 2257
rect 2081 2252 2534 2257
rect 2569 2252 2646 2257
rect 497 2242 686 2247
rect 705 2237 710 2252
rect 785 2247 790 2252
rect 2569 2247 2574 2252
rect 785 2242 1118 2247
rect 1145 2242 1270 2247
rect 1297 2242 1422 2247
rect 1449 2242 1550 2247
rect 1809 2242 2070 2247
rect 2241 2242 2302 2247
rect 2345 2242 2406 2247
rect 2449 2242 2574 2247
rect 2641 2247 2646 2252
rect 2641 2242 2982 2247
rect 1265 2237 1270 2242
rect 2089 2237 2222 2242
rect 417 2232 486 2237
rect 569 2232 710 2237
rect 785 2232 982 2237
rect 1065 2232 1166 2237
rect 1265 2232 1302 2237
rect 1385 2232 1654 2237
rect 1673 2232 1782 2237
rect 1833 2232 2094 2237
rect 2217 2232 2246 2237
rect 2353 2232 2478 2237
rect 3057 2232 3118 2237
rect 481 2227 574 2232
rect 1777 2227 1782 2232
rect 2689 2227 2790 2232
rect 393 2222 430 2227
rect 593 2222 814 2227
rect 929 2222 998 2227
rect 1137 2222 1230 2227
rect 1313 2222 1558 2227
rect 1585 2222 1638 2227
rect 1657 2222 1766 2227
rect 1777 2222 2182 2227
rect 2233 2222 2366 2227
rect 2585 2222 2694 2227
rect 2785 2222 2814 2227
rect 2905 2222 3046 2227
rect 3129 2222 3206 2227
rect 1017 2217 1118 2222
rect 1249 2217 1318 2222
rect 257 2197 262 2217
rect 321 2212 422 2217
rect 521 2212 806 2217
rect 825 2212 1022 2217
rect 1113 2212 1254 2217
rect 1377 2212 1398 2217
rect 1433 2212 2494 2217
rect 2569 2212 2622 2217
rect 2705 2212 2854 2217
rect 2977 2212 3286 2217
rect 801 2207 806 2212
rect 1393 2207 1398 2212
rect 2873 2207 2982 2212
rect 481 2202 758 2207
rect 801 2202 982 2207
rect 993 2202 1158 2207
rect 1185 2202 1246 2207
rect 1297 2202 1366 2207
rect 1393 2202 1430 2207
rect 1441 2202 1494 2207
rect 81 2192 262 2197
rect 513 2192 686 2197
rect 705 2192 838 2197
rect 913 2192 942 2197
rect 833 2187 838 2192
rect 977 2187 982 2202
rect 1185 2197 1190 2202
rect 1505 2197 1510 2207
rect 1681 2202 1774 2207
rect 1849 2202 1894 2207
rect 1929 2202 1990 2207
rect 2049 2202 2118 2207
rect 2177 2202 2598 2207
rect 2689 2202 2878 2207
rect 2993 2202 3142 2207
rect 3281 2202 3286 2212
rect 3313 2202 3398 2207
rect 1017 2192 1070 2197
rect 1081 2192 1190 2197
rect 1201 2192 1278 2197
rect 1289 2192 1622 2197
rect 1737 2192 1766 2197
rect 1897 2192 1934 2197
rect 1969 2192 2030 2197
rect 2161 2192 2310 2197
rect 2481 2192 2742 2197
rect 2865 2192 3006 2197
rect 3041 2192 3078 2197
rect 1201 2187 1206 2192
rect 1785 2187 1878 2192
rect 2361 2187 2462 2192
rect 89 2182 118 2187
rect 273 2182 614 2187
rect 641 2182 718 2187
rect 785 2182 822 2187
rect 833 2182 966 2187
rect 977 2182 1206 2187
rect 1217 2182 1238 2187
rect 1377 2182 1454 2187
rect 1465 2182 1542 2187
rect 113 2177 278 2182
rect 641 2177 646 2182
rect 785 2177 790 2182
rect 1425 2177 1430 2182
rect 1537 2177 1542 2182
rect 1601 2182 1630 2187
rect 1729 2182 1790 2187
rect 1873 2182 1942 2187
rect 1953 2182 2150 2187
rect 2177 2182 2262 2187
rect 2337 2182 2366 2187
rect 2457 2182 2654 2187
rect 2809 2182 2870 2187
rect 2913 2182 3070 2187
rect 3337 2182 3382 2187
rect 1601 2177 1606 2182
rect 1953 2177 1958 2182
rect 521 2172 646 2177
rect 657 2172 790 2177
rect 849 2172 982 2177
rect 1001 2172 1030 2177
rect 1121 2172 1150 2177
rect 1161 2172 1398 2177
rect 1425 2172 1518 2177
rect 1537 2172 1606 2177
rect 1721 2172 1806 2177
rect 1825 2172 1958 2177
rect 2041 2172 2566 2177
rect 2673 2172 2774 2177
rect 2801 2172 2910 2177
rect 3025 2172 3110 2177
rect 3129 2172 3214 2177
rect 185 2162 262 2167
rect 281 2162 606 2167
rect 649 2162 806 2167
rect 281 2157 286 2162
rect 849 2157 854 2172
rect 1393 2167 1398 2172
rect 2673 2167 2678 2172
rect 865 2162 1262 2167
rect 1393 2162 1438 2167
rect 1745 2162 1910 2167
rect 2017 2162 2246 2167
rect 2289 2162 2678 2167
rect 2769 2167 2774 2172
rect 3129 2167 3134 2172
rect 2769 2162 3134 2167
rect 3209 2167 3214 2172
rect 3209 2162 3238 2167
rect 1457 2157 1550 2162
rect 233 2152 286 2157
rect 417 2152 550 2157
rect 609 2152 702 2157
rect 737 2152 854 2157
rect 937 2152 1078 2157
rect 1129 2152 1158 2157
rect 1169 2152 1366 2157
rect 1401 2152 1462 2157
rect 1545 2152 1574 2157
rect 1633 2152 1694 2157
rect 1721 2152 2454 2157
rect 2641 2152 2766 2157
rect 2785 2152 3246 2157
rect 3337 2152 3366 2157
rect 609 2147 614 2152
rect 2473 2147 2574 2152
rect 2785 2147 2790 2152
rect 193 2142 614 2147
rect 625 2142 670 2147
rect 793 2142 1118 2147
rect 1153 2142 1294 2147
rect 1305 2142 1534 2147
rect 1553 2142 1590 2147
rect 1625 2142 1774 2147
rect 1873 2142 1902 2147
rect 2009 2142 2478 2147
rect 2569 2142 2598 2147
rect 2609 2142 2790 2147
rect 2809 2142 2878 2147
rect 2889 2142 2982 2147
rect 3065 2142 3166 2147
rect 3177 2142 3254 2147
rect 3265 2142 3350 2147
rect 3361 2142 3366 2152
rect 1553 2137 1558 2142
rect 3249 2137 3254 2142
rect 137 2132 1558 2137
rect 1697 2132 1846 2137
rect 1857 2132 1990 2137
rect 2153 2132 2214 2137
rect 1473 2127 1478 2132
rect 2057 2127 2134 2132
rect 2225 2127 2230 2137
rect 2281 2132 2334 2137
rect 2369 2132 3198 2137
rect 3249 2132 3334 2137
rect 3345 2132 3350 2142
rect 3361 2132 3398 2137
rect 249 2122 318 2127
rect 369 2117 374 2127
rect 385 2122 550 2127
rect 641 2122 694 2127
rect 833 2117 838 2127
rect 849 2122 934 2127
rect 1025 2122 1046 2127
rect 1057 2122 1438 2127
rect 1473 2122 1494 2127
rect 1569 2122 1654 2127
rect 1777 2122 1798 2127
rect 1865 2122 2062 2127
rect 2129 2122 2286 2127
rect 2337 2122 2430 2127
rect 2513 2122 2550 2127
rect 2705 2122 2742 2127
rect 2841 2122 3126 2127
rect 3177 2122 3270 2127
rect 3321 2122 3414 2127
rect 2569 2117 2686 2122
rect 3121 2117 3126 2122
rect 97 2112 254 2117
rect 369 2112 678 2117
rect 721 2112 766 2117
rect 833 2112 1046 2117
rect 1129 2112 1166 2117
rect 1193 2112 1238 2117
rect 1337 2112 1614 2117
rect 1761 2112 1798 2117
rect 1921 2112 1966 2117
rect 2073 2112 2118 2117
rect 2129 2112 2574 2117
rect 2681 2112 2990 2117
rect 3041 2112 3102 2117
rect 3121 2112 3166 2117
rect 3185 2112 3222 2117
rect 3305 2112 3406 2117
rect 2129 2107 2134 2112
rect 225 2102 542 2107
rect 641 2102 686 2107
rect 809 2102 1678 2107
rect 1745 2102 1830 2107
rect 1873 2102 2078 2107
rect 2105 2102 2134 2107
rect 2177 2102 2414 2107
rect 2449 2102 2478 2107
rect 2553 2102 2958 2107
rect 3041 2102 3062 2107
rect 3081 2102 3102 2107
rect 3233 2102 3286 2107
rect 169 2092 726 2097
rect 745 2092 894 2097
rect 905 2092 942 2097
rect 1025 2092 1158 2097
rect 1217 2092 2014 2097
rect 2225 2092 2270 2097
rect 2281 2092 2446 2097
rect 2489 2092 2518 2097
rect 2545 2092 3110 2097
rect 3145 2092 3398 2097
rect 2033 2087 2174 2092
rect 2513 2087 2518 2092
rect 89 2082 238 2087
rect 409 2082 574 2087
rect 601 2082 710 2087
rect 785 2082 854 2087
rect 905 2082 1350 2087
rect 1433 2082 1542 2087
rect 1793 2082 1934 2087
rect 1953 2082 2038 2087
rect 2169 2082 2198 2087
rect 2233 2082 2502 2087
rect 2513 2082 2622 2087
rect 2689 2082 3078 2087
rect 3329 2082 3358 2087
rect 785 2077 790 2082
rect 1561 2077 1678 2082
rect 3073 2077 3270 2082
rect 3329 2077 3334 2082
rect 265 2072 654 2077
rect 721 2072 790 2077
rect 801 2072 1150 2077
rect 1185 2072 1374 2077
rect 1513 2072 1566 2077
rect 1673 2072 1702 2077
rect 1713 2072 1790 2077
rect 1809 2072 1902 2077
rect 2009 2072 2142 2077
rect 2185 2072 2494 2077
rect 2505 2072 2942 2077
rect 3001 2072 3054 2077
rect 3265 2072 3334 2077
rect 649 2067 726 2072
rect 1697 2067 1702 2072
rect 369 2062 502 2067
rect 777 2062 1686 2067
rect 1697 2062 2046 2067
rect 2073 2062 2246 2067
rect 2553 2062 2742 2067
rect 3017 2062 3062 2067
rect 3121 2062 3246 2067
rect 529 2057 614 2062
rect 2241 2057 2558 2062
rect 377 2052 534 2057
rect 609 2052 710 2057
rect 825 2052 1286 2057
rect 1281 2047 1286 2052
rect 1369 2052 1406 2057
rect 1521 2052 1750 2057
rect 1761 2052 2086 2057
rect 2153 2052 2222 2057
rect 2577 2052 2670 2057
rect 2721 2052 2814 2057
rect 2977 2052 3022 2057
rect 1369 2047 1374 2052
rect 105 2042 214 2047
rect 225 2042 294 2047
rect 337 2042 598 2047
rect 681 2042 974 2047
rect 1001 2042 1078 2047
rect 1089 2042 1118 2047
rect 1137 2042 1166 2047
rect 1177 2042 1262 2047
rect 1281 2042 1374 2047
rect 1665 2042 2142 2047
rect 2233 2042 2590 2047
rect 2641 2042 2686 2047
rect 2753 2042 2806 2047
rect 3073 2042 3174 2047
rect 2137 2037 2238 2042
rect 2929 2037 3030 2042
rect 3073 2037 3078 2042
rect 121 2032 238 2037
rect 409 2032 454 2037
rect 473 2032 526 2037
rect 545 2032 654 2037
rect 809 2032 926 2037
rect 945 2032 1238 2037
rect 1393 2032 1566 2037
rect 1713 2032 1806 2037
rect 1817 2032 1846 2037
rect 1865 2032 1894 2037
rect 1993 2032 2046 2037
rect 2065 2032 2094 2037
rect 2257 2032 2286 2037
rect 2393 2032 2454 2037
rect 2617 2032 2934 2037
rect 3025 2032 3078 2037
rect 3169 2037 3174 2042
rect 3169 2032 3254 2037
rect 673 2027 790 2032
rect 945 2027 950 2032
rect 1841 2027 1846 2032
rect 1889 2027 1998 2032
rect 209 2022 678 2027
rect 785 2022 950 2027
rect 977 2022 1198 2027
rect 1217 2022 1270 2027
rect 1441 2022 1478 2027
rect 1649 2022 1750 2027
rect 1769 2022 1830 2027
rect 1841 2022 1862 2027
rect 2017 2022 2158 2027
rect 2177 2022 2254 2027
rect 2273 2022 2398 2027
rect 2593 2022 2678 2027
rect 2697 2022 3214 2027
rect 3257 2022 3294 2027
rect 169 2012 302 2017
rect 465 2012 574 2017
rect 657 2012 774 2017
rect 801 2012 870 2017
rect 961 2012 1006 2017
rect 1081 2012 1294 2017
rect 1361 2012 1462 2017
rect 1569 2012 1822 2017
rect 1937 2012 2014 2017
rect 2025 2012 2062 2017
rect 2081 2012 2246 2017
rect 2257 2012 2342 2017
rect 2377 2012 2518 2017
rect 2561 2012 2662 2017
rect 769 2007 774 2012
rect 2673 2007 2678 2022
rect 2713 2012 2894 2017
rect 2953 2012 3094 2017
rect 3089 2007 3190 2012
rect 121 2002 206 2007
rect 249 2002 406 2007
rect 417 2002 742 2007
rect 769 2002 1350 2007
rect 1449 2002 1726 2007
rect 1745 2002 2654 2007
rect 2673 2002 2830 2007
rect 2985 2002 3054 2007
rect 3185 2002 3270 2007
rect 417 1997 422 2002
rect 1345 1997 1454 2002
rect 105 1992 158 1997
rect 289 1992 422 1997
rect 465 1992 574 1997
rect 721 1992 1318 1997
rect 1473 1992 1518 1997
rect 1633 1992 2310 1997
rect 2329 1992 2454 1997
rect 2529 1992 2694 1997
rect 2993 1992 3238 1997
rect 2449 1987 2454 1992
rect 65 1982 158 1987
rect 329 1982 534 1987
rect 593 1982 822 1987
rect 841 1982 918 1987
rect 929 1982 1006 1987
rect 1033 1982 1054 1987
rect 1065 1982 1182 1987
rect 1217 1982 1262 1987
rect 1409 1982 1614 1987
rect 1729 1982 2022 1987
rect 2033 1982 2070 1987
rect 2129 1982 2278 1987
rect 2337 1982 2358 1987
rect 2393 1982 2430 1987
rect 2449 1982 2558 1987
rect 2609 1982 2822 1987
rect 2833 1982 2870 1987
rect 3001 1982 3054 1987
rect 913 1977 918 1982
rect 289 1972 398 1977
rect 409 1972 486 1977
rect 553 1972 894 1977
rect 913 1972 1054 1977
rect 1193 1972 1366 1977
rect 1073 1967 1174 1972
rect 217 1962 278 1967
rect 465 1962 486 1967
rect 585 1962 630 1967
rect 713 1962 918 1967
rect 937 1962 1078 1967
rect 1169 1962 1294 1967
rect 1409 1962 1414 1982
rect 2817 1977 2822 1982
rect 1441 1972 1526 1977
rect 1569 1972 1774 1977
rect 1873 1972 1942 1977
rect 1953 1972 1982 1977
rect 2001 1972 2030 1977
rect 2041 1972 2646 1977
rect 2665 1972 2726 1977
rect 2817 1972 3310 1977
rect 2641 1967 2646 1972
rect 1449 1962 1670 1967
rect 1785 1962 2470 1967
rect 2505 1962 2590 1967
rect 2641 1962 2910 1967
rect 3017 1962 3062 1967
rect 3153 1962 3182 1967
rect 505 1957 590 1962
rect 153 1952 510 1957
rect 601 1952 806 1957
rect 833 1952 902 1957
rect 913 1947 918 1962
rect 1313 1957 1414 1962
rect 961 1952 1102 1957
rect 1145 1952 1318 1957
rect 1425 1952 1502 1957
rect 1681 1952 2598 1957
rect 2801 1952 2830 1957
rect 3001 1952 3262 1957
rect 1521 1947 1646 1952
rect 2617 1947 2726 1952
rect 209 1942 270 1947
rect 409 1942 462 1947
rect 513 1942 574 1947
rect 777 1942 846 1947
rect 857 1942 878 1947
rect 913 1942 1030 1947
rect 1185 1942 1262 1947
rect 1313 1942 1526 1947
rect 1641 1942 1902 1947
rect 1937 1942 2366 1947
rect 2441 1942 2622 1947
rect 2721 1942 2966 1947
rect 3033 1942 3062 1947
rect 321 1937 414 1942
rect 1049 1937 1166 1942
rect 273 1932 326 1937
rect 433 1932 670 1937
rect 801 1932 1054 1937
rect 1161 1932 1542 1937
rect 1561 1932 1630 1937
rect 689 1927 782 1932
rect 1713 1927 1822 1932
rect 1937 1927 1942 1942
rect 3057 1937 3062 1942
rect 3145 1942 3174 1947
rect 3145 1937 3150 1942
rect 97 1922 342 1927
rect 377 1922 526 1927
rect 561 1922 694 1927
rect 777 1922 862 1927
rect 913 1922 942 1927
rect 977 1922 1094 1927
rect 1129 1922 1158 1927
rect 1233 1922 1558 1927
rect 1585 1922 1718 1927
rect 1817 1922 1942 1927
rect 1985 1932 2710 1937
rect 3057 1932 3150 1937
rect 3177 1932 3214 1937
rect 1985 1922 1990 1932
rect 1996 1922 2094 1927
rect 2177 1922 2334 1927
rect 2353 1922 2470 1927
rect 2561 1922 2670 1927
rect 2801 1922 2918 1927
rect 2937 1922 2990 1927
rect 449 1912 542 1917
rect 577 1912 854 1917
rect 881 1912 1190 1917
rect 1321 1912 1350 1917
rect 1417 1912 1518 1917
rect 1529 1912 1550 1917
rect 1585 1912 1590 1922
rect 1996 1917 2001 1922
rect 1729 1912 2001 1917
rect 2009 1912 2118 1917
rect 2137 1912 2550 1917
rect 2649 1912 2702 1917
rect 3033 1912 3110 1917
rect 3185 1912 3230 1917
rect 849 1907 854 1912
rect 2113 1907 2118 1912
rect 3281 1907 3286 1937
rect 3425 1922 3504 1927
rect 3297 1912 3406 1917
rect 185 1902 262 1907
rect 273 1902 310 1907
rect 361 1902 662 1907
rect 681 1902 758 1907
rect 849 1902 990 1907
rect 1065 1902 1238 1907
rect 1281 1902 1326 1907
rect 1377 1902 1430 1907
rect 1617 1902 1654 1907
rect 1809 1902 1854 1907
rect 1873 1902 2102 1907
rect 2113 1902 2174 1907
rect 2233 1902 2278 1907
rect 2289 1902 2350 1907
rect 2393 1902 2438 1907
rect 2561 1902 2638 1907
rect 1281 1897 1286 1902
rect 1873 1897 1878 1902
rect 2633 1897 2638 1902
rect 2713 1902 2830 1907
rect 3281 1902 3318 1907
rect 3353 1902 3414 1907
rect 2713 1897 2718 1902
rect 489 1892 542 1897
rect 553 1892 726 1897
rect 745 1892 1102 1897
rect 1217 1892 1286 1897
rect 1305 1892 1342 1897
rect 1425 1892 1494 1897
rect 1521 1892 1542 1897
rect 1585 1892 1742 1897
rect 1833 1892 1878 1897
rect 1897 1892 2038 1897
rect 2065 1892 2182 1897
rect 2249 1892 2390 1897
rect 2425 1892 2454 1897
rect 2513 1892 2614 1897
rect 2633 1892 2718 1897
rect 1217 1887 1222 1892
rect 3313 1887 3318 1902
rect 3345 1892 3382 1897
rect 377 1882 462 1887
rect 481 1882 670 1887
rect 785 1882 926 1887
rect 961 1882 1070 1887
rect 1081 1882 1150 1887
rect 1161 1882 1222 1887
rect 1257 1882 1670 1887
rect 1793 1882 2014 1887
rect 2025 1882 2054 1887
rect 2065 1882 2126 1887
rect 2169 1882 2310 1887
rect 2377 1882 2462 1887
rect 2569 1882 2598 1887
rect 3313 1882 3350 1887
rect 3377 1882 3382 1892
rect 377 1877 382 1882
rect 97 1872 174 1877
rect 353 1872 382 1877
rect 457 1877 462 1882
rect 1689 1877 1798 1882
rect 2049 1877 2054 1882
rect 457 1872 582 1877
rect 601 1872 942 1877
rect 1025 1872 1358 1877
rect 1369 1872 1422 1877
rect 1497 1872 1694 1877
rect 1817 1872 1862 1877
rect 1905 1872 2014 1877
rect 2049 1872 2446 1877
rect 2577 1872 2614 1877
rect 97 1837 102 1872
rect 281 1862 870 1867
rect 897 1862 1398 1867
rect 1545 1862 1606 1867
rect 1697 1862 1758 1867
rect 1817 1862 1870 1867
rect 1953 1862 2102 1867
rect 2185 1862 2222 1867
rect 2281 1862 2358 1867
rect 2401 1862 2630 1867
rect 2729 1862 2766 1867
rect 2785 1862 2878 1867
rect 2785 1857 2790 1862
rect 129 1852 166 1857
rect 561 1852 790 1857
rect 817 1852 934 1857
rect 945 1852 982 1857
rect 1041 1852 1142 1857
rect 1153 1852 1206 1857
rect 1297 1852 1526 1857
rect 1705 1852 2246 1857
rect 2345 1852 2422 1857
rect 2441 1852 2470 1857
rect 2481 1852 2790 1857
rect 2873 1857 2878 1862
rect 2921 1862 3022 1867
rect 2921 1857 2926 1862
rect 2873 1852 2926 1857
rect 3017 1857 3022 1862
rect 3017 1852 3046 1857
rect 209 1847 542 1852
rect 2241 1847 2326 1852
rect 121 1842 150 1847
rect 185 1842 214 1847
rect 537 1842 1334 1847
rect 1345 1842 1438 1847
rect 1465 1842 1510 1847
rect 1577 1842 2046 1847
rect 2073 1842 2118 1847
rect 2129 1842 2174 1847
rect 2321 1842 2886 1847
rect 3065 1842 3166 1847
rect 3185 1842 3206 1847
rect 2905 1837 3070 1842
rect 3161 1837 3166 1842
rect 65 1832 134 1837
rect 209 1832 238 1837
rect 273 1832 654 1837
rect 785 1832 918 1837
rect 945 1832 1478 1837
rect 1633 1832 1662 1837
rect 1681 1832 1710 1837
rect 1817 1832 2910 1837
rect 3161 1832 3206 1837
rect 81 1822 150 1827
rect 225 1822 254 1827
rect 217 1812 278 1817
rect 353 1812 358 1832
rect 673 1827 766 1832
rect 1705 1827 1822 1832
rect 409 1822 534 1827
rect 545 1822 678 1827
rect 761 1822 838 1827
rect 921 1822 1046 1827
rect 1065 1822 1662 1827
rect 1841 1822 1982 1827
rect 2009 1822 2686 1827
rect 2697 1822 2734 1827
rect 2753 1822 2854 1827
rect 2865 1822 3102 1827
rect 545 1817 550 1822
rect 2865 1817 2870 1822
rect 433 1812 518 1817
rect 529 1812 550 1817
rect 569 1812 670 1817
rect 729 1812 750 1817
rect 793 1812 814 1817
rect 833 1812 1230 1817
rect 1241 1812 1350 1817
rect 1377 1812 1398 1817
rect 1505 1812 1534 1817
rect 1633 1812 1846 1817
rect 1905 1812 2038 1817
rect 2145 1812 2198 1817
rect 2273 1812 2374 1817
rect 2489 1812 2870 1817
rect 2889 1812 3158 1817
rect 3177 1812 3230 1817
rect 193 1802 270 1807
rect 505 1802 598 1807
rect 673 1802 726 1807
rect 833 1802 838 1812
rect 1529 1807 1638 1812
rect 1841 1807 1846 1812
rect 849 1802 1462 1807
rect 1657 1802 1782 1807
rect 1841 1802 1862 1807
rect 2137 1802 2246 1807
rect 353 1797 486 1802
rect 1457 1797 1462 1802
rect 1857 1797 1862 1802
rect 2009 1797 2118 1802
rect 2241 1797 2246 1802
rect 2273 1797 2278 1812
rect 2353 1802 2422 1807
rect 2433 1802 2470 1807
rect 2481 1802 2534 1807
rect 2577 1802 2622 1807
rect 2689 1802 2798 1807
rect 2945 1802 3102 1807
rect 2353 1797 2358 1802
rect 2481 1797 2486 1802
rect 2945 1797 2950 1802
rect 3153 1797 3158 1812
rect 3185 1802 3270 1807
rect 3345 1802 3422 1807
rect 3265 1797 3270 1802
rect 113 1792 190 1797
rect 233 1792 286 1797
rect 329 1792 358 1797
rect 481 1792 886 1797
rect 913 1792 958 1797
rect 985 1792 1110 1797
rect 1137 1792 1214 1797
rect 1257 1792 1446 1797
rect 1457 1792 1526 1797
rect 1585 1792 1710 1797
rect 1745 1792 1838 1797
rect 1857 1792 1942 1797
rect 1985 1792 2014 1797
rect 2113 1792 2222 1797
rect 2241 1792 2278 1797
rect 2305 1792 2358 1797
rect 2377 1792 2486 1797
rect 2497 1792 2614 1797
rect 2649 1792 2694 1797
rect 2729 1792 2766 1797
rect 2833 1792 2950 1797
rect 3009 1792 3126 1797
rect 3153 1792 3230 1797
rect 3265 1792 3294 1797
rect 1105 1787 1110 1792
rect 145 1782 174 1787
rect 337 1782 822 1787
rect 857 1782 926 1787
rect 1105 1782 1206 1787
rect 1233 1782 1310 1787
rect 1353 1782 1582 1787
rect 1601 1782 1726 1787
rect 1737 1782 1822 1787
rect 1833 1782 1910 1787
rect 1929 1782 2958 1787
rect 2969 1782 3038 1787
rect 953 1777 1086 1782
rect 321 1772 350 1777
rect 465 1772 958 1777
rect 1081 1772 1270 1777
rect 1353 1772 1614 1777
rect 1657 1772 1710 1777
rect 1729 1772 2142 1777
rect 2201 1772 2398 1777
rect 2465 1772 2502 1777
rect 2537 1772 2750 1777
rect 2849 1772 2878 1777
rect 3217 1772 3246 1777
rect 345 1767 470 1772
rect 1265 1767 1358 1772
rect 489 1762 526 1767
rect 545 1762 574 1767
rect 585 1762 918 1767
rect 945 1762 1102 1767
rect 1113 1762 1246 1767
rect 1377 1762 1422 1767
rect 1465 1762 1510 1767
rect 1521 1762 1694 1767
rect 1753 1762 1798 1767
rect 1817 1762 1958 1767
rect 2081 1762 2126 1767
rect 2145 1762 2222 1767
rect 2233 1762 2294 1767
rect 2313 1762 2702 1767
rect 2753 1762 2790 1767
rect 2825 1762 2854 1767
rect 2881 1762 2990 1767
rect 3177 1762 3398 1767
rect 2289 1757 2294 1762
rect 201 1752 238 1757
rect 401 1752 462 1757
rect 641 1752 1230 1757
rect 1297 1752 1366 1757
rect 1401 1752 1630 1757
rect 1689 1752 2014 1757
rect 2025 1752 2174 1757
rect 2241 1752 2278 1757
rect 2289 1752 2334 1757
rect 2361 1752 2398 1757
rect 2441 1752 2494 1757
rect 2553 1752 2598 1757
rect 2721 1752 2742 1757
rect 2785 1752 2830 1757
rect 2905 1752 2998 1757
rect 3257 1752 3310 1757
rect 3409 1752 3438 1757
rect 3305 1747 3414 1752
rect 217 1742 294 1747
rect 337 1742 422 1747
rect 489 1742 518 1747
rect 537 1742 614 1747
rect 649 1742 846 1747
rect 889 1742 1318 1747
rect 1449 1742 1670 1747
rect 1785 1742 1806 1747
rect 1865 1742 2054 1747
rect 2065 1742 2174 1747
rect 2193 1742 2926 1747
rect 2969 1742 3086 1747
rect 3209 1742 3286 1747
rect 609 1737 614 1742
rect 1313 1737 1454 1742
rect 2193 1737 2198 1742
rect 321 1732 366 1737
rect 385 1732 526 1737
rect 609 1732 646 1737
rect 673 1732 750 1737
rect 833 1732 966 1737
rect 1001 1732 1086 1737
rect 1161 1732 1294 1737
rect 1473 1732 1590 1737
rect 1657 1732 1702 1737
rect 1841 1732 1878 1737
rect 1889 1732 1966 1737
rect 2017 1732 2198 1737
rect 2241 1732 3006 1737
rect 3041 1732 3062 1737
rect 3233 1732 3366 1737
rect 129 1722 358 1727
rect 513 1722 582 1727
rect 673 1722 678 1732
rect 1721 1727 1822 1732
rect 689 1722 742 1727
rect 785 1722 942 1727
rect 953 1722 1390 1727
rect 1449 1722 1606 1727
rect 1625 1722 1726 1727
rect 1817 1722 3302 1727
rect 137 1712 198 1717
rect 273 1712 326 1717
rect 393 1712 1526 1717
rect 1729 1712 1782 1717
rect 1793 1712 1870 1717
rect 1897 1712 1982 1717
rect 2009 1712 2166 1717
rect 2345 1712 2366 1717
rect 2433 1712 2462 1717
rect 2473 1712 2550 1717
rect 2665 1712 2742 1717
rect 2825 1712 2870 1717
rect 2961 1712 3230 1717
rect 2961 1707 2966 1712
rect 209 1702 390 1707
rect 417 1702 446 1707
rect 505 1702 686 1707
rect 729 1702 806 1707
rect 865 1702 1022 1707
rect 1049 1702 1086 1707
rect 1097 1702 1318 1707
rect 1417 1702 1510 1707
rect 1585 1702 1694 1707
rect 1737 1702 2246 1707
rect 2337 1702 2502 1707
rect 2593 1702 2702 1707
rect 2801 1702 2966 1707
rect 2985 1702 3190 1707
rect 3209 1702 3278 1707
rect 289 1692 318 1697
rect 441 1692 574 1697
rect 697 1692 774 1697
rect 817 1692 998 1697
rect 1017 1692 1118 1697
rect 1129 1692 1158 1697
rect 1169 1692 1214 1697
rect 1449 1692 1718 1697
rect 1825 1692 2206 1697
rect 2401 1692 2422 1697
rect 2465 1692 2614 1697
rect 2697 1692 2814 1697
rect 2945 1692 2990 1697
rect 3073 1692 3110 1697
rect 313 1687 446 1692
rect 2401 1687 2406 1692
rect 137 1682 222 1687
rect 465 1682 1302 1687
rect 1321 1682 1422 1687
rect 1441 1682 1534 1687
rect 1577 1682 1638 1687
rect 1713 1682 1750 1687
rect 1833 1682 1910 1687
rect 1961 1682 2118 1687
rect 2185 1682 2222 1687
rect 2345 1682 2406 1687
rect 2609 1682 2646 1687
rect 1321 1677 1326 1682
rect 89 1672 126 1677
rect 121 1667 126 1672
rect 185 1672 326 1677
rect 417 1672 502 1677
rect 537 1672 702 1677
rect 761 1672 886 1677
rect 897 1672 1030 1677
rect 1121 1672 1326 1677
rect 1417 1677 1422 1682
rect 2641 1677 2646 1682
rect 2729 1682 2758 1687
rect 3041 1682 3158 1687
rect 2729 1677 2734 1682
rect 1417 1672 2446 1677
rect 2465 1672 2582 1677
rect 2641 1672 2734 1677
rect 2761 1672 2822 1677
rect 3065 1672 3134 1677
rect 185 1667 190 1672
rect 897 1667 902 1672
rect 2465 1667 2470 1672
rect 121 1662 190 1667
rect 225 1662 294 1667
rect 409 1662 782 1667
rect 841 1662 902 1667
rect 929 1662 1166 1667
rect 1297 1662 1334 1667
rect 1345 1662 1422 1667
rect 1505 1662 1606 1667
rect 1617 1662 1798 1667
rect 1905 1662 1950 1667
rect 1985 1662 2054 1667
rect 2129 1662 2374 1667
rect 2417 1662 2470 1667
rect 2577 1667 2582 1672
rect 2577 1662 2622 1667
rect 3169 1662 3342 1667
rect 289 1657 294 1662
rect 1185 1657 1270 1662
rect 1601 1657 1606 1662
rect 2417 1657 2422 1662
rect 209 1652 270 1657
rect 289 1652 422 1657
rect 513 1652 1190 1657
rect 1265 1652 1454 1657
rect 1473 1652 1534 1657
rect 1601 1652 1694 1657
rect 1705 1652 2014 1657
rect 2033 1652 2062 1657
rect 2137 1652 2294 1657
rect 2329 1652 2422 1657
rect 2465 1652 2566 1657
rect 2873 1652 3046 1657
rect 3073 1652 3206 1657
rect 417 1647 518 1652
rect 129 1642 230 1647
rect 297 1642 398 1647
rect 537 1642 654 1647
rect 665 1642 702 1647
rect 889 1642 1078 1647
rect 1201 1642 1254 1647
rect 1369 1642 1766 1647
rect 1857 1642 2574 1647
rect 2641 1642 2830 1647
rect 721 1637 814 1642
rect 1761 1637 1862 1642
rect 2641 1637 2646 1642
rect 169 1632 222 1637
rect 305 1632 438 1637
rect 601 1632 726 1637
rect 809 1632 838 1637
rect 913 1632 998 1637
rect 1033 1632 1070 1637
rect 1305 1632 1390 1637
rect 1481 1632 1502 1637
rect 1529 1632 1558 1637
rect 1577 1632 1742 1637
rect 1881 1632 1966 1637
rect 2073 1632 2102 1637
rect 2233 1632 2318 1637
rect 2345 1632 2374 1637
rect 2409 1632 2646 1637
rect 2825 1637 2830 1642
rect 2873 1637 2878 1652
rect 2825 1632 2878 1637
rect 3041 1637 3046 1652
rect 3041 1632 3078 1637
rect 465 1627 582 1632
rect 993 1627 998 1632
rect 2097 1627 2238 1632
rect 89 1622 174 1627
rect 201 1622 310 1627
rect 369 1622 470 1627
rect 577 1622 926 1627
rect 993 1622 1054 1627
rect 1185 1622 1238 1627
rect 1313 1617 1318 1627
rect 1449 1622 1550 1627
rect 1657 1622 2070 1627
rect 2257 1622 2486 1627
rect 2521 1622 2654 1627
rect 2689 1622 2710 1627
rect 2801 1622 2878 1627
rect 2921 1622 2974 1627
rect 3009 1622 3062 1627
rect 1545 1617 1662 1622
rect 2257 1617 2262 1622
rect 2481 1617 2486 1622
rect 65 1612 142 1617
rect 185 1612 214 1617
rect 481 1612 590 1617
rect 625 1612 830 1617
rect 929 1612 1038 1617
rect 1185 1612 1230 1617
rect 1313 1612 1430 1617
rect 1465 1612 1526 1617
rect 65 1607 70 1612
rect 209 1607 214 1612
rect 313 1607 462 1612
rect 825 1607 934 1612
rect 1681 1607 1686 1617
rect 1697 1612 1806 1617
rect 1889 1612 1942 1617
rect 2017 1612 2262 1617
rect 2273 1612 2470 1617
rect 2481 1612 3038 1617
rect 3073 1607 3078 1632
rect 3169 1622 3262 1627
rect 3089 1612 3422 1617
rect 65 1602 94 1607
rect 113 1602 150 1607
rect 209 1602 270 1607
rect 289 1602 318 1607
rect 457 1602 534 1607
rect 745 1602 806 1607
rect 953 1602 982 1607
rect 1105 1602 1198 1607
rect 1321 1602 1686 1607
rect 1745 1602 1774 1607
rect 1897 1602 2142 1607
rect 2153 1602 2326 1607
rect 2345 1602 2430 1607
rect 2449 1602 2614 1607
rect 2721 1602 2766 1607
rect 2849 1602 2974 1607
rect 2985 1602 3038 1607
rect 3073 1602 3270 1607
rect 81 1592 134 1597
rect 145 1577 150 1602
rect 289 1597 294 1602
rect 553 1597 662 1602
rect 2321 1597 2326 1602
rect 2449 1597 2454 1602
rect 2609 1597 2614 1602
rect 257 1592 294 1597
rect 313 1592 558 1597
rect 657 1592 686 1597
rect 737 1592 822 1597
rect 865 1592 942 1597
rect 953 1592 1006 1597
rect 1137 1592 1342 1597
rect 1665 1592 1726 1597
rect 1801 1592 1934 1597
rect 1969 1592 2006 1597
rect 2025 1592 2054 1597
rect 2185 1592 2262 1597
rect 2321 1592 2454 1597
rect 2489 1592 2598 1597
rect 2609 1592 2710 1597
rect 2777 1592 2870 1597
rect 2889 1592 3142 1597
rect 3217 1592 3286 1597
rect 3297 1592 3398 1597
rect 737 1587 742 1592
rect 1369 1587 1478 1592
rect 1969 1587 1974 1592
rect 2705 1587 2782 1592
rect 2865 1587 2870 1592
rect 3281 1587 3286 1592
rect 305 1582 398 1587
rect 449 1582 502 1587
rect 545 1582 598 1587
rect 625 1582 766 1587
rect 785 1582 1006 1587
rect 1025 1582 1118 1587
rect 1169 1582 1270 1587
rect 1345 1582 1374 1587
rect 1473 1582 1566 1587
rect 1657 1582 1758 1587
rect 1825 1582 1854 1587
rect 1905 1582 1974 1587
rect 2001 1582 2078 1587
rect 2129 1582 2214 1587
rect 2241 1582 2342 1587
rect 2393 1582 2422 1587
rect 2441 1582 2526 1587
rect 2865 1582 2910 1587
rect 2961 1582 3094 1587
rect 3281 1582 3334 1587
rect 1025 1577 1030 1582
rect 121 1572 150 1577
rect 305 1572 334 1577
rect 353 1572 806 1577
rect 889 1572 950 1577
rect 977 1572 1030 1577
rect 1113 1577 1118 1582
rect 1113 1572 1462 1577
rect 1681 1572 1782 1577
rect 1849 1572 1918 1577
rect 1937 1572 2022 1577
rect 2089 1572 2134 1577
rect 2145 1572 2222 1577
rect 2241 1572 2294 1577
rect 2305 1572 2462 1577
rect 2489 1572 2510 1577
rect 2593 1572 2638 1577
rect 2729 1572 2830 1577
rect 3001 1572 3102 1577
rect 3361 1572 3430 1577
rect 145 1567 150 1572
rect 2729 1567 2734 1572
rect 145 1562 238 1567
rect 289 1562 326 1567
rect 361 1562 734 1567
rect 817 1562 1158 1567
rect 1209 1562 1294 1567
rect 1313 1562 1398 1567
rect 1737 1562 2734 1567
rect 2825 1567 2830 1572
rect 2825 1562 2854 1567
rect 3185 1562 3278 1567
rect 233 1557 238 1562
rect 233 1552 622 1557
rect 705 1552 814 1557
rect 921 1552 1174 1557
rect 1209 1552 1254 1557
rect 1273 1552 1390 1557
rect 1521 1552 1614 1557
rect 1625 1552 1670 1557
rect 1721 1552 1838 1557
rect 1897 1552 2006 1557
rect 2025 1552 2534 1557
rect 2569 1552 2638 1557
rect 2745 1552 2934 1557
rect 2945 1552 3070 1557
rect 3241 1552 3278 1557
rect 3313 1552 3342 1557
rect 809 1547 926 1552
rect 2001 1547 2006 1552
rect 2945 1547 2950 1552
rect 49 1542 134 1547
rect 297 1542 366 1547
rect 377 1542 438 1547
rect 473 1542 494 1547
rect 553 1542 622 1547
rect 673 1542 726 1547
rect 737 1542 790 1547
rect 945 1542 1030 1547
rect 1097 1542 1134 1547
rect 1225 1542 1262 1547
rect 1329 1542 1374 1547
rect 1529 1542 1942 1547
rect 2001 1542 2782 1547
rect 2873 1542 2950 1547
rect 3281 1542 3310 1547
rect 3321 1542 3350 1547
rect 49 1407 54 1542
rect 2777 1537 2878 1542
rect 153 1532 222 1537
rect 593 1532 894 1537
rect 905 1532 1126 1537
rect 1161 1532 1270 1537
rect 1281 1532 1350 1537
rect 1409 1532 1502 1537
rect 1681 1532 1774 1537
rect 1785 1532 2206 1537
rect 2257 1532 2366 1537
rect 2385 1532 2614 1537
rect 2657 1532 2686 1537
rect 2713 1532 2758 1537
rect 2937 1532 2990 1537
rect 297 1527 542 1532
rect 1409 1527 1414 1532
rect 1497 1527 1646 1532
rect 2657 1527 2662 1532
rect 129 1522 158 1527
rect 153 1517 158 1522
rect 233 1522 302 1527
rect 537 1522 566 1527
rect 585 1522 1006 1527
rect 1105 1522 1414 1527
rect 1641 1522 2510 1527
rect 2521 1522 2662 1527
rect 2681 1522 2854 1527
rect 2881 1522 3030 1527
rect 3273 1522 3374 1527
rect 233 1517 238 1522
rect 561 1517 566 1522
rect 3273 1517 3278 1522
rect 113 1487 118 1517
rect 153 1512 238 1517
rect 313 1512 502 1517
rect 561 1512 1630 1517
rect 1721 1512 1822 1517
rect 1865 1512 2758 1517
rect 2769 1512 3086 1517
rect 3185 1512 3278 1517
rect 3369 1517 3374 1522
rect 3369 1512 3398 1517
rect 497 1507 502 1512
rect 2769 1507 2774 1512
rect 281 1502 478 1507
rect 497 1502 558 1507
rect 577 1502 622 1507
rect 817 1502 1542 1507
rect 1633 1502 1790 1507
rect 1849 1502 1990 1507
rect 2033 1502 2062 1507
rect 2081 1502 2774 1507
rect 2833 1502 3006 1507
rect 681 1497 750 1502
rect 3001 1497 3006 1502
rect 3065 1502 3206 1507
rect 3289 1502 3438 1507
rect 3065 1497 3070 1502
rect 281 1492 646 1497
rect 657 1492 686 1497
rect 745 1492 814 1497
rect 873 1492 1094 1497
rect 1121 1492 1142 1497
rect 1249 1492 1742 1497
rect 1753 1492 1926 1497
rect 1953 1492 2014 1497
rect 2057 1492 2078 1497
rect 2097 1492 2134 1497
rect 2209 1492 2254 1497
rect 2305 1492 2334 1497
rect 2345 1492 2446 1497
rect 2481 1492 2566 1497
rect 2681 1492 2766 1497
rect 3001 1492 3070 1497
rect 641 1487 646 1492
rect 81 1482 118 1487
rect 217 1482 246 1487
rect 329 1482 358 1487
rect 409 1482 534 1487
rect 601 1482 630 1487
rect 641 1482 734 1487
rect 897 1482 926 1487
rect 1025 1482 1294 1487
rect 1345 1482 2470 1487
rect 241 1477 334 1482
rect 729 1477 902 1482
rect 2465 1477 2470 1482
rect 2553 1482 2582 1487
rect 3089 1482 3198 1487
rect 2553 1477 2558 1482
rect 2737 1477 2830 1482
rect 65 1472 134 1477
rect 417 1472 494 1477
rect 577 1472 598 1477
rect 1033 1472 1142 1477
rect 1201 1472 1254 1477
rect 1521 1472 1574 1477
rect 1697 1472 1854 1477
rect 1937 1472 2054 1477
rect 2065 1472 2422 1477
rect 2465 1472 2558 1477
rect 2713 1472 2742 1477
rect 2825 1472 2854 1477
rect 617 1467 710 1472
rect 1137 1467 1142 1472
rect 1273 1467 1502 1472
rect 2065 1467 2070 1472
rect 89 1462 238 1467
rect 297 1462 342 1467
rect 377 1462 430 1467
rect 449 1462 518 1467
rect 529 1462 622 1467
rect 705 1462 734 1467
rect 777 1462 830 1467
rect 961 1462 990 1467
rect 1041 1462 1118 1467
rect 1137 1462 1278 1467
rect 1497 1462 1558 1467
rect 1769 1462 1942 1467
rect 1953 1462 2070 1467
rect 2137 1462 2342 1467
rect 2761 1462 2886 1467
rect 2993 1462 3030 1467
rect 1609 1457 1750 1462
rect 2641 1457 2742 1462
rect 241 1452 326 1457
rect 377 1452 478 1457
rect 497 1452 710 1457
rect 873 1452 1614 1457
rect 1745 1452 2446 1457
rect 2617 1452 2646 1457
rect 2737 1452 2846 1457
rect 3009 1452 3062 1457
rect 177 1442 206 1447
rect 257 1442 310 1447
rect 337 1442 414 1447
rect 457 1442 574 1447
rect 81 1432 142 1437
rect 177 1427 182 1442
rect 625 1437 630 1447
rect 641 1442 806 1447
rect 881 1442 1414 1447
rect 1433 1442 1542 1447
rect 1617 1442 1886 1447
rect 1961 1442 2054 1447
rect 2065 1442 2174 1447
rect 2233 1442 2270 1447
rect 2289 1442 2310 1447
rect 2393 1442 2414 1447
rect 2433 1442 2502 1447
rect 2537 1442 2870 1447
rect 2945 1442 3078 1447
rect 3137 1442 3230 1447
rect 2945 1437 2950 1442
rect 193 1432 222 1437
rect 393 1432 630 1437
rect 665 1432 750 1437
rect 865 1432 1022 1437
rect 1049 1432 1270 1437
rect 1329 1432 1582 1437
rect 1713 1432 1934 1437
rect 1985 1432 2294 1437
rect 2305 1432 2950 1437
rect 2961 1432 3014 1437
rect 217 1427 398 1432
rect 2305 1427 2310 1432
rect 113 1422 150 1427
rect 177 1422 198 1427
rect 417 1422 438 1427
rect 497 1422 590 1427
rect 793 1422 918 1427
rect 929 1422 966 1427
rect 977 1422 1078 1427
rect 1153 1422 1294 1427
rect 1313 1422 1406 1427
rect 1449 1422 1494 1427
rect 145 1407 150 1422
rect 193 1417 198 1422
rect 681 1417 774 1422
rect 1073 1417 1078 1422
rect 1313 1417 1318 1422
rect 1681 1417 1686 1427
rect 1977 1422 2126 1427
rect 2153 1422 2310 1427
rect 2345 1422 2374 1427
rect 2465 1422 2654 1427
rect 2745 1422 2774 1427
rect 2937 1422 2966 1427
rect 3041 1422 3062 1427
rect 3185 1422 3302 1427
rect 3385 1422 3414 1427
rect 1833 1417 1902 1422
rect 2769 1417 2942 1422
rect 3185 1417 3190 1422
rect 193 1412 238 1417
rect 265 1412 326 1417
rect 385 1412 478 1417
rect 513 1412 646 1417
rect 657 1412 686 1417
rect 769 1412 1006 1417
rect 1073 1412 1126 1417
rect 1185 1412 1318 1417
rect 1345 1412 1446 1417
rect 1457 1412 1502 1417
rect 1569 1412 1838 1417
rect 1897 1412 2358 1417
rect 2401 1412 2622 1417
rect 3001 1412 3046 1417
rect 3145 1412 3190 1417
rect 321 1407 326 1412
rect 657 1407 662 1412
rect 2353 1407 2358 1412
rect 49 1402 70 1407
rect 89 1402 118 1407
rect 145 1402 166 1407
rect 257 1402 302 1407
rect 321 1402 662 1407
rect 721 1402 814 1407
rect 849 1402 1062 1407
rect 1137 1402 1558 1407
rect 1721 1402 1750 1407
rect 1849 1402 1886 1407
rect 1985 1402 2262 1407
rect 2297 1402 2334 1407
rect 2353 1402 2678 1407
rect 2697 1402 2766 1407
rect 2833 1402 2894 1407
rect 2905 1402 2942 1407
rect 3161 1402 3294 1407
rect 161 1397 166 1402
rect 81 1392 142 1397
rect 161 1392 214 1397
rect 249 1392 310 1397
rect 353 1392 574 1397
rect 689 1392 838 1397
rect 849 1387 854 1402
rect 1553 1397 1726 1402
rect 977 1392 1166 1397
rect 1177 1392 1310 1397
rect 1361 1392 1390 1397
rect 1417 1392 1478 1397
rect 1785 1392 1870 1397
rect 1913 1392 2982 1397
rect 3241 1392 3294 1397
rect 3321 1392 3406 1397
rect 1177 1387 1182 1392
rect 89 1382 198 1387
rect 225 1382 694 1387
rect 713 1382 742 1387
rect 769 1382 854 1387
rect 921 1382 1038 1387
rect 1065 1382 1086 1387
rect 1121 1382 1182 1387
rect 1193 1382 1558 1387
rect 1609 1382 1750 1387
rect 1833 1382 2150 1387
rect 2233 1382 2438 1387
rect 2465 1382 2502 1387
rect 2561 1382 2822 1387
rect 2841 1382 3038 1387
rect 3233 1382 3422 1387
rect 737 1377 742 1382
rect 1609 1377 1614 1382
rect 337 1372 358 1377
rect 377 1372 414 1377
rect 545 1372 726 1377
rect 737 1372 838 1377
rect 969 1372 1086 1377
rect 1113 1372 1542 1377
rect 1585 1372 1614 1377
rect 1745 1377 1750 1382
rect 2817 1377 2822 1382
rect 1745 1372 2142 1377
rect 2249 1372 2358 1377
rect 2369 1372 2654 1377
rect 2681 1372 2718 1377
rect 2817 1372 2926 1377
rect 3017 1372 3062 1377
rect 3177 1372 3270 1377
rect 433 1367 510 1372
rect 1537 1367 1542 1372
rect 2353 1367 2358 1372
rect 305 1362 438 1367
rect 505 1362 822 1367
rect 1001 1362 1126 1367
rect 1177 1362 1286 1367
rect 1321 1362 1526 1367
rect 1537 1362 1630 1367
rect 1649 1362 1734 1367
rect 1849 1362 1894 1367
rect 1969 1362 2126 1367
rect 2193 1362 2238 1367
rect 2289 1362 2342 1367
rect 2353 1362 2390 1367
rect 2441 1362 2502 1367
rect 2537 1362 2662 1367
rect 2721 1362 2822 1367
rect 2833 1362 2910 1367
rect 2921 1362 3014 1367
rect 1281 1357 1286 1362
rect 1649 1357 1654 1362
rect 2497 1357 2502 1362
rect 3009 1357 3014 1362
rect 3073 1362 3102 1367
rect 3073 1357 3078 1362
rect 185 1352 494 1357
rect 561 1352 926 1357
rect 937 1352 1198 1357
rect 1233 1352 1262 1357
rect 1281 1352 1654 1357
rect 1721 1352 1926 1357
rect 1937 1352 2086 1357
rect 2105 1352 2486 1357
rect 2497 1352 2814 1357
rect 2905 1352 2990 1357
rect 3009 1352 3078 1357
rect 3233 1352 3286 1357
rect 81 1342 158 1347
rect 337 1342 430 1347
rect 609 1342 630 1347
rect 689 1342 910 1347
rect 953 1342 1022 1347
rect 1097 1342 1614 1347
rect 1801 1342 1838 1347
rect 1921 1342 1926 1352
rect 2481 1347 2486 1352
rect 2041 1342 2174 1347
rect 2265 1342 2286 1347
rect 2305 1342 2390 1347
rect 2409 1342 2462 1347
rect 2481 1342 2566 1347
rect 2625 1342 2742 1347
rect 2761 1342 2870 1347
rect 3153 1342 3270 1347
rect 1609 1337 1710 1342
rect 1801 1337 1806 1342
rect 1921 1337 2022 1342
rect 2785 1337 2790 1342
rect 201 1332 230 1337
rect 225 1327 230 1332
rect 289 1332 318 1337
rect 385 1332 422 1337
rect 585 1332 646 1337
rect 705 1332 742 1337
rect 793 1332 822 1337
rect 937 1332 1030 1337
rect 1137 1332 1158 1337
rect 1185 1332 1326 1337
rect 1361 1332 1478 1337
rect 1561 1332 1590 1337
rect 1705 1332 1806 1337
rect 2017 1332 2646 1337
rect 2761 1332 2790 1337
rect 2841 1332 2982 1337
rect 3193 1332 3350 1337
rect 289 1327 294 1332
rect 817 1327 942 1332
rect 1361 1327 1366 1332
rect 1473 1327 1566 1332
rect 2641 1327 2766 1332
rect 225 1322 294 1327
rect 593 1322 726 1327
rect 961 1322 1366 1327
rect 1385 1322 1438 1327
rect 1601 1322 1662 1327
rect 1825 1322 2046 1327
rect 2153 1322 2310 1327
rect 2385 1322 2462 1327
rect 2545 1322 2622 1327
rect 2961 1322 3038 1327
rect 3201 1322 3270 1327
rect 2785 1317 2966 1322
rect 625 1312 854 1317
rect 953 1312 1614 1317
rect 1673 1312 1918 1317
rect 2129 1312 2214 1317
rect 2265 1312 2398 1317
rect 2449 1312 2790 1317
rect 2985 1312 3190 1317
rect 105 1302 206 1307
rect 505 1302 574 1307
rect 705 1302 734 1307
rect 929 1302 974 1307
rect 1081 1302 1166 1307
rect 1361 1302 1422 1307
rect 1449 1302 1486 1307
rect 1585 1302 1590 1312
rect 1609 1307 1678 1312
rect 1937 1307 2110 1312
rect 1801 1302 1942 1307
rect 2105 1302 2406 1307
rect 2417 1302 2582 1307
rect 2745 1302 3046 1307
rect 105 1297 110 1302
rect 81 1292 110 1297
rect 201 1297 206 1302
rect 201 1292 230 1297
rect 449 1292 510 1297
rect 705 1292 710 1302
rect 849 1292 950 1297
rect 1073 1292 1142 1297
rect 1193 1292 1222 1297
rect 1241 1292 1310 1297
rect 1409 1292 1638 1297
rect 1657 1292 1758 1297
rect 1865 1292 2150 1297
rect 2193 1292 2310 1297
rect 2321 1292 2734 1297
rect 2793 1292 2966 1297
rect 1241 1287 1246 1292
rect 105 1282 294 1287
rect 409 1282 558 1287
rect 985 1282 1246 1287
rect 1305 1287 1310 1292
rect 1657 1287 1662 1292
rect 1305 1282 1398 1287
rect 1553 1282 1662 1287
rect 1753 1287 1758 1292
rect 2321 1287 2326 1292
rect 2729 1287 2798 1292
rect 1753 1282 1902 1287
rect 1913 1282 2326 1287
rect 2385 1282 2518 1287
rect 1393 1277 1558 1282
rect 209 1272 238 1277
rect 305 1272 398 1277
rect 569 1272 598 1277
rect 801 1272 918 1277
rect 977 1272 1102 1277
rect 1121 1272 1294 1277
rect 1577 1272 1742 1277
rect 1865 1272 1894 1277
rect 1921 1272 2614 1277
rect 2633 1272 2758 1277
rect 233 1267 310 1272
rect 393 1267 574 1272
rect 1737 1267 1870 1272
rect 609 1262 790 1267
rect 881 1262 1030 1267
rect 1153 1262 1510 1267
rect 1665 1262 1718 1267
rect 233 1252 302 1257
rect 369 1252 390 1257
rect 409 1252 534 1257
rect 409 1247 414 1252
rect 369 1242 414 1247
rect 529 1247 534 1252
rect 609 1247 614 1262
rect 785 1257 886 1262
rect 1025 1257 1158 1262
rect 1921 1257 1926 1272
rect 2633 1267 2638 1272
rect 1977 1262 2406 1267
rect 2433 1262 2638 1267
rect 2753 1267 2758 1272
rect 2753 1262 2878 1267
rect 905 1252 1006 1257
rect 1177 1252 1302 1257
rect 1457 1252 1654 1257
rect 1713 1252 1926 1257
rect 1937 1252 2110 1257
rect 2217 1252 2238 1257
rect 2249 1252 2286 1257
rect 2305 1252 2366 1257
rect 2441 1252 2470 1257
rect 2481 1252 2518 1257
rect 2641 1252 2742 1257
rect 2993 1252 3062 1257
rect 1329 1247 1438 1252
rect 529 1242 614 1247
rect 665 1242 718 1247
rect 817 1242 942 1247
rect 1057 1242 1110 1247
rect 1201 1242 1334 1247
rect 1433 1242 1582 1247
rect 1601 1242 2998 1247
rect 2993 1237 2998 1242
rect 145 1232 518 1237
rect 585 1232 670 1237
rect 753 1232 814 1237
rect 1041 1232 1150 1237
rect 1201 1232 1238 1237
rect 1345 1232 1566 1237
rect 1745 1232 1918 1237
rect 2065 1232 2198 1237
rect 2209 1232 2246 1237
rect 2257 1232 2342 1237
rect 2369 1232 2542 1237
rect 2673 1232 2766 1237
rect 2993 1232 3086 1237
rect 3161 1232 3310 1237
rect 105 1222 198 1227
rect 433 1222 1086 1227
rect 1241 1222 1326 1227
rect 137 1212 278 1217
rect 329 1212 414 1217
rect 153 1202 182 1207
rect 329 1202 422 1207
rect 177 1197 182 1202
rect 241 1197 334 1202
rect 433 1197 438 1222
rect 1345 1217 1350 1232
rect 1537 1227 1542 1232
rect 1585 1227 1726 1232
rect 1745 1227 1750 1232
rect 1937 1227 2046 1232
rect 2561 1227 2654 1232
rect 1377 1222 1462 1227
rect 1537 1222 1590 1227
rect 1721 1222 1774 1227
rect 1793 1222 1942 1227
rect 2041 1222 2470 1227
rect 2521 1222 2566 1227
rect 2649 1222 2678 1227
rect 2777 1222 2934 1227
rect 3041 1222 3118 1227
rect 3169 1222 3206 1227
rect 2673 1217 2782 1222
rect 513 1212 654 1217
rect 721 1212 758 1217
rect 769 1212 814 1217
rect 1169 1212 1350 1217
rect 1417 1212 2654 1217
rect 2817 1212 2846 1217
rect 2945 1212 3062 1217
rect 3121 1212 3190 1217
rect 3329 1212 3334 1237
rect 753 1207 758 1212
rect 833 1207 934 1212
rect 993 1207 1150 1212
rect 2841 1207 2950 1212
rect 457 1202 566 1207
rect 753 1202 838 1207
rect 929 1202 958 1207
rect 969 1202 998 1207
rect 1145 1202 1630 1207
rect 1745 1202 1822 1207
rect 1881 1202 2014 1207
rect 2057 1202 2142 1207
rect 2161 1202 2230 1207
rect 2305 1202 2518 1207
rect 2665 1202 2718 1207
rect 2537 1197 2638 1202
rect 177 1192 246 1197
rect 353 1192 414 1197
rect 433 1192 478 1197
rect 489 1192 990 1197
rect 1001 1192 1526 1197
rect 313 1182 526 1187
rect 705 1182 798 1187
rect 865 1182 966 1187
rect 1105 1182 1262 1187
rect 1369 1182 1510 1187
rect 977 1177 1110 1182
rect 1257 1177 1374 1182
rect 1521 1177 1526 1192
rect 1553 1192 2542 1197
rect 2633 1192 2662 1197
rect 2737 1192 2806 1197
rect 2865 1192 3006 1197
rect 3193 1192 3302 1197
rect 1553 1187 1558 1192
rect 2737 1187 2742 1192
rect 1537 1182 1558 1187
rect 1601 1182 2742 1187
rect 2801 1187 2806 1192
rect 2801 1182 2830 1187
rect 2977 1182 3006 1187
rect 3025 1182 3094 1187
rect 3201 1182 3270 1187
rect 3025 1177 3030 1182
rect 265 1172 358 1177
rect 377 1172 494 1177
rect 561 1172 622 1177
rect 681 1172 982 1177
rect 1129 1172 1238 1177
rect 1521 1172 1822 1177
rect 1913 1172 2822 1177
rect 2849 1172 2950 1177
rect 2969 1172 3030 1177
rect 3089 1177 3094 1182
rect 3089 1172 3118 1177
rect 561 1167 566 1172
rect 2849 1167 2854 1172
rect 113 1162 190 1167
rect 289 1162 318 1167
rect 417 1162 566 1167
rect 585 1162 614 1167
rect 777 1162 838 1167
rect 865 1162 950 1167
rect 1017 1162 1934 1167
rect 1969 1162 2126 1167
rect 2153 1162 2198 1167
rect 2217 1162 2262 1167
rect 2321 1162 2342 1167
rect 2401 1162 2470 1167
rect 2585 1162 2854 1167
rect 2945 1167 2950 1172
rect 2945 1162 3134 1167
rect 313 1157 422 1162
rect 609 1157 782 1162
rect 497 1152 582 1157
rect 801 1152 862 1157
rect 897 1152 926 1157
rect 953 1152 1006 1157
rect 1121 1152 1206 1157
rect 1217 1152 1446 1157
rect 1457 1152 1990 1157
rect 2041 1152 2190 1157
rect 2201 1152 2246 1157
rect 2257 1152 2558 1157
rect 2617 1152 2662 1157
rect 2689 1152 2766 1157
rect 2785 1152 2870 1157
rect 2897 1152 2966 1157
rect 3129 1152 3190 1157
rect 3281 1152 3342 1157
rect 185 1142 350 1147
rect 385 1142 542 1147
rect 617 1142 694 1147
rect 185 1137 190 1142
rect 81 1132 126 1137
rect 161 1132 190 1137
rect 345 1137 350 1142
rect 345 1132 742 1137
rect 81 1107 86 1132
rect 897 1127 902 1152
rect 1001 1147 1126 1152
rect 1201 1147 1206 1152
rect 921 1142 982 1147
rect 1201 1142 1262 1147
rect 1457 1142 1462 1152
rect 2257 1147 2262 1152
rect 2785 1147 2790 1152
rect 1521 1142 1582 1147
rect 1609 1142 1654 1147
rect 1697 1142 1782 1147
rect 1873 1142 2110 1147
rect 2169 1142 2262 1147
rect 2273 1142 2382 1147
rect 2457 1142 2478 1147
rect 2489 1142 2790 1147
rect 2841 1142 2950 1147
rect 1281 1137 1462 1142
rect 2961 1137 2966 1152
rect 2977 1142 3182 1147
rect 3265 1142 3294 1147
rect 3265 1137 3270 1142
rect 1025 1132 1286 1137
rect 1537 1132 1566 1137
rect 1753 1132 1798 1137
rect 1825 1132 2894 1137
rect 2961 1132 3006 1137
rect 3225 1132 3270 1137
rect 3345 1132 3366 1137
rect 3345 1127 3350 1132
rect 185 1122 254 1127
rect 289 1122 334 1127
rect 417 1122 446 1127
rect 545 1122 574 1127
rect 625 1122 670 1127
rect 713 1122 806 1127
rect 873 1122 1070 1127
rect 1137 1122 1270 1127
rect 1329 1122 1606 1127
rect 1721 1122 1774 1127
rect 1881 1122 1990 1127
rect 2049 1122 2086 1127
rect 2097 1122 2470 1127
rect 2625 1122 2966 1127
rect 3281 1122 3350 1127
rect 3369 1122 3398 1127
rect 441 1117 550 1122
rect 801 1117 806 1122
rect 105 1112 142 1117
rect 169 1112 302 1117
rect 337 1112 398 1117
rect 593 1112 790 1117
rect 801 1112 854 1117
rect 929 1112 1022 1117
rect 1041 1112 1238 1117
rect 1265 1112 1270 1122
rect 2489 1117 2606 1122
rect 1377 1112 1414 1117
rect 1473 1112 1566 1117
rect 1705 1112 2494 1117
rect 2601 1112 2782 1117
rect 2825 1112 2902 1117
rect 3073 1112 3238 1117
rect 3249 1112 3294 1117
rect 3361 1112 3414 1117
rect 1585 1107 1686 1112
rect 81 1102 126 1107
rect 185 1102 246 1107
rect 289 1102 326 1107
rect 353 1102 414 1107
rect 465 1102 574 1107
rect 625 1102 774 1107
rect 889 1102 958 1107
rect 1017 1102 1398 1107
rect 1505 1102 1590 1107
rect 1681 1102 2038 1107
rect 2105 1102 2182 1107
rect 2193 1102 2278 1107
rect 2297 1102 2598 1107
rect 2649 1102 2710 1107
rect 2809 1102 2998 1107
rect 3153 1102 3318 1107
rect 465 1097 470 1102
rect 305 1092 334 1097
rect 329 1087 334 1092
rect 393 1092 470 1097
rect 569 1097 574 1102
rect 569 1092 1134 1097
rect 1153 1092 1246 1097
rect 393 1087 398 1092
rect 1393 1087 1398 1102
rect 2273 1097 2278 1102
rect 1473 1092 1494 1097
rect 1537 1092 1806 1097
rect 1833 1092 1910 1097
rect 1937 1092 2046 1097
rect 2065 1092 2198 1097
rect 2273 1092 2430 1097
rect 2441 1092 2542 1097
rect 2673 1092 2798 1097
rect 2953 1092 2982 1097
rect 3137 1092 3206 1097
rect 3257 1092 3278 1097
rect 3289 1092 3326 1097
rect 1937 1087 1942 1092
rect 2793 1087 2958 1092
rect 329 1082 398 1087
rect 481 1082 702 1087
rect 753 1082 894 1087
rect 929 1082 1318 1087
rect 1393 1082 1718 1087
rect 1753 1082 1942 1087
rect 1961 1082 2310 1087
rect 2625 1082 2646 1087
rect 2329 1077 2454 1082
rect 417 1072 502 1077
rect 545 1072 734 1077
rect 769 1072 910 1077
rect 1105 1072 1790 1077
rect 1817 1072 1870 1077
rect 1905 1072 1974 1077
rect 2041 1072 2334 1077
rect 2449 1072 2646 1077
rect 2689 1072 2798 1077
rect 2881 1072 3142 1077
rect 929 1067 1086 1072
rect 497 1062 534 1067
rect 601 1062 934 1067
rect 1081 1062 1270 1067
rect 1561 1062 1614 1067
rect 1625 1062 2062 1067
rect 2097 1062 2438 1067
rect 2793 1062 2950 1067
rect 1265 1057 1542 1062
rect 2457 1057 2774 1062
rect 505 1052 550 1057
rect 889 1052 1150 1057
rect 1537 1052 2462 1057
rect 2769 1052 2942 1057
rect 665 1047 870 1052
rect 377 1042 494 1047
rect 489 1037 494 1042
rect 561 1042 670 1047
rect 865 1042 1430 1047
rect 1441 1042 3006 1047
rect 3249 1042 3358 1047
rect 561 1037 566 1042
rect 489 1032 566 1037
rect 681 1032 750 1037
rect 793 1032 1078 1037
rect 1225 1032 1382 1037
rect 1393 1032 1550 1037
rect 1673 1032 2894 1037
rect 3169 1032 3214 1037
rect 3361 1032 3422 1037
rect 1073 1027 1230 1032
rect 1393 1027 1398 1032
rect 1545 1027 1678 1032
rect 233 1022 334 1027
rect 353 1022 374 1027
rect 625 1022 710 1027
rect 809 1022 934 1027
rect 969 1022 1054 1027
rect 1249 1022 1286 1027
rect 1361 1022 1422 1027
rect 1449 1022 1502 1027
rect 1697 1022 1790 1027
rect 1849 1022 1902 1027
rect 1953 1022 2142 1027
rect 2185 1022 2406 1027
rect 2433 1022 2478 1027
rect 2553 1022 2598 1027
rect 2641 1022 2686 1027
rect 3145 1022 3198 1027
rect 3345 1022 3382 1027
rect 233 1017 238 1022
rect 169 1012 238 1017
rect 329 1017 334 1022
rect 625 1017 630 1022
rect 929 1017 934 1022
rect 329 1012 510 1017
rect 593 1012 630 1017
rect 873 1012 918 1017
rect 929 1012 1414 1017
rect 1577 1012 1798 1017
rect 1817 1012 2038 1017
rect 2049 1012 2110 1017
rect 2201 1012 2222 1017
rect 2233 1012 2614 1017
rect 2705 1012 2734 1017
rect 2801 1012 2982 1017
rect 3297 1012 3382 1017
rect 729 1007 822 1012
rect 2033 1007 2038 1012
rect 705 1002 734 1007
rect 817 1002 1102 1007
rect 1153 1002 1350 1007
rect 1361 1002 1390 1007
rect 1481 1002 1558 1007
rect 1705 1002 1838 1007
rect 1849 1002 1870 1007
rect 2033 1002 2254 1007
rect 2297 1002 2454 1007
rect 273 997 382 1002
rect 1345 997 1350 1002
rect 1889 997 1998 1002
rect 249 992 278 997
rect 377 992 446 997
rect 465 992 678 997
rect 753 992 806 997
rect 913 992 1102 997
rect 1161 992 1326 997
rect 1345 992 1454 997
rect 1465 992 1894 997
rect 1993 992 2670 997
rect 465 987 470 992
rect 113 982 470 987
rect 449 972 654 977
rect 305 967 430 972
rect 673 967 678 992
rect 689 982 950 987
rect 1145 982 1318 987
rect 1377 982 1606 987
rect 969 977 1094 982
rect 1601 977 1606 982
rect 1713 982 1982 987
rect 2057 982 2302 987
rect 2313 982 2494 987
rect 1713 977 1718 982
rect 2705 977 2710 1012
rect 3097 992 3198 997
rect 3257 992 3358 997
rect 2721 982 2758 987
rect 3057 982 3110 987
rect 3257 982 3366 987
rect 753 972 782 977
rect 913 972 974 977
rect 1089 972 1206 977
rect 1289 972 1582 977
rect 1601 972 1718 977
rect 1737 972 2006 977
rect 2057 972 2110 977
rect 2129 972 2294 977
rect 2369 972 2662 977
rect 2705 972 2734 977
rect 2777 972 3022 977
rect 3321 972 3342 977
rect 753 967 758 972
rect 1201 967 1294 972
rect 2777 967 2782 972
rect 3073 967 3166 972
rect 281 962 310 967
rect 425 962 462 967
rect 673 962 758 967
rect 881 962 966 967
rect 1001 962 1094 967
rect 1145 962 1182 967
rect 1313 962 1446 967
rect 1497 962 1542 967
rect 1769 962 1886 967
rect 1945 962 1998 967
rect 2009 962 2054 967
rect 2073 962 2206 967
rect 2265 962 2334 967
rect 2369 962 2782 967
rect 3009 962 3078 967
rect 3161 962 3190 967
rect 497 957 598 962
rect 97 952 118 957
rect 209 952 238 957
rect 249 952 286 957
rect 297 952 358 957
rect 385 952 502 957
rect 593 952 622 957
rect 777 952 854 957
rect 865 952 894 957
rect 1113 952 1198 957
rect 1209 952 1286 957
rect 1441 952 1622 957
rect 1633 952 1790 957
rect 1809 952 2294 957
rect 2401 952 2822 957
rect 2961 952 2990 957
rect 3089 952 3190 957
rect 113 942 278 947
rect 289 942 526 947
rect 585 942 806 947
rect 825 942 918 947
rect 937 942 1054 947
rect 1073 942 1182 947
rect 1329 942 1694 947
rect 1721 942 1766 947
rect 1913 942 2046 947
rect 2065 942 2238 947
rect 2265 942 2326 947
rect 913 937 918 942
rect 1761 937 1886 942
rect 193 932 262 937
rect 353 932 390 937
rect 457 932 486 937
rect 665 932 814 937
rect 825 932 862 937
rect 913 932 1190 937
rect 1201 932 1446 937
rect 1457 932 1742 937
rect 1881 932 2006 937
rect 2177 932 2286 937
rect 2345 932 2390 937
rect 257 927 262 932
rect 481 927 566 932
rect 1185 927 1190 932
rect 1441 927 1446 932
rect 2025 927 2158 932
rect 2401 927 2406 952
rect 2433 942 2478 947
rect 2489 942 2590 947
rect 2673 942 2702 947
rect 2801 942 2934 947
rect 2697 937 2806 942
rect 2497 932 2582 937
rect 2881 932 2942 937
rect 3321 932 3398 937
rect 257 922 382 927
rect 561 922 902 927
rect 1057 922 1094 927
rect 1185 922 1246 927
rect 1353 922 1430 927
rect 1441 922 1710 927
rect 1785 922 2030 927
rect 2153 922 2406 927
rect 1241 917 1358 922
rect 1425 917 1430 922
rect 2577 917 2582 932
rect 2593 922 2630 927
rect 2761 922 2830 927
rect 2849 922 3030 927
rect 3313 922 3414 927
rect 2761 917 2766 922
rect 353 912 430 917
rect 809 912 1006 917
rect 1153 912 1222 917
rect 1425 912 1910 917
rect 1961 912 2062 917
rect 2089 912 2142 917
rect 2209 912 2326 917
rect 2353 912 2374 917
rect 2425 912 2558 917
rect 2577 912 2614 917
rect 2649 912 2718 917
rect 2737 912 2766 917
rect 2825 917 2830 922
rect 2825 912 2910 917
rect 2961 912 3062 917
rect 3105 912 3246 917
rect 3321 912 3350 917
rect 561 907 686 912
rect 2425 907 2430 912
rect 457 902 566 907
rect 681 902 710 907
rect 833 902 894 907
rect 953 902 1326 907
rect 1385 902 1462 907
rect 1473 902 1518 907
rect 1609 902 1862 907
rect 1937 902 2430 907
rect 2553 907 2558 912
rect 2553 902 2918 907
rect 1473 897 1478 902
rect 1857 897 1862 902
rect 337 892 358 897
rect 577 892 862 897
rect 1161 892 1398 897
rect 1457 892 1478 897
rect 1497 892 1542 897
rect 1713 892 1838 897
rect 1857 892 2198 897
rect 2209 892 2262 897
rect 2329 892 2462 897
rect 2497 892 2566 897
rect 2617 892 2750 897
rect 2825 892 3030 897
rect 401 887 494 892
rect 1049 887 1142 892
rect 1561 887 1694 892
rect 3025 887 3030 892
rect 3113 892 3142 897
rect 3113 887 3118 892
rect 377 882 406 887
rect 489 882 950 887
rect 1025 882 1054 887
rect 1137 882 1222 887
rect 1401 882 1566 887
rect 1689 882 2838 887
rect 3025 882 3118 887
rect 1241 877 1382 882
rect 305 872 478 877
rect 473 867 478 872
rect 593 872 862 877
rect 961 872 1246 877
rect 1377 872 2222 877
rect 2369 872 2710 877
rect 593 867 598 872
rect 857 867 966 872
rect 2705 867 2710 872
rect 2977 872 3006 877
rect 2977 867 2982 872
rect 233 862 454 867
rect 473 862 598 867
rect 617 862 838 867
rect 1065 862 1446 867
rect 1465 862 1534 867
rect 1641 862 1758 867
rect 1809 862 1902 867
rect 2041 862 2118 867
rect 2129 862 2174 867
rect 2193 862 2310 867
rect 2329 862 2670 867
rect 2705 862 2982 867
rect 1921 857 2022 862
rect 2305 857 2310 862
rect 217 852 270 857
rect 321 852 430 857
rect 625 852 854 857
rect 953 852 1190 857
rect 1217 852 1478 857
rect 1561 852 1614 857
rect 1641 852 1926 857
rect 2017 852 2286 857
rect 2305 852 2518 857
rect 2545 852 2566 857
rect 2585 852 2686 857
rect 625 847 630 852
rect 97 842 630 847
rect 649 842 846 847
rect 865 842 942 847
rect 1001 842 1414 847
rect 1521 842 1670 847
rect 1849 842 1918 847
rect 1969 842 2166 847
rect 2249 842 2542 847
rect 97 817 102 842
rect 113 832 206 837
rect 329 832 374 837
rect 593 832 686 837
rect 705 832 798 837
rect 817 832 862 837
rect 897 832 1078 837
rect 1113 832 1198 837
rect 1297 832 1486 837
rect 1521 827 1526 842
rect 1689 837 1830 842
rect 2161 837 2254 842
rect 1537 832 1694 837
rect 1825 832 1870 837
rect 2025 832 2142 837
rect 2273 832 2438 837
rect 2457 832 2630 837
rect 2873 832 3110 837
rect 3353 832 3406 837
rect 1889 827 2030 832
rect 193 822 446 827
rect 457 822 518 827
rect 561 822 598 827
rect 657 822 1222 827
rect 1241 822 1270 827
rect 1313 822 1406 827
rect 1417 822 1526 827
rect 1537 822 1590 827
rect 1657 822 1894 827
rect 2049 822 2310 827
rect 2385 822 2646 827
rect 3201 822 3230 827
rect 3297 822 3414 827
rect 1265 817 1270 822
rect 97 812 118 817
rect 529 812 1270 817
rect 1377 817 1382 822
rect 1537 817 1542 822
rect 2305 817 2310 822
rect 1377 812 1542 817
rect 1609 812 2030 817
rect 2081 812 2174 817
rect 2305 812 2574 817
rect 2769 812 2854 817
rect 3385 812 3504 817
rect 337 807 470 812
rect 529 807 534 812
rect 2593 807 2686 812
rect 2769 807 2774 812
rect 185 802 206 807
rect 273 802 342 807
rect 465 802 534 807
rect 545 802 582 807
rect 657 802 774 807
rect 817 802 990 807
rect 1049 802 1318 807
rect 1401 802 1678 807
rect 1897 802 1934 807
rect 2049 802 2182 807
rect 2297 802 2438 807
rect 2497 802 2598 807
rect 2681 802 2774 807
rect 2849 807 2854 812
rect 2849 802 3006 807
rect 177 792 222 797
rect 257 792 310 797
rect 337 792 454 797
rect 561 792 670 797
rect 817 787 822 802
rect 1761 797 1878 802
rect 833 792 1270 797
rect 1289 792 1598 797
rect 1689 792 1766 797
rect 1873 792 2670 797
rect 3297 792 3374 797
rect 1593 787 1694 792
rect 2809 787 2886 792
rect 3297 787 3302 792
rect 3369 787 3374 792
rect 3473 792 3504 797
rect 3473 787 3478 792
rect 105 782 262 787
rect 353 782 470 787
rect 633 782 822 787
rect 937 782 1134 787
rect 1217 782 1574 787
rect 1777 782 2310 787
rect 2457 782 2494 787
rect 2553 782 2646 787
rect 2785 782 2814 787
rect 2881 782 3046 787
rect 3257 782 3302 787
rect 3313 782 3342 787
rect 3369 782 3478 787
rect 1129 777 1222 782
rect 2329 777 2438 782
rect 225 772 310 777
rect 329 772 526 777
rect 577 772 598 777
rect 665 772 1110 777
rect 1241 772 1302 777
rect 1313 772 1366 777
rect 1401 772 1486 777
rect 1569 772 1638 777
rect 1897 772 1934 777
rect 2113 772 2190 777
rect 2305 772 2334 777
rect 2433 772 2590 777
rect 2841 772 2870 777
rect 1721 767 1878 772
rect 1929 767 2118 772
rect 2185 767 2310 772
rect 2865 767 2870 772
rect 2985 772 3014 777
rect 2985 767 2990 772
rect 393 762 534 767
rect 609 762 710 767
rect 729 762 814 767
rect 841 762 1038 767
rect 1089 762 1182 767
rect 1257 762 1558 767
rect 1697 762 1726 767
rect 1873 762 1910 767
rect 2137 762 2166 767
rect 2329 762 2406 767
rect 2425 762 2534 767
rect 2569 762 2742 767
rect 2865 762 2990 767
rect 2737 757 2742 762
rect 49 752 118 757
rect 409 752 486 757
rect 625 752 854 757
rect 1233 752 1406 757
rect 1441 752 2038 757
rect 2241 752 2310 757
rect 2409 752 2654 757
rect 2737 752 2766 757
rect 49 737 54 752
rect 313 747 390 752
rect 2241 747 2246 752
rect 65 742 110 747
rect 225 742 318 747
rect 385 742 526 747
rect 617 742 686 747
rect 801 742 830 747
rect 897 742 926 747
rect 1137 742 1174 747
rect 1201 742 1278 747
rect 1361 742 1590 747
rect 1737 742 1822 747
rect 1849 742 1950 747
rect 2217 742 2246 747
rect 2305 747 2310 752
rect 2305 742 2422 747
rect 2473 742 2494 747
rect 2545 742 2574 747
rect 2665 742 2726 747
rect 3113 742 3166 747
rect 3201 742 3270 747
rect 1169 737 1174 742
rect 49 732 70 737
rect 329 732 470 737
rect 497 732 566 737
rect 633 727 638 737
rect 713 732 958 737
rect 977 732 1062 737
rect 1121 732 1158 737
rect 1169 732 1838 737
rect 1881 732 2070 737
rect 2089 732 2254 737
rect 2281 732 2382 737
rect 977 727 982 732
rect 97 722 118 727
rect 185 722 214 727
rect 249 722 494 727
rect 633 722 686 727
rect 785 722 830 727
rect 865 722 982 727
rect 1057 727 1062 732
rect 2401 727 2510 732
rect 1057 722 1614 727
rect 1649 722 2006 727
rect 2169 722 2406 727
rect 2505 722 2534 727
rect 2545 722 2550 742
rect 2569 737 2670 742
rect 3201 737 3206 742
rect 3177 732 3206 737
rect 3265 737 3270 742
rect 3265 732 3366 737
rect 2657 722 2694 727
rect 2049 717 2150 722
rect 161 712 246 717
rect 289 712 326 717
rect 401 712 654 717
rect 985 712 1046 717
rect 1137 712 1166 717
rect 1289 712 2054 717
rect 2145 712 2750 717
rect 2825 712 2950 717
rect 2969 712 3070 717
rect 3169 712 3254 717
rect 177 702 230 707
rect 241 702 246 712
rect 305 702 342 707
rect 377 702 526 707
rect 617 702 646 707
rect 729 702 774 707
rect 793 702 966 707
rect 1145 702 1174 707
rect 1241 702 1286 707
rect 1297 702 1878 707
rect 2065 702 2454 707
rect 2529 702 2742 707
rect 3089 702 3206 707
rect 3281 702 3342 707
rect 225 697 230 702
rect 337 697 342 702
rect 521 697 622 702
rect 793 697 798 702
rect 961 697 1126 702
rect 1873 697 2070 702
rect 225 692 254 697
rect 337 692 374 697
rect 481 692 502 697
rect 721 692 798 697
rect 1121 692 1238 697
rect 1273 692 1366 697
rect 1409 692 1494 697
rect 1545 692 1598 697
rect 1641 692 1750 697
rect 1817 692 1854 697
rect 2089 692 2182 697
rect 2201 692 2718 697
rect 3121 692 3222 697
rect 3217 687 3222 692
rect 3321 692 3350 697
rect 3321 687 3326 692
rect 409 682 614 687
rect 649 682 750 687
rect 761 682 1246 687
rect 1281 682 1470 687
rect 1625 682 1726 687
rect 1769 682 1798 687
rect 1817 682 1958 687
rect 1993 682 2110 687
rect 2153 682 2422 687
rect 2657 682 2766 687
rect 3217 682 3326 687
rect 545 672 838 677
rect 1001 672 1054 677
rect 1089 672 1302 677
rect 1393 672 1614 677
rect 1697 672 1846 677
rect 2097 672 2486 677
rect 833 667 1006 672
rect 1297 667 1398 672
rect 1609 667 1702 672
rect 1841 667 2102 672
rect 657 662 814 667
rect 1153 662 1198 667
rect 1209 662 1278 667
rect 1417 662 1478 667
rect 1721 662 1822 667
rect 2121 662 2198 667
rect 2209 662 2246 667
rect 2329 662 2494 667
rect 3017 662 3198 667
rect 1025 657 1134 662
rect 345 652 486 657
rect 505 652 638 657
rect 697 652 1030 657
rect 1129 652 2446 657
rect 2505 652 2574 657
rect 505 647 510 652
rect 433 642 510 647
rect 633 647 638 652
rect 2441 647 2510 652
rect 3017 647 3022 662
rect 633 642 854 647
rect 1041 642 1182 647
rect 1329 642 1406 647
rect 1449 642 1478 647
rect 921 637 1022 642
rect 1201 637 1278 642
rect 1329 637 1334 642
rect 1601 637 1606 647
rect 1705 642 1854 647
rect 2105 642 2374 647
rect 2385 642 2422 647
rect 2601 642 2678 647
rect 2801 642 3022 647
rect 3193 647 3198 662
rect 3193 642 3222 647
rect 2385 637 2390 642
rect 97 632 198 637
rect 329 632 726 637
rect 809 632 862 637
rect 897 632 926 637
rect 1017 632 1110 637
rect 1129 632 1206 637
rect 1273 632 1334 637
rect 1353 632 1390 637
rect 1601 632 2390 637
rect 2489 632 2550 637
rect 2577 632 2646 637
rect 3033 632 3190 637
rect 3313 632 3406 637
rect 3313 627 3318 632
rect 65 622 110 627
rect 289 622 350 627
rect 489 622 518 627
rect 617 622 798 627
rect 889 622 1014 627
rect 1193 622 1262 627
rect 1409 622 1462 627
rect 1521 622 1614 627
rect 1625 622 1678 627
rect 1745 622 1910 627
rect 2209 622 2310 627
rect 2457 622 2542 627
rect 3137 622 3318 627
rect 3361 622 3414 627
rect 513 617 622 622
rect 793 617 894 622
rect 3137 617 3142 622
rect 209 612 318 617
rect 337 612 470 617
rect 641 612 750 617
rect 913 612 1286 617
rect 1305 612 1662 617
rect 1793 612 1902 617
rect 2273 612 2446 617
rect 2505 612 2534 617
rect 2593 612 2630 617
rect 2937 612 3142 617
rect 3153 612 3198 617
rect 961 607 966 612
rect 2169 607 2254 612
rect 2289 607 2294 612
rect 2441 607 2510 612
rect 3297 607 3302 617
rect 513 602 558 607
rect 689 597 694 607
rect 857 602 918 607
rect 961 602 990 607
rect 1257 602 1334 607
rect 1393 602 1510 607
rect 1521 602 1638 607
rect 1745 602 1782 607
rect 1145 597 1238 602
rect 1393 597 1398 602
rect 281 592 382 597
rect 393 592 446 597
rect 513 592 542 597
rect 593 592 982 597
rect 1041 592 1150 597
rect 1233 592 1398 597
rect 1505 597 1510 602
rect 1745 597 1750 602
rect 1505 592 1750 597
rect 1777 597 1782 602
rect 1849 602 2038 607
rect 2049 602 2174 607
rect 2249 602 2294 607
rect 2929 602 3350 607
rect 1849 597 1854 602
rect 2033 597 2038 602
rect 1777 592 1854 597
rect 1873 592 1942 597
rect 2033 592 2086 597
rect 2185 592 2222 597
rect 2241 592 2302 597
rect 2321 592 2478 597
rect 2705 592 2766 597
rect 3073 592 3190 597
rect 3345 592 3350 602
rect 2081 587 2166 592
rect 2321 587 2326 592
rect 473 582 534 587
rect 577 582 726 587
rect 817 582 1030 587
rect 1161 582 1574 587
rect 1929 582 2070 587
rect 2161 582 2190 587
rect 2265 582 2326 587
rect 2473 587 2478 592
rect 2473 582 2502 587
rect 2689 582 2774 587
rect 2905 582 3014 587
rect 3057 582 3222 587
rect 1049 577 1142 582
rect 1569 577 1574 582
rect 289 572 326 577
rect 353 572 406 577
rect 545 572 1054 577
rect 1137 572 1502 577
rect 1529 572 1550 577
rect 1569 572 1758 577
rect 1777 572 1846 577
rect 1921 572 1998 577
rect 2065 572 2462 577
rect 2569 572 2638 577
rect 1753 567 1758 572
rect 2569 567 2574 572
rect 265 562 342 567
rect 337 557 342 562
rect 417 562 542 567
rect 561 562 702 567
rect 849 562 1046 567
rect 1081 562 1350 567
rect 1361 562 1494 567
rect 1753 562 2334 567
rect 2385 562 2406 567
rect 2545 562 2574 567
rect 2633 567 2638 572
rect 3097 567 3238 572
rect 2633 562 2662 567
rect 2865 562 3054 567
rect 3073 562 3102 567
rect 3233 562 3438 567
rect 417 557 422 562
rect 1345 557 1350 562
rect 1513 557 1598 562
rect 2865 557 2870 562
rect 201 552 246 557
rect 337 552 422 557
rect 569 552 1022 557
rect 1145 552 1214 557
rect 1345 552 1518 557
rect 1593 552 2686 557
rect 2705 552 2870 557
rect 3049 557 3054 562
rect 3049 552 3222 557
rect 1017 547 1150 552
rect 1233 547 1326 552
rect 249 542 310 547
rect 545 542 902 547
rect 961 542 998 547
rect 1169 542 1238 547
rect 1321 542 1422 547
rect 1457 542 1582 547
rect 1817 542 2006 547
rect 2129 542 2334 547
rect 2353 542 2486 547
rect 2529 542 2606 547
rect 2353 537 2358 542
rect 2705 537 2710 552
rect 3249 547 3358 552
rect 2865 542 3254 547
rect 3353 542 3422 547
rect 249 532 286 537
rect 425 532 518 537
rect 681 532 758 537
rect 769 532 1046 537
rect 1065 532 1142 537
rect 1217 532 1358 537
rect 1369 532 1398 537
rect 1441 532 1566 537
rect 1697 532 2166 537
rect 2185 532 2358 537
rect 2449 532 2574 537
rect 2617 532 2710 537
rect 3121 532 3246 537
rect 3265 532 3326 537
rect 3361 532 3406 537
rect 537 527 662 532
rect 769 527 774 532
rect 1041 527 1046 532
rect 1585 527 1678 532
rect 2369 527 2454 532
rect 217 522 270 527
rect 393 522 542 527
rect 657 522 774 527
rect 841 522 1014 527
rect 1041 522 1590 527
rect 1673 522 2086 527
rect 2185 522 2206 527
rect 2289 522 2374 527
rect 2593 522 2654 527
rect 2777 522 2838 527
rect 2473 517 2598 522
rect 2833 517 2838 522
rect 2969 522 3174 527
rect 3233 522 3278 527
rect 2969 517 2974 522
rect 3169 517 3174 522
rect 177 512 230 517
rect 297 512 638 517
rect 649 512 686 517
rect 697 512 1110 517
rect 1153 512 1214 517
rect 1393 512 1622 517
rect 1649 512 1686 517
rect 1729 512 1862 517
rect 1929 512 1974 517
rect 2025 512 2110 517
rect 2153 512 2278 517
rect 2305 512 2430 517
rect 2449 512 2478 517
rect 2665 512 2726 517
rect 2833 512 2974 517
rect 3017 512 3142 517
rect 3169 512 3190 517
rect 225 507 230 512
rect 1233 507 1374 512
rect 1857 507 1862 512
rect 3185 507 3190 512
rect 3289 512 3342 517
rect 3289 507 3294 512
rect 225 502 374 507
rect 513 502 558 507
rect 697 502 1238 507
rect 1369 502 1662 507
rect 1801 502 1838 507
rect 1857 502 1974 507
rect 1985 502 2062 507
rect 2185 502 2214 507
rect 2257 502 2302 507
rect 2409 502 2438 507
rect 2489 502 2534 507
rect 2753 502 2814 507
rect 3033 502 3102 507
rect 3185 502 3294 507
rect 3329 502 3382 507
rect 369 497 518 502
rect 593 497 702 502
rect 1681 497 1774 502
rect 153 492 350 497
rect 537 492 598 497
rect 721 492 1166 497
rect 1217 492 1406 497
rect 1625 492 1686 497
rect 1769 492 1798 497
rect 1809 492 2318 497
rect 2441 492 2606 497
rect 3313 492 3422 497
rect 1425 487 1606 492
rect 137 482 166 487
rect 161 467 166 482
rect 289 482 414 487
rect 481 482 686 487
rect 753 482 854 487
rect 865 482 1430 487
rect 1601 482 1902 487
rect 2009 482 2054 487
rect 2233 482 2462 487
rect 2489 482 2518 487
rect 2625 482 2710 487
rect 3129 482 3262 487
rect 289 467 294 482
rect 865 477 870 482
rect 2625 477 2630 482
rect 313 472 366 477
rect 601 472 870 477
rect 905 472 982 477
rect 1105 472 1334 477
rect 1425 472 1478 477
rect 1497 472 1646 477
rect 1657 472 1734 477
rect 1769 472 1814 477
rect 1889 472 2150 477
rect 2257 472 2630 477
rect 2705 477 2710 482
rect 2705 472 2734 477
rect 2753 472 2918 477
rect 505 467 582 472
rect 1329 467 1430 472
rect 1473 467 1478 472
rect 2753 467 2758 472
rect 161 462 294 467
rect 361 462 510 467
rect 577 462 830 467
rect 857 462 934 467
rect 961 462 1310 467
rect 1473 462 1774 467
rect 1785 462 1894 467
rect 2281 462 2542 467
rect 2729 462 2758 467
rect 2913 467 2918 472
rect 2913 462 2942 467
rect 1937 457 2262 462
rect 2537 457 2542 462
rect 2641 457 2734 462
rect 521 452 758 457
rect 929 452 974 457
rect 1049 452 1302 457
rect 1377 452 1590 457
rect 1601 452 1862 457
rect 1913 452 1942 457
rect 2257 452 2510 457
rect 2537 452 2646 457
rect 2777 452 2894 457
rect 753 447 934 452
rect 2777 447 2782 452
rect 281 442 614 447
rect 657 442 734 447
rect 953 442 974 447
rect 1113 442 2518 447
rect 2673 442 2782 447
rect 2889 447 2894 452
rect 2889 442 3022 447
rect 281 437 286 442
rect 161 432 286 437
rect 409 432 486 437
rect 593 432 742 437
rect 817 432 894 437
rect 993 432 1198 437
rect 1281 432 1446 437
rect 1521 432 1926 437
rect 1945 432 2038 437
rect 2049 432 2158 437
rect 2185 432 2246 437
rect 2281 432 2654 437
rect 2713 432 2742 437
rect 737 427 742 432
rect 1521 427 1526 432
rect 1921 427 1926 432
rect 2737 427 2742 432
rect 2801 432 2878 437
rect 2801 427 2806 432
rect 2921 427 3054 432
rect 97 422 214 427
rect 209 417 214 422
rect 289 422 606 427
rect 737 422 854 427
rect 953 422 1030 427
rect 1145 422 1270 427
rect 1337 422 1526 427
rect 1593 422 1806 427
rect 1857 422 1886 427
rect 1921 422 2126 427
rect 2377 422 2494 427
rect 2737 422 2806 427
rect 2897 422 2926 427
rect 3049 422 3078 427
rect 3161 422 3222 427
rect 289 417 294 422
rect 625 417 718 422
rect 1025 417 1126 422
rect 1265 417 1342 422
rect 105 412 142 417
rect 209 412 294 417
rect 313 412 630 417
rect 713 412 998 417
rect 1121 412 1190 417
rect 1361 412 1934 417
rect 2201 412 2310 417
rect 993 407 998 412
rect 1953 407 2182 412
rect 2329 407 2518 412
rect 129 402 166 407
rect 409 402 438 407
rect 585 402 982 407
rect 993 402 1230 407
rect 1249 402 1342 407
rect 1401 402 1958 407
rect 2177 402 2334 407
rect 2513 402 2542 407
rect 433 397 590 402
rect 2593 397 2598 417
rect 2825 412 2878 417
rect 2889 412 3030 417
rect 3065 412 3190 417
rect 3209 412 3310 417
rect 3385 402 3438 407
rect 609 392 1142 397
rect 1153 392 1318 397
rect 1393 392 1630 397
rect 1873 392 2686 397
rect 2745 392 2814 397
rect 1625 387 1878 392
rect 2809 387 2814 392
rect 2929 392 2982 397
rect 2929 387 2934 392
rect 73 382 230 387
rect 497 382 694 387
rect 881 382 990 387
rect 1009 382 1246 387
rect 1297 382 1502 387
rect 1569 382 1606 387
rect 1897 382 2054 387
rect 2129 382 2198 387
rect 2345 382 2478 387
rect 2497 382 2526 387
rect 2217 377 2318 382
rect 2521 377 2526 382
rect 2601 382 2630 387
rect 2657 382 2742 387
rect 2809 382 2934 387
rect 2601 377 2606 382
rect 249 372 366 377
rect 385 372 494 377
rect 585 372 710 377
rect 841 372 1134 377
rect 1257 372 1590 377
rect 1601 372 1710 377
rect 1801 372 2110 377
rect 2145 372 2222 377
rect 2313 372 2342 377
rect 249 367 254 372
rect 129 362 254 367
rect 361 367 366 372
rect 2337 367 2342 372
rect 2417 372 2446 377
rect 2521 372 2606 377
rect 2977 377 2982 392
rect 3089 392 3142 397
rect 3089 377 3094 392
rect 3137 387 3142 392
rect 3209 392 3430 397
rect 3209 387 3214 392
rect 3137 382 3214 387
rect 2977 372 3094 377
rect 2417 367 2422 372
rect 361 362 702 367
rect 769 362 830 367
rect 1009 362 1486 367
rect 1497 362 1542 367
rect 1721 362 1846 367
rect 2097 362 2318 367
rect 2337 362 2422 367
rect 857 357 990 362
rect 1841 357 2102 362
rect 241 352 790 357
rect 801 352 862 357
rect 985 352 1158 357
rect 1169 352 1246 357
rect 1265 352 1398 357
rect 1409 352 1622 357
rect 2121 352 2166 357
rect 2209 352 2262 357
rect 2689 352 2782 357
rect 2809 352 3342 357
rect 801 347 806 352
rect 1153 347 1158 352
rect 1393 347 1398 352
rect 1641 347 1822 352
rect 297 342 454 347
rect 473 342 542 347
rect 673 342 806 347
rect 817 342 958 347
rect 1001 342 1102 347
rect 1153 342 1382 347
rect 1393 342 1646 347
rect 1817 342 1846 347
rect 1865 342 1974 347
rect 1993 342 2110 347
rect 561 337 654 342
rect 1377 337 1382 342
rect 1865 337 1870 342
rect 193 332 278 337
rect 361 332 414 337
rect 433 332 566 337
rect 649 332 1166 337
rect 1217 327 1222 337
rect 1265 332 1286 337
rect 1329 327 1334 337
rect 1377 332 1430 337
rect 1481 332 1870 337
rect 1969 337 1974 342
rect 1969 332 1998 337
rect 2105 332 2134 337
rect 2409 332 2558 337
rect 2577 332 2646 337
rect 1993 327 2110 332
rect 2577 327 2582 332
rect 289 322 390 327
rect 409 322 478 327
rect 513 322 1334 327
rect 1417 322 1502 327
rect 1721 322 1974 327
rect 2513 322 2582 327
rect 2641 327 2646 332
rect 2641 322 2670 327
rect 2785 322 3134 327
rect 385 317 390 322
rect 513 317 518 322
rect 1521 317 1702 322
rect 105 312 334 317
rect 385 312 486 317
rect 497 312 518 317
rect 529 312 654 317
rect 665 312 870 317
rect 865 307 870 312
rect 1017 312 1406 317
rect 1505 312 1526 317
rect 1697 312 2094 317
rect 2137 312 2246 317
rect 2537 312 2574 317
rect 1017 307 1022 312
rect 1401 307 1510 312
rect 2785 307 2790 322
rect 3129 317 3134 322
rect 3129 312 3158 317
rect 225 302 254 307
rect 481 302 718 307
rect 249 297 486 302
rect 713 297 718 302
rect 817 302 846 307
rect 865 302 1022 307
rect 1081 302 1214 307
rect 1249 302 1358 307
rect 1529 302 2222 307
rect 2577 302 2790 307
rect 2809 302 2918 307
rect 817 297 822 302
rect 1249 297 1254 302
rect 2809 297 2814 302
rect 505 292 598 297
rect 713 292 822 297
rect 1041 292 1134 297
rect 1145 292 1254 297
rect 1257 292 1422 297
rect 1593 292 1702 297
rect 2017 292 2502 297
rect 2625 292 2654 297
rect 1257 287 1262 292
rect 1441 287 1574 292
rect 1697 287 2022 292
rect 2649 287 2654 292
rect 2721 292 2814 297
rect 2721 287 2726 292
rect 273 282 518 287
rect 1161 282 1262 287
rect 1273 282 1446 287
rect 1569 282 1678 287
rect 2041 282 2174 287
rect 2649 282 2726 287
rect 2785 282 2894 287
rect 2913 277 2918 302
rect 3169 292 3222 297
rect 3169 277 3174 292
rect 529 272 798 277
rect 1017 272 1526 277
rect 1569 272 1614 277
rect 1801 272 2022 277
rect 2065 272 2110 277
rect 2913 272 3174 277
rect 465 267 534 272
rect 1801 267 1806 272
rect 2129 267 2254 272
rect 257 262 470 267
rect 769 262 942 267
rect 1137 262 1542 267
rect 1553 262 1806 267
rect 1889 262 2134 267
rect 2249 262 2430 267
rect 369 252 398 257
rect 393 247 398 252
rect 481 252 582 257
rect 793 252 1014 257
rect 1049 252 1086 257
rect 481 247 486 252
rect 1137 247 1142 262
rect 1537 257 1542 262
rect 1161 252 1334 257
rect 1537 252 2238 257
rect 2385 252 2414 257
rect 1353 247 1478 252
rect 2385 247 2390 252
rect 393 242 486 247
rect 601 242 750 247
rect 849 242 1142 247
rect 1281 242 1358 247
rect 1473 242 1502 247
rect 1537 242 1846 247
rect 1881 242 2174 247
rect 2249 242 2390 247
rect 2409 242 2446 247
rect 601 237 606 242
rect 745 237 830 242
rect 1161 237 1262 242
rect 2169 237 2254 242
rect 249 232 358 237
rect 561 232 606 237
rect 825 232 1166 237
rect 1257 232 2150 237
rect 2401 232 2510 237
rect 3089 232 3182 237
rect 377 222 542 227
rect 561 222 598 227
rect 681 222 822 227
rect 865 222 926 227
rect 1033 222 1534 227
rect 1625 222 1742 227
rect 1761 222 1950 227
rect 2057 222 2166 227
rect 2209 222 2318 227
rect 2545 222 2758 227
rect 2769 222 2862 227
rect 2929 222 3030 227
rect 377 217 382 222
rect 185 212 318 217
rect 345 212 382 217
rect 537 217 542 222
rect 921 217 1038 222
rect 2209 217 2214 222
rect 537 212 902 217
rect 1249 212 1406 217
rect 1417 212 1846 217
rect 2001 212 2030 217
rect 2057 212 2214 217
rect 2313 217 2318 222
rect 2753 217 2758 222
rect 2313 212 2350 217
rect 2753 212 2782 217
rect 2865 212 3358 217
rect 2777 207 2870 212
rect 89 202 398 207
rect 433 202 646 207
rect 665 202 1334 207
rect 1345 202 1886 207
rect 2041 202 2134 207
rect 2225 202 2302 207
rect 2481 202 2534 207
rect 2129 197 2134 202
rect 2529 197 2534 202
rect 2649 202 2678 207
rect 2889 202 2950 207
rect 3041 202 3070 207
rect 3321 202 3438 207
rect 2649 197 2654 202
rect 2945 197 3046 202
rect 169 192 198 197
rect 193 187 198 192
rect 305 192 462 197
rect 569 192 710 197
rect 745 192 1006 197
rect 1209 192 1246 197
rect 1257 192 1486 197
rect 1593 192 1702 197
rect 1793 192 1918 197
rect 1929 192 2118 197
rect 2129 192 2262 197
rect 2345 192 2478 197
rect 2529 192 2654 197
rect 2721 192 2926 197
rect 3193 192 3222 197
rect 305 187 310 192
rect 3217 187 3222 192
rect 3305 192 3334 197
rect 3305 187 3310 192
rect 193 182 310 187
rect 361 182 390 187
rect 473 182 590 187
rect 665 182 758 187
rect 969 182 1022 187
rect 1081 182 2078 187
rect 2209 182 2286 187
rect 2737 182 2766 187
rect 385 177 478 182
rect 753 177 758 182
rect 849 177 974 182
rect 2073 177 2214 182
rect 2761 177 2766 182
rect 2833 182 2926 187
rect 2953 182 3102 187
rect 3217 182 3310 187
rect 2833 177 2838 182
rect 753 172 854 177
rect 993 172 1182 177
rect 1193 172 1374 177
rect 1441 172 1582 177
rect 1849 172 1878 177
rect 2025 172 2054 177
rect 2233 172 2406 177
rect 2761 172 2838 177
rect 1873 167 1966 172
rect 2025 167 2030 172
rect 329 162 430 167
rect 497 162 534 167
rect 553 162 702 167
rect 873 162 974 167
rect 1185 162 1246 167
rect 1345 162 1846 167
rect 1961 162 2030 167
rect 2145 162 2254 167
rect 529 157 534 162
rect 993 157 1102 162
rect 209 152 310 157
rect 529 152 566 157
rect 721 152 790 157
rect 929 152 998 157
rect 1097 152 1126 157
rect 1225 152 1302 157
rect 1489 152 1574 157
rect 1809 152 1942 157
rect 2273 152 2478 157
rect 2857 152 3022 157
rect 209 147 214 152
rect 305 147 486 152
rect 721 147 726 152
rect 1641 147 1790 152
rect 2273 147 2278 152
rect 2857 147 2862 152
rect 65 142 214 147
rect 481 142 726 147
rect 737 142 1462 147
rect 1537 142 1646 147
rect 1785 142 1998 147
rect 2089 142 2278 147
rect 2385 142 2470 147
rect 2721 142 2862 147
rect 3017 147 3022 152
rect 3017 142 3126 147
rect 225 132 598 137
rect 809 132 1062 137
rect 1073 132 1446 137
rect 1457 132 1462 142
rect 1657 132 1854 137
rect 1881 132 1950 137
rect 1961 132 2382 137
rect 2561 132 2638 137
rect 593 127 814 132
rect 1457 127 1542 132
rect 2721 127 2726 142
rect 2873 132 2958 137
rect 2953 127 2958 132
rect 417 122 574 127
rect 937 122 1062 127
rect 1177 122 1206 127
rect 1217 122 1262 127
rect 1537 122 1606 127
rect 1617 122 2190 127
rect 2305 122 2390 127
rect 2513 122 2582 127
rect 2609 122 2726 127
rect 2905 122 2950 127
rect 2953 122 3006 127
rect 569 117 574 122
rect 849 117 942 122
rect 1057 117 1182 122
rect 1305 117 1438 122
rect 2945 117 2950 122
rect 337 112 422 117
rect 433 112 542 117
rect 569 112 854 117
rect 961 112 1038 117
rect 1281 112 1310 117
rect 1433 112 1558 117
rect 1761 112 1838 117
rect 1889 112 2358 117
rect 2553 112 2582 117
rect 433 107 438 112
rect 1577 107 1742 112
rect 1889 107 1894 112
rect 2577 107 2582 112
rect 2665 112 2694 117
rect 2745 112 2814 117
rect 2865 112 2934 117
rect 2945 112 2982 117
rect 3329 112 3382 117
rect 2665 107 2670 112
rect 161 102 326 107
rect 321 97 326 102
rect 385 102 438 107
rect 497 102 550 107
rect 385 97 390 102
rect 545 97 550 102
rect 873 102 990 107
rect 1153 102 1582 107
rect 1737 102 1894 107
rect 2033 102 2166 107
rect 2369 102 2462 107
rect 2577 102 2670 107
rect 873 97 878 102
rect 1153 97 1158 102
rect 1913 97 2014 102
rect 2161 97 2270 102
rect 2369 97 2374 102
rect 321 92 390 97
rect 409 92 438 97
rect 433 87 438 92
rect 497 92 526 97
rect 545 92 878 97
rect 897 92 1158 97
rect 1169 92 1294 97
rect 1401 92 1630 97
rect 1673 92 1918 97
rect 2009 92 2142 97
rect 2265 92 2374 97
rect 2921 92 3374 97
rect 497 87 502 92
rect 433 82 502 87
rect 953 82 1054 87
rect 1513 82 2246 87
rect 913 72 942 77
rect 937 57 942 72
rect 1209 72 1750 77
rect 2257 72 2718 77
rect 1209 67 1214 72
rect 1745 67 2126 72
rect 2257 67 2262 72
rect 1065 62 1214 67
rect 1409 62 1438 67
rect 1561 62 1726 67
rect 2121 62 2262 67
rect 1065 57 1070 62
rect 1433 57 1566 62
rect 937 52 1070 57
rect 1313 52 1398 57
rect 1393 47 1398 52
rect 1737 52 2102 57
rect 1737 47 1742 52
rect 1233 42 1302 47
rect 1393 42 1742 47
rect 2113 42 2486 47
rect 1297 27 1302 42
rect 2113 27 2118 42
rect 1297 22 2118 27
use AND2X2  AND2X2_0
timestamp 1712622712
transform 1 0 2632 0 -1 1170
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1712622712
transform 1 0 1368 0 -1 1170
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1712622712
transform 1 0 2864 0 -1 170
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1712622712
transform 1 0 1416 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1712622712
transform 1 0 1392 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1712622712
transform 1 0 1360 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1712622712
transform 1 0 2272 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1712622712
transform 1 0 1552 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1712622712
transform 1 0 1048 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1712622712
transform 1 0 2656 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1712622712
transform 1 0 1080 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1712622712
transform 1 0 2608 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1712622712
transform 1 0 2688 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1712622712
transform 1 0 848 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1712622712
transform 1 0 2272 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1712622712
transform 1 0 1584 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1712622712
transform 1 0 1472 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1712622712
transform 1 0 1760 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1712622712
transform 1 0 112 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1712622712
transform 1 0 1208 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_20
timestamp 1712622712
transform 1 0 1728 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1712622712
transform 1 0 1040 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1712622712
transform 1 0 1584 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_23
timestamp 1712622712
transform 1 0 3176 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1712622712
transform 1 0 3280 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_25
timestamp 1712622712
transform 1 0 2664 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_26
timestamp 1712622712
transform 1 0 2768 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_27
timestamp 1712622712
transform 1 0 2056 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_28
timestamp 1712622712
transform 1 0 816 0 -1 3170
box -8 -3 40 105
use AND2X2  AND2X2_29
timestamp 1712622712
transform 1 0 2104 0 -1 3170
box -8 -3 40 105
use AND2X2  AND2X2_30
timestamp 1712622712
transform 1 0 3032 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_31
timestamp 1712622712
transform 1 0 2912 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_32
timestamp 1712622712
transform 1 0 1856 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_33
timestamp 1712622712
transform 1 0 496 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_34
timestamp 1712622712
transform 1 0 928 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_35
timestamp 1712622712
transform 1 0 1384 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_36
timestamp 1712622712
transform 1 0 3272 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_37
timestamp 1712622712
transform 1 0 3344 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_38
timestamp 1712622712
transform 1 0 3280 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_39
timestamp 1712622712
transform 1 0 3368 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_40
timestamp 1712622712
transform 1 0 2856 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_41
timestamp 1712622712
transform 1 0 2888 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_42
timestamp 1712622712
transform 1 0 3064 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_43
timestamp 1712622712
transform 1 0 3312 0 1 570
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1712622712
transform 1 0 3120 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1712622712
transform 1 0 208 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1712622712
transform 1 0 416 0 -1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1712622712
transform 1 0 1624 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1712622712
transform 1 0 528 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1712622712
transform 1 0 2368 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1712622712
transform 1 0 488 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1712622712
transform 1 0 776 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1712622712
transform 1 0 392 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1712622712
transform 1 0 2080 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1712622712
transform 1 0 856 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1712622712
transform 1 0 2384 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1712622712
transform 1 0 88 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1712622712
transform 1 0 1240 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1712622712
transform 1 0 1896 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1712622712
transform 1 0 1120 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1712622712
transform 1 0 1216 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1712622712
transform 1 0 888 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1712622712
transform 1 0 816 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1712622712
transform 1 0 816 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1712622712
transform 1 0 1024 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1712622712
transform 1 0 1272 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1712622712
transform 1 0 1648 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1712622712
transform 1 0 1832 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1712622712
transform 1 0 1752 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1712622712
transform 1 0 1648 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1712622712
transform 1 0 1432 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_27
timestamp 1712622712
transform 1 0 2192 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_28
timestamp 1712622712
transform 1 0 2424 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_29
timestamp 1712622712
transform 1 0 2568 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_30
timestamp 1712622712
transform 1 0 2064 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_31
timestamp 1712622712
transform 1 0 3080 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_32
timestamp 1712622712
transform 1 0 2960 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_33
timestamp 1712622712
transform 1 0 2880 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_34
timestamp 1712622712
transform 1 0 2624 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_35
timestamp 1712622712
transform 1 0 2792 0 1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_36
timestamp 1712622712
transform 1 0 2616 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_37
timestamp 1712622712
transform 1 0 2632 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_38
timestamp 1712622712
transform 1 0 1776 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_39
timestamp 1712622712
transform 1 0 1728 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_40
timestamp 1712622712
transform 1 0 824 0 1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_41
timestamp 1712622712
transform 1 0 864 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_42
timestamp 1712622712
transform 1 0 2528 0 -1 3170
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1712622712
transform 1 0 1464 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1712622712
transform 1 0 1048 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1712622712
transform 1 0 664 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1712622712
transform 1 0 1080 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1712622712
transform 1 0 200 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1712622712
transform 1 0 224 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1712622712
transform 1 0 184 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1712622712
transform 1 0 2232 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1712622712
transform 1 0 2344 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1712622712
transform 1 0 2072 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1712622712
transform 1 0 944 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1712622712
transform 1 0 2224 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1712622712
transform 1 0 1552 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1712622712
transform 1 0 856 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1712622712
transform 1 0 408 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1712622712
transform 1 0 408 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1712622712
transform 1 0 440 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1712622712
transform 1 0 960 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1712622712
transform 1 0 464 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1712622712
transform 1 0 2224 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1712622712
transform 1 0 1720 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1712622712
transform 1 0 1920 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1712622712
transform 1 0 2560 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1712622712
transform 1 0 2616 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1712622712
transform 1 0 1048 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1712622712
transform 1 0 520 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1712622712
transform 1 0 488 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1712622712
transform 1 0 736 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1712622712
transform 1 0 1024 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1712622712
transform 1 0 488 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1712622712
transform 1 0 1856 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1712622712
transform 1 0 2368 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1712622712
transform 1 0 2384 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1712622712
transform 1 0 2240 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1712622712
transform 1 0 1560 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1712622712
transform 1 0 1224 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1712622712
transform 1 0 928 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1712622712
transform 1 0 712 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1712622712
transform 1 0 928 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1712622712
transform 1 0 600 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1712622712
transform 1 0 552 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1712622712
transform 1 0 1392 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1712622712
transform 1 0 2232 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1712622712
transform 1 0 1976 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1712622712
transform 1 0 2416 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1712622712
transform 1 0 2008 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1712622712
transform 1 0 1584 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1712622712
transform 1 0 496 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1712622712
transform 1 0 1520 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1712622712
transform 1 0 368 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1712622712
transform 1 0 360 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1712622712
transform 1 0 336 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1712622712
transform 1 0 2632 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1712622712
transform 1 0 2176 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1712622712
transform 1 0 1856 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_55
timestamp 1712622712
transform 1 0 1200 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1712622712
transform 1 0 2440 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_57
timestamp 1712622712
transform 1 0 1592 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_58
timestamp 1712622712
transform 1 0 2192 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_59
timestamp 1712622712
transform 1 0 1952 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_60
timestamp 1712622712
transform 1 0 2200 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_61
timestamp 1712622712
transform 1 0 2024 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_62
timestamp 1712622712
transform 1 0 192 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_63
timestamp 1712622712
transform 1 0 672 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_64
timestamp 1712622712
transform 1 0 288 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_65
timestamp 1712622712
transform 1 0 128 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_66
timestamp 1712622712
transform 1 0 376 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_67
timestamp 1712622712
transform 1 0 248 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_68
timestamp 1712622712
transform 1 0 328 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_69
timestamp 1712622712
transform 1 0 432 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_70
timestamp 1712622712
transform 1 0 1464 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_71
timestamp 1712622712
transform 1 0 1272 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1712622712
transform 1 0 2360 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_73
timestamp 1712622712
transform 1 0 1808 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_74
timestamp 1712622712
transform 1 0 2232 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_75
timestamp 1712622712
transform 1 0 2376 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_76
timestamp 1712622712
transform 1 0 96 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_77
timestamp 1712622712
transform 1 0 736 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_78
timestamp 1712622712
transform 1 0 136 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_79
timestamp 1712622712
transform 1 0 216 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_80
timestamp 1712622712
transform 1 0 1120 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_81
timestamp 1712622712
transform 1 0 1944 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_82
timestamp 1712622712
transform 1 0 2160 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_83
timestamp 1712622712
transform 1 0 2224 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_84
timestamp 1712622712
transform 1 0 1584 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_85
timestamp 1712622712
transform 1 0 1928 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_86
timestamp 1712622712
transform 1 0 1424 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_87
timestamp 1712622712
transform 1 0 1592 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_88
timestamp 1712622712
transform 1 0 1200 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_89
timestamp 1712622712
transform 1 0 1408 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_90
timestamp 1712622712
transform 1 0 1176 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_91
timestamp 1712622712
transform 1 0 1432 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_92
timestamp 1712622712
transform 1 0 808 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_93
timestamp 1712622712
transform 1 0 984 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_94
timestamp 1712622712
transform 1 0 1392 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_95
timestamp 1712622712
transform 1 0 1304 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_96
timestamp 1712622712
transform 1 0 720 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_97
timestamp 1712622712
transform 1 0 912 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_98
timestamp 1712622712
transform 1 0 648 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_99
timestamp 1712622712
transform 1 0 568 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_100
timestamp 1712622712
transform 1 0 448 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_101
timestamp 1712622712
transform 1 0 656 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_102
timestamp 1712622712
transform 1 0 376 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_103
timestamp 1712622712
transform 1 0 264 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_104
timestamp 1712622712
transform 1 0 368 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_105
timestamp 1712622712
transform 1 0 560 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_106
timestamp 1712622712
transform 1 0 208 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_107
timestamp 1712622712
transform 1 0 88 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_108
timestamp 1712622712
transform 1 0 416 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_109
timestamp 1712622712
transform 1 0 552 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_110
timestamp 1712622712
transform 1 0 264 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_111
timestamp 1712622712
transform 1 0 96 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_112
timestamp 1712622712
transform 1 0 1024 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_113
timestamp 1712622712
transform 1 0 416 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_114
timestamp 1712622712
transform 1 0 552 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_115
timestamp 1712622712
transform 1 0 240 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_116
timestamp 1712622712
transform 1 0 96 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_117
timestamp 1712622712
transform 1 0 448 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_118
timestamp 1712622712
transform 1 0 544 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_119
timestamp 1712622712
transform 1 0 240 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_120
timestamp 1712622712
transform 1 0 88 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_121
timestamp 1712622712
transform 1 0 408 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_122
timestamp 1712622712
transform 1 0 512 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_123
timestamp 1712622712
transform 1 0 184 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_124
timestamp 1712622712
transform 1 0 104 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_125
timestamp 1712622712
transform 1 0 480 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_126
timestamp 1712622712
transform 1 0 560 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_127
timestamp 1712622712
transform 1 0 200 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_128
timestamp 1712622712
transform 1 0 96 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_129
timestamp 1712622712
transform 1 0 432 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_130
timestamp 1712622712
transform 1 0 776 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_131
timestamp 1712622712
transform 1 0 232 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_132
timestamp 1712622712
transform 1 0 104 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_133
timestamp 1712622712
transform 1 0 512 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_134
timestamp 1712622712
transform 1 0 664 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_135
timestamp 1712622712
transform 1 0 320 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_136
timestamp 1712622712
transform 1 0 504 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_137
timestamp 1712622712
transform 1 0 920 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_138
timestamp 1712622712
transform 1 0 960 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_139
timestamp 1712622712
transform 1 0 864 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_140
timestamp 1712622712
transform 1 0 792 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_141
timestamp 1712622712
transform 1 0 1160 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_142
timestamp 1712622712
transform 1 0 1128 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_143
timestamp 1712622712
transform 1 0 1080 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_144
timestamp 1712622712
transform 1 0 1024 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_145
timestamp 1712622712
transform 1 0 1056 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_146
timestamp 1712622712
transform 1 0 1288 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_147
timestamp 1712622712
transform 1 0 1456 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_148
timestamp 1712622712
transform 1 0 1456 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_149
timestamp 1712622712
transform 1 0 1488 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_150
timestamp 1712622712
transform 1 0 1848 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_151
timestamp 1712622712
transform 1 0 1792 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_152
timestamp 1712622712
transform 1 0 1736 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_153
timestamp 1712622712
transform 1 0 1712 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_154
timestamp 1712622712
transform 1 0 2088 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_155
timestamp 1712622712
transform 1 0 1912 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_156
timestamp 1712622712
transform 1 0 2280 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_157
timestamp 1712622712
transform 1 0 2136 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_158
timestamp 1712622712
transform 1 0 2376 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_159
timestamp 1712622712
transform 1 0 2304 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_160
timestamp 1712622712
transform 1 0 2312 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_161
timestamp 1712622712
transform 1 0 2192 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_162
timestamp 1712622712
transform 1 0 2536 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_163
timestamp 1712622712
transform 1 0 2456 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_164
timestamp 1712622712
transform 1 0 2336 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_165
timestamp 1712622712
transform 1 0 2192 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_166
timestamp 1712622712
transform 1 0 2496 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_167
timestamp 1712622712
transform 1 0 2440 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_168
timestamp 1712622712
transform 1 0 2184 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_169
timestamp 1712622712
transform 1 0 2072 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_170
timestamp 1712622712
transform 1 0 2560 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_171
timestamp 1712622712
transform 1 0 2440 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_172
timestamp 1712622712
transform 1 0 2224 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_173
timestamp 1712622712
transform 1 0 2096 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_174
timestamp 1712622712
transform 1 0 1592 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_175
timestamp 1712622712
transform 1 0 1744 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_176
timestamp 1712622712
transform 1 0 1696 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_177
timestamp 1712622712
transform 1 0 1792 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_178
timestamp 1712622712
transform 1 0 1800 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_179
timestamp 1712622712
transform 1 0 1760 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_180
timestamp 1712622712
transform 1 0 1912 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_181
timestamp 1712622712
transform 1 0 2008 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_182
timestamp 1712622712
transform 1 0 1912 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_183
timestamp 1712622712
transform 1 0 1872 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_184
timestamp 1712622712
transform 1 0 2144 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_185
timestamp 1712622712
transform 1 0 2312 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_186
timestamp 1712622712
transform 1 0 2168 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_187
timestamp 1712622712
transform 1 0 2136 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_188
timestamp 1712622712
transform 1 0 2336 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_189
timestamp 1712622712
transform 1 0 2448 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_190
timestamp 1712622712
transform 1 0 2328 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_191
timestamp 1712622712
transform 1 0 2272 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_192
timestamp 1712622712
transform 1 0 2552 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_193
timestamp 1712622712
transform 1 0 2032 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_194
timestamp 1712622712
transform 1 0 1712 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_195
timestamp 1712622712
transform 1 0 2696 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_196
timestamp 1712622712
transform 1 0 3024 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_197
timestamp 1712622712
transform 1 0 2896 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_198
timestamp 1712622712
transform 1 0 3096 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_199
timestamp 1712622712
transform 1 0 2960 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_200
timestamp 1712622712
transform 1 0 2952 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_201
timestamp 1712622712
transform 1 0 2848 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_202
timestamp 1712622712
transform 1 0 2776 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_203
timestamp 1712622712
transform 1 0 2768 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_204
timestamp 1712622712
transform 1 0 2912 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_205
timestamp 1712622712
transform 1 0 2968 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_206
timestamp 1712622712
transform 1 0 3072 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_207
timestamp 1712622712
transform 1 0 3304 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_208
timestamp 1712622712
transform 1 0 3376 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_209
timestamp 1712622712
transform 1 0 3328 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_210
timestamp 1712622712
transform 1 0 2520 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_211
timestamp 1712622712
transform 1 0 2432 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_212
timestamp 1712622712
transform 1 0 1992 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_213
timestamp 1712622712
transform 1 0 2296 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_214
timestamp 1712622712
transform 1 0 2272 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_215
timestamp 1712622712
transform 1 0 2344 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_216
timestamp 1712622712
transform 1 0 2192 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_217
timestamp 1712622712
transform 1 0 2304 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_218
timestamp 1712622712
transform 1 0 2112 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_219
timestamp 1712622712
transform 1 0 2200 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_220
timestamp 1712622712
transform 1 0 1792 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_221
timestamp 1712622712
transform 1 0 1808 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_222
timestamp 1712622712
transform 1 0 1920 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_223
timestamp 1712622712
transform 1 0 1864 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_224
timestamp 1712622712
transform 1 0 1688 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_225
timestamp 1712622712
transform 1 0 1744 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_226
timestamp 1712622712
transform 1 0 1616 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_227
timestamp 1712622712
transform 1 0 1640 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_228
timestamp 1712622712
transform 1 0 1448 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_229
timestamp 1712622712
transform 1 0 1632 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_230
timestamp 1712622712
transform 1 0 1336 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_231
timestamp 1712622712
transform 1 0 1552 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_232
timestamp 1712622712
transform 1 0 1240 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_233
timestamp 1712622712
transform 1 0 1568 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_234
timestamp 1712622712
transform 1 0 1176 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_235
timestamp 1712622712
transform 1 0 1512 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_236
timestamp 1712622712
transform 1 0 1120 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_237
timestamp 1712622712
transform 1 0 1336 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_238
timestamp 1712622712
transform 1 0 944 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_239
timestamp 1712622712
transform 1 0 1224 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_240
timestamp 1712622712
transform 1 0 536 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_241
timestamp 1712622712
transform 1 0 1120 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_242
timestamp 1712622712
transform 1 0 640 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_243
timestamp 1712622712
transform 1 0 1008 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_244
timestamp 1712622712
transform 1 0 512 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_245
timestamp 1712622712
transform 1 0 736 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_246
timestamp 1712622712
transform 1 0 448 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_247
timestamp 1712622712
transform 1 0 680 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_248
timestamp 1712622712
transform 1 0 440 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_249
timestamp 1712622712
transform 1 0 640 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_250
timestamp 1712622712
transform 1 0 480 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_251
timestamp 1712622712
transform 1 0 680 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_252
timestamp 1712622712
transform 1 0 584 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_253
timestamp 1712622712
transform 1 0 736 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_254
timestamp 1712622712
transform 1 0 648 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_255
timestamp 1712622712
transform 1 0 672 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_256
timestamp 1712622712
transform 1 0 832 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_257
timestamp 1712622712
transform 1 0 624 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_258
timestamp 1712622712
transform 1 0 952 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_259
timestamp 1712622712
transform 1 0 704 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_260
timestamp 1712622712
transform 1 0 3328 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_261
timestamp 1712622712
transform 1 0 2216 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_262
timestamp 1712622712
transform 1 0 1960 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_263
timestamp 1712622712
transform 1 0 2136 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_264
timestamp 1712622712
transform 1 0 2384 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_265
timestamp 1712622712
transform 1 0 2504 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_266
timestamp 1712622712
transform 1 0 2592 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_267
timestamp 1712622712
transform 1 0 2744 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_268
timestamp 1712622712
transform 1 0 1144 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_269
timestamp 1712622712
transform 1 0 872 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_270
timestamp 1712622712
transform 1 0 2824 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_271
timestamp 1712622712
transform 1 0 712 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_272
timestamp 1712622712
transform 1 0 616 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_273
timestamp 1712622712
transform 1 0 496 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_274
timestamp 1712622712
transform 1 0 408 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_275
timestamp 1712622712
transform 1 0 328 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_276
timestamp 1712622712
transform 1 0 296 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_277
timestamp 1712622712
transform 1 0 232 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_278
timestamp 1712622712
transform 1 0 88 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_279
timestamp 1712622712
transform 1 0 152 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_280
timestamp 1712622712
transform 1 0 800 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_281
timestamp 1712622712
transform 1 0 2880 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_282
timestamp 1712622712
transform 1 0 952 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_283
timestamp 1712622712
transform 1 0 1200 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_284
timestamp 1712622712
transform 1 0 1440 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_285
timestamp 1712622712
transform 1 0 1496 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_286
timestamp 1712622712
transform 1 0 1584 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_287
timestamp 1712622712
transform 1 0 1656 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_288
timestamp 1712622712
transform 1 0 1752 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_289
timestamp 1712622712
transform 1 0 1832 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_290
timestamp 1712622712
transform 1 0 2032 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_291
timestamp 1712622712
transform 1 0 2312 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_292
timestamp 1712622712
transform 1 0 2664 0 -1 2570
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1712622712
transform 1 0 2088 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1712622712
transform 1 0 1912 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1712622712
transform 1 0 3408 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1712622712
transform 1 0 3144 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1712622712
transform 1 0 2688 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1712622712
transform 1 0 2720 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1712622712
transform 1 0 3200 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1712622712
transform 1 0 3128 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1712622712
transform 1 0 1744 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1712622712
transform 1 0 2936 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1712622712
transform 1 0 3072 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1712622712
transform 1 0 3232 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1712622712
transform 1 0 3208 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1712622712
transform 1 0 2320 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1712622712
transform 1 0 2136 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1712622712
transform 1 0 2296 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1712622712
transform 1 0 1888 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1712622712
transform 1 0 1720 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1712622712
transform 1 0 1736 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1712622712
transform 1 0 3184 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1712622712
transform 1 0 2448 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_21
timestamp 1712622712
transform 1 0 2792 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_22
timestamp 1712622712
transform 1 0 2976 0 1 2770
box -5 -3 28 105
use BUFX2  BUFX2_23
timestamp 1712622712
transform 1 0 3168 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1712622712
transform 1 0 3000 0 -1 2970
box -5 -3 28 105
use BUFX2  BUFX2_25
timestamp 1712622712
transform 1 0 2272 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_26
timestamp 1712622712
transform 1 0 2408 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_27
timestamp 1712622712
transform 1 0 2112 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_28
timestamp 1712622712
transform 1 0 2448 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_29
timestamp 1712622712
transform 1 0 2264 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_30
timestamp 1712622712
transform 1 0 2384 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_31
timestamp 1712622712
transform 1 0 1616 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_32
timestamp 1712622712
transform 1 0 3216 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_33
timestamp 1712622712
transform 1 0 1672 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_34
timestamp 1712622712
transform 1 0 3088 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_35
timestamp 1712622712
transform 1 0 2656 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_36
timestamp 1712622712
transform 1 0 1712 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_37
timestamp 1712622712
transform 1 0 1928 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_38
timestamp 1712622712
transform 1 0 2856 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_39
timestamp 1712622712
transform 1 0 1584 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_40
timestamp 1712622712
transform 1 0 1448 0 -1 2970
box -5 -3 28 105
use BUFX2  BUFX2_41
timestamp 1712622712
transform 1 0 1304 0 -1 2970
box -5 -3 28 105
use BUFX2  BUFX2_42
timestamp 1712622712
transform 1 0 1696 0 -1 1770
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1712622712
transform 1 0 3328 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1712622712
transform 1 0 3312 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1712622712
transform 1 0 3096 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1712622712
transform 1 0 3152 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1712622712
transform 1 0 2800 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1712622712
transform 1 0 2920 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1712622712
transform 1 0 3040 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1712622712
transform 1 0 3184 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1712622712
transform 1 0 3328 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1712622712
transform 1 0 2776 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1712622712
transform 1 0 2744 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1712622712
transform 1 0 2968 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1712622712
transform 1 0 3048 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1712622712
transform 1 0 3048 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1712622712
transform 1 0 3328 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1712622712
transform 1 0 3224 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1712622712
transform 1 0 3104 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1712622712
transform 1 0 2944 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1712622712
transform 1 0 2736 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1712622712
transform 1 0 3112 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1712622712
transform 1 0 3336 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1712622712
transform 1 0 1152 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1712622712
transform 1 0 856 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1712622712
transform 1 0 744 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1712622712
transform 1 0 632 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1712622712
transform 1 0 416 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1712622712
transform 1 0 304 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1712622712
transform 1 0 200 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1712622712
transform 1 0 192 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1712622712
transform 1 0 128 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1712622712
transform 1 0 80 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1712622712
transform 1 0 88 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1712622712
transform 1 0 528 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1712622712
transform 1 0 968 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1712622712
transform 1 0 1024 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1712622712
transform 1 0 1256 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1712622712
transform 1 0 1360 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1712622712
transform 1 0 1464 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1712622712
transform 1 0 1520 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1712622712
transform 1 0 1632 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1712622712
transform 1 0 1768 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1712622712
transform 1 0 1968 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1712622712
transform 1 0 2264 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1712622712
transform 1 0 2168 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1712622712
transform 1 0 1872 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1712622712
transform 1 0 2072 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1712622712
transform 1 0 2368 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1712622712
transform 1 0 2464 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1712622712
transform 1 0 2560 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1712622712
transform 1 0 2760 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1712622712
transform 1 0 2960 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1712622712
transform 1 0 2856 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1712622712
transform 1 0 2664 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1712622712
transform 1 0 2896 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1712622712
transform 1 0 952 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1712622712
transform 1 0 768 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1712622712
transform 1 0 424 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1712622712
transform 1 0 464 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1712622712
transform 1 0 304 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1712622712
transform 1 0 248 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1712622712
transform 1 0 264 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1712622712
transform 1 0 200 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1712622712
transform 1 0 80 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1712622712
transform 1 0 136 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1712622712
transform 1 0 80 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1712622712
transform 1 0 1056 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1712622712
transform 1 0 1016 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1712622712
transform 1 0 1200 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1712622712
transform 1 0 1376 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1712622712
transform 1 0 1352 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1712622712
transform 1 0 1472 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1712622712
transform 1 0 1520 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1712622712
transform 1 0 1832 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1712622712
transform 1 0 1680 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1712622712
transform 1 0 1976 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1712622712
transform 1 0 2144 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1712622712
transform 1 0 2240 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1712622712
transform 1 0 2056 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1712622712
transform 1 0 2416 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1712622712
transform 1 0 2728 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1712622712
transform 1 0 2680 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1712622712
transform 1 0 2600 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1712622712
transform 1 0 2808 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1712622712
transform 1 0 3096 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1712622712
transform 1 0 2888 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1712622712
transform 1 0 2592 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1712622712
transform 1 0 3104 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1712622712
transform 1 0 2992 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1712622712
transform 1 0 1104 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1712622712
transform 1 0 784 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1712622712
transform 1 0 672 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1712622712
transform 1 0 568 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1712622712
transform 1 0 368 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1712622712
transform 1 0 352 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1712622712
transform 1 0 304 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1712622712
transform 1 0 232 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1712622712
transform 1 0 192 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1712622712
transform 1 0 80 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1712622712
transform 1 0 112 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1712622712
transform 1 0 888 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1712622712
transform 1 0 992 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1712622712
transform 1 0 1208 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1712622712
transform 1 0 1320 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1712622712
transform 1 0 1416 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1712622712
transform 1 0 1568 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1712622712
transform 1 0 1680 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1712622712
transform 1 0 1904 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1712622712
transform 1 0 1792 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1712622712
transform 1 0 2024 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1712622712
transform 1 0 2144 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1712622712
transform 1 0 2208 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1712622712
transform 1 0 1896 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1712622712
transform 1 0 2344 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1712622712
transform 1 0 2456 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1712622712
transform 1 0 2520 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1712622712
transform 1 0 2568 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1712622712
transform 1 0 2752 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1712622712
transform 1 0 2944 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1712622712
transform 1 0 2880 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1712622712
transform 1 0 2640 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1712622712
transform 1 0 3336 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1712622712
transform 1 0 3296 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1712622712
transform 1 0 3200 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1712622712
transform 1 0 3232 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1712622712
transform 1 0 3232 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1712622712
transform 1 0 3056 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1712622712
transform 1 0 3160 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1712622712
transform 1 0 3336 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_128
timestamp 1712622712
transform 1 0 3328 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1712622712
transform 1 0 3336 0 -1 2570
box -8 -3 104 105
use FILL  FILL_0
timestamp 1712622712
transform 1 0 3424 0 1 3170
box -8 -3 16 105
use FILL  FILL_1
timestamp 1712622712
transform 1 0 3416 0 1 3170
box -8 -3 16 105
use FILL  FILL_2
timestamp 1712622712
transform 1 0 3360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3
timestamp 1712622712
transform 1 0 3320 0 1 3170
box -8 -3 16 105
use FILL  FILL_4
timestamp 1712622712
transform 1 0 3296 0 1 3170
box -8 -3 16 105
use FILL  FILL_5
timestamp 1712622712
transform 1 0 3192 0 1 3170
box -8 -3 16 105
use FILL  FILL_6
timestamp 1712622712
transform 1 0 3088 0 1 3170
box -8 -3 16 105
use FILL  FILL_7
timestamp 1712622712
transform 1 0 3080 0 1 3170
box -8 -3 16 105
use FILL  FILL_8
timestamp 1712622712
transform 1 0 3072 0 1 3170
box -8 -3 16 105
use FILL  FILL_9
timestamp 1712622712
transform 1 0 3064 0 1 3170
box -8 -3 16 105
use FILL  FILL_10
timestamp 1712622712
transform 1 0 2952 0 1 3170
box -8 -3 16 105
use FILL  FILL_11
timestamp 1712622712
transform 1 0 2912 0 1 3170
box -8 -3 16 105
use FILL  FILL_12
timestamp 1712622712
transform 1 0 2904 0 1 3170
box -8 -3 16 105
use FILL  FILL_13
timestamp 1712622712
transform 1 0 2864 0 1 3170
box -8 -3 16 105
use FILL  FILL_14
timestamp 1712622712
transform 1 0 2856 0 1 3170
box -8 -3 16 105
use FILL  FILL_15
timestamp 1712622712
transform 1 0 2848 0 1 3170
box -8 -3 16 105
use FILL  FILL_16
timestamp 1712622712
transform 1 0 2784 0 1 3170
box -8 -3 16 105
use FILL  FILL_17
timestamp 1712622712
transform 1 0 2776 0 1 3170
box -8 -3 16 105
use FILL  FILL_18
timestamp 1712622712
transform 1 0 2672 0 1 3170
box -8 -3 16 105
use FILL  FILL_19
timestamp 1712622712
transform 1 0 2664 0 1 3170
box -8 -3 16 105
use FILL  FILL_20
timestamp 1712622712
transform 1 0 2600 0 1 3170
box -8 -3 16 105
use FILL  FILL_21
timestamp 1712622712
transform 1 0 2592 0 1 3170
box -8 -3 16 105
use FILL  FILL_22
timestamp 1712622712
transform 1 0 2584 0 1 3170
box -8 -3 16 105
use FILL  FILL_23
timestamp 1712622712
transform 1 0 2528 0 1 3170
box -8 -3 16 105
use FILL  FILL_24
timestamp 1712622712
transform 1 0 2520 0 1 3170
box -8 -3 16 105
use FILL  FILL_25
timestamp 1712622712
transform 1 0 2488 0 1 3170
box -8 -3 16 105
use FILL  FILL_26
timestamp 1712622712
transform 1 0 2480 0 1 3170
box -8 -3 16 105
use FILL  FILL_27
timestamp 1712622712
transform 1 0 2440 0 1 3170
box -8 -3 16 105
use FILL  FILL_28
timestamp 1712622712
transform 1 0 2416 0 1 3170
box -8 -3 16 105
use FILL  FILL_29
timestamp 1712622712
transform 1 0 2384 0 1 3170
box -8 -3 16 105
use FILL  FILL_30
timestamp 1712622712
transform 1 0 2344 0 1 3170
box -8 -3 16 105
use FILL  FILL_31
timestamp 1712622712
transform 1 0 2336 0 1 3170
box -8 -3 16 105
use FILL  FILL_32
timestamp 1712622712
transform 1 0 2288 0 1 3170
box -8 -3 16 105
use FILL  FILL_33
timestamp 1712622712
transform 1 0 2248 0 1 3170
box -8 -3 16 105
use FILL  FILL_34
timestamp 1712622712
transform 1 0 2240 0 1 3170
box -8 -3 16 105
use FILL  FILL_35
timestamp 1712622712
transform 1 0 2232 0 1 3170
box -8 -3 16 105
use FILL  FILL_36
timestamp 1712622712
transform 1 0 2224 0 1 3170
box -8 -3 16 105
use FILL  FILL_37
timestamp 1712622712
transform 1 0 2136 0 1 3170
box -8 -3 16 105
use FILL  FILL_38
timestamp 1712622712
transform 1 0 2128 0 1 3170
box -8 -3 16 105
use FILL  FILL_39
timestamp 1712622712
transform 1 0 2120 0 1 3170
box -8 -3 16 105
use FILL  FILL_40
timestamp 1712622712
transform 1 0 2048 0 1 3170
box -8 -3 16 105
use FILL  FILL_41
timestamp 1712622712
transform 1 0 2008 0 1 3170
box -8 -3 16 105
use FILL  FILL_42
timestamp 1712622712
transform 1 0 1968 0 1 3170
box -8 -3 16 105
use FILL  FILL_43
timestamp 1712622712
transform 1 0 1960 0 1 3170
box -8 -3 16 105
use FILL  FILL_44
timestamp 1712622712
transform 1 0 1896 0 1 3170
box -8 -3 16 105
use FILL  FILL_45
timestamp 1712622712
transform 1 0 1888 0 1 3170
box -8 -3 16 105
use FILL  FILL_46
timestamp 1712622712
transform 1 0 1832 0 1 3170
box -8 -3 16 105
use FILL  FILL_47
timestamp 1712622712
transform 1 0 1824 0 1 3170
box -8 -3 16 105
use FILL  FILL_48
timestamp 1712622712
transform 1 0 1792 0 1 3170
box -8 -3 16 105
use FILL  FILL_49
timestamp 1712622712
transform 1 0 1752 0 1 3170
box -8 -3 16 105
use FILL  FILL_50
timestamp 1712622712
transform 1 0 1720 0 1 3170
box -8 -3 16 105
use FILL  FILL_51
timestamp 1712622712
transform 1 0 1712 0 1 3170
box -8 -3 16 105
use FILL  FILL_52
timestamp 1712622712
transform 1 0 1704 0 1 3170
box -8 -3 16 105
use FILL  FILL_53
timestamp 1712622712
transform 1 0 1632 0 1 3170
box -8 -3 16 105
use FILL  FILL_54
timestamp 1712622712
transform 1 0 1624 0 1 3170
box -8 -3 16 105
use FILL  FILL_55
timestamp 1712622712
transform 1 0 1616 0 1 3170
box -8 -3 16 105
use FILL  FILL_56
timestamp 1712622712
transform 1 0 1608 0 1 3170
box -8 -3 16 105
use FILL  FILL_57
timestamp 1712622712
transform 1 0 1576 0 1 3170
box -8 -3 16 105
use FILL  FILL_58
timestamp 1712622712
transform 1 0 1552 0 1 3170
box -8 -3 16 105
use FILL  FILL_59
timestamp 1712622712
transform 1 0 1512 0 1 3170
box -8 -3 16 105
use FILL  FILL_60
timestamp 1712622712
transform 1 0 1472 0 1 3170
box -8 -3 16 105
use FILL  FILL_61
timestamp 1712622712
transform 1 0 1464 0 1 3170
box -8 -3 16 105
use FILL  FILL_62
timestamp 1712622712
transform 1 0 1456 0 1 3170
box -8 -3 16 105
use FILL  FILL_63
timestamp 1712622712
transform 1 0 1448 0 1 3170
box -8 -3 16 105
use FILL  FILL_64
timestamp 1712622712
transform 1 0 1376 0 1 3170
box -8 -3 16 105
use FILL  FILL_65
timestamp 1712622712
transform 1 0 1368 0 1 3170
box -8 -3 16 105
use FILL  FILL_66
timestamp 1712622712
transform 1 0 1344 0 1 3170
box -8 -3 16 105
use FILL  FILL_67
timestamp 1712622712
transform 1 0 1304 0 1 3170
box -8 -3 16 105
use FILL  FILL_68
timestamp 1712622712
transform 1 0 1296 0 1 3170
box -8 -3 16 105
use FILL  FILL_69
timestamp 1712622712
transform 1 0 1264 0 1 3170
box -8 -3 16 105
use FILL  FILL_70
timestamp 1712622712
transform 1 0 1256 0 1 3170
box -8 -3 16 105
use FILL  FILL_71
timestamp 1712622712
transform 1 0 1232 0 1 3170
box -8 -3 16 105
use FILL  FILL_72
timestamp 1712622712
transform 1 0 1192 0 1 3170
box -8 -3 16 105
use FILL  FILL_73
timestamp 1712622712
transform 1 0 1184 0 1 3170
box -8 -3 16 105
use FILL  FILL_74
timestamp 1712622712
transform 1 0 1176 0 1 3170
box -8 -3 16 105
use FILL  FILL_75
timestamp 1712622712
transform 1 0 1168 0 1 3170
box -8 -3 16 105
use FILL  FILL_76
timestamp 1712622712
transform 1 0 1096 0 1 3170
box -8 -3 16 105
use FILL  FILL_77
timestamp 1712622712
transform 1 0 1088 0 1 3170
box -8 -3 16 105
use FILL  FILL_78
timestamp 1712622712
transform 1 0 1080 0 1 3170
box -8 -3 16 105
use FILL  FILL_79
timestamp 1712622712
transform 1 0 1072 0 1 3170
box -8 -3 16 105
use FILL  FILL_80
timestamp 1712622712
transform 1 0 984 0 1 3170
box -8 -3 16 105
use FILL  FILL_81
timestamp 1712622712
transform 1 0 976 0 1 3170
box -8 -3 16 105
use FILL  FILL_82
timestamp 1712622712
transform 1 0 968 0 1 3170
box -8 -3 16 105
use FILL  FILL_83
timestamp 1712622712
transform 1 0 960 0 1 3170
box -8 -3 16 105
use FILL  FILL_84
timestamp 1712622712
transform 1 0 872 0 1 3170
box -8 -3 16 105
use FILL  FILL_85
timestamp 1712622712
transform 1 0 864 0 1 3170
box -8 -3 16 105
use FILL  FILL_86
timestamp 1712622712
transform 1 0 856 0 1 3170
box -8 -3 16 105
use FILL  FILL_87
timestamp 1712622712
transform 1 0 816 0 1 3170
box -8 -3 16 105
use FILL  FILL_88
timestamp 1712622712
transform 1 0 808 0 1 3170
box -8 -3 16 105
use FILL  FILL_89
timestamp 1712622712
transform 1 0 744 0 1 3170
box -8 -3 16 105
use FILL  FILL_90
timestamp 1712622712
transform 1 0 736 0 1 3170
box -8 -3 16 105
use FILL  FILL_91
timestamp 1712622712
transform 1 0 728 0 1 3170
box -8 -3 16 105
use FILL  FILL_92
timestamp 1712622712
transform 1 0 720 0 1 3170
box -8 -3 16 105
use FILL  FILL_93
timestamp 1712622712
transform 1 0 632 0 1 3170
box -8 -3 16 105
use FILL  FILL_94
timestamp 1712622712
transform 1 0 624 0 1 3170
box -8 -3 16 105
use FILL  FILL_95
timestamp 1712622712
transform 1 0 616 0 1 3170
box -8 -3 16 105
use FILL  FILL_96
timestamp 1712622712
transform 1 0 608 0 1 3170
box -8 -3 16 105
use FILL  FILL_97
timestamp 1712622712
transform 1 0 600 0 1 3170
box -8 -3 16 105
use FILL  FILL_98
timestamp 1712622712
transform 1 0 528 0 1 3170
box -8 -3 16 105
use FILL  FILL_99
timestamp 1712622712
transform 1 0 488 0 1 3170
box -8 -3 16 105
use FILL  FILL_100
timestamp 1712622712
transform 1 0 480 0 1 3170
box -8 -3 16 105
use FILL  FILL_101
timestamp 1712622712
transform 1 0 432 0 1 3170
box -8 -3 16 105
use FILL  FILL_102
timestamp 1712622712
transform 1 0 424 0 1 3170
box -8 -3 16 105
use FILL  FILL_103
timestamp 1712622712
transform 1 0 416 0 1 3170
box -8 -3 16 105
use FILL  FILL_104
timestamp 1712622712
transform 1 0 360 0 1 3170
box -8 -3 16 105
use FILL  FILL_105
timestamp 1712622712
transform 1 0 352 0 1 3170
box -8 -3 16 105
use FILL  FILL_106
timestamp 1712622712
transform 1 0 344 0 1 3170
box -8 -3 16 105
use FILL  FILL_107
timestamp 1712622712
transform 1 0 240 0 1 3170
box -8 -3 16 105
use FILL  FILL_108
timestamp 1712622712
transform 1 0 232 0 1 3170
box -8 -3 16 105
use FILL  FILL_109
timestamp 1712622712
transform 1 0 128 0 1 3170
box -8 -3 16 105
use FILL  FILL_110
timestamp 1712622712
transform 1 0 120 0 1 3170
box -8 -3 16 105
use FILL  FILL_111
timestamp 1712622712
transform 1 0 112 0 1 3170
box -8 -3 16 105
use FILL  FILL_112
timestamp 1712622712
transform 1 0 104 0 1 3170
box -8 -3 16 105
use FILL  FILL_113
timestamp 1712622712
transform 1 0 96 0 1 3170
box -8 -3 16 105
use FILL  FILL_114
timestamp 1712622712
transform 1 0 72 0 1 3170
box -8 -3 16 105
use FILL  FILL_115
timestamp 1712622712
transform 1 0 3424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_116
timestamp 1712622712
transform 1 0 3392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_117
timestamp 1712622712
transform 1 0 3288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_118
timestamp 1712622712
transform 1 0 3280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_119
timestamp 1712622712
transform 1 0 3272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_120
timestamp 1712622712
transform 1 0 3200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_121
timestamp 1712622712
transform 1 0 3192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_122
timestamp 1712622712
transform 1 0 3168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_123
timestamp 1712622712
transform 1 0 3160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_124
timestamp 1712622712
transform 1 0 3152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_125
timestamp 1712622712
transform 1 0 3128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_126
timestamp 1712622712
transform 1 0 3088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_127
timestamp 1712622712
transform 1 0 3080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_128
timestamp 1712622712
transform 1 0 3072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_129
timestamp 1712622712
transform 1 0 3040 0 -1 3170
box -8 -3 16 105
use FILL  FILL_130
timestamp 1712622712
transform 1 0 3008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_131
timestamp 1712622712
transform 1 0 3000 0 -1 3170
box -8 -3 16 105
use FILL  FILL_132
timestamp 1712622712
transform 1 0 2992 0 -1 3170
box -8 -3 16 105
use FILL  FILL_133
timestamp 1712622712
transform 1 0 2968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_134
timestamp 1712622712
transform 1 0 2928 0 -1 3170
box -8 -3 16 105
use FILL  FILL_135
timestamp 1712622712
transform 1 0 2920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_136
timestamp 1712622712
transform 1 0 2912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_137
timestamp 1712622712
transform 1 0 2904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_138
timestamp 1712622712
transform 1 0 2832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_139
timestamp 1712622712
transform 1 0 2824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_140
timestamp 1712622712
transform 1 0 2816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_141
timestamp 1712622712
transform 1 0 2808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_142
timestamp 1712622712
transform 1 0 2784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_143
timestamp 1712622712
transform 1 0 2776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_144
timestamp 1712622712
transform 1 0 2712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_145
timestamp 1712622712
transform 1 0 2704 0 -1 3170
box -8 -3 16 105
use FILL  FILL_146
timestamp 1712622712
transform 1 0 2696 0 -1 3170
box -8 -3 16 105
use FILL  FILL_147
timestamp 1712622712
transform 1 0 2688 0 -1 3170
box -8 -3 16 105
use FILL  FILL_148
timestamp 1712622712
transform 1 0 2680 0 -1 3170
box -8 -3 16 105
use FILL  FILL_149
timestamp 1712622712
transform 1 0 2608 0 -1 3170
box -8 -3 16 105
use FILL  FILL_150
timestamp 1712622712
transform 1 0 2600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_151
timestamp 1712622712
transform 1 0 2592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_152
timestamp 1712622712
transform 1 0 2584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_153
timestamp 1712622712
transform 1 0 2520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_154
timestamp 1712622712
transform 1 0 2512 0 -1 3170
box -8 -3 16 105
use FILL  FILL_155
timestamp 1712622712
transform 1 0 2504 0 -1 3170
box -8 -3 16 105
use FILL  FILL_156
timestamp 1712622712
transform 1 0 2480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_157
timestamp 1712622712
transform 1 0 2472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_158
timestamp 1712622712
transform 1 0 2464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_159
timestamp 1712622712
transform 1 0 2408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_160
timestamp 1712622712
transform 1 0 2400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_161
timestamp 1712622712
transform 1 0 2392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_162
timestamp 1712622712
transform 1 0 2384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_163
timestamp 1712622712
transform 1 0 2296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_164
timestamp 1712622712
transform 1 0 2288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_165
timestamp 1712622712
transform 1 0 2280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_166
timestamp 1712622712
transform 1 0 2272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_167
timestamp 1712622712
transform 1 0 2192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_168
timestamp 1712622712
transform 1 0 2184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_169
timestamp 1712622712
transform 1 0 2176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_170
timestamp 1712622712
transform 1 0 2168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_171
timestamp 1712622712
transform 1 0 2096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_172
timestamp 1712622712
transform 1 0 2088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_173
timestamp 1712622712
transform 1 0 2056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_174
timestamp 1712622712
transform 1 0 2048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_175
timestamp 1712622712
transform 1 0 2024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_176
timestamp 1712622712
transform 1 0 1984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_177
timestamp 1712622712
transform 1 0 1976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_178
timestamp 1712622712
transform 1 0 1936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_179
timestamp 1712622712
transform 1 0 1928 0 -1 3170
box -8 -3 16 105
use FILL  FILL_180
timestamp 1712622712
transform 1 0 1920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_181
timestamp 1712622712
transform 1 0 1856 0 -1 3170
box -8 -3 16 105
use FILL  FILL_182
timestamp 1712622712
transform 1 0 1848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_183
timestamp 1712622712
transform 1 0 1824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_184
timestamp 1712622712
transform 1 0 1816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_185
timestamp 1712622712
transform 1 0 1808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_186
timestamp 1712622712
transform 1 0 1768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_187
timestamp 1712622712
transform 1 0 1760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_188
timestamp 1712622712
transform 1 0 1720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_189
timestamp 1712622712
transform 1 0 1712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_190
timestamp 1712622712
transform 1 0 1704 0 -1 3170
box -8 -3 16 105
use FILL  FILL_191
timestamp 1712622712
transform 1 0 1696 0 -1 3170
box -8 -3 16 105
use FILL  FILL_192
timestamp 1712622712
transform 1 0 1624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_193
timestamp 1712622712
transform 1 0 1616 0 -1 3170
box -8 -3 16 105
use FILL  FILL_194
timestamp 1712622712
transform 1 0 1608 0 -1 3170
box -8 -3 16 105
use FILL  FILL_195
timestamp 1712622712
transform 1 0 1600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_196
timestamp 1712622712
transform 1 0 1592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_197
timestamp 1712622712
transform 1 0 1544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_198
timestamp 1712622712
transform 1 0 1504 0 -1 3170
box -8 -3 16 105
use FILL  FILL_199
timestamp 1712622712
transform 1 0 1496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_200
timestamp 1712622712
transform 1 0 1488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_201
timestamp 1712622712
transform 1 0 1480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_202
timestamp 1712622712
transform 1 0 1472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_203
timestamp 1712622712
transform 1 0 1408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_204
timestamp 1712622712
transform 1 0 1400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_205
timestamp 1712622712
transform 1 0 1392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_206
timestamp 1712622712
transform 1 0 1384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_207
timestamp 1712622712
transform 1 0 1376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_208
timestamp 1712622712
transform 1 0 1296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_209
timestamp 1712622712
transform 1 0 1288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_210
timestamp 1712622712
transform 1 0 1280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_211
timestamp 1712622712
transform 1 0 1272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_212
timestamp 1712622712
transform 1 0 1264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_213
timestamp 1712622712
transform 1 0 1184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_214
timestamp 1712622712
transform 1 0 1176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_215
timestamp 1712622712
transform 1 0 1168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_216
timestamp 1712622712
transform 1 0 1160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_217
timestamp 1712622712
transform 1 0 1080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_218
timestamp 1712622712
transform 1 0 1072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_219
timestamp 1712622712
transform 1 0 1064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_220
timestamp 1712622712
transform 1 0 1056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_221
timestamp 1712622712
transform 1 0 1048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_222
timestamp 1712622712
transform 1 0 984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_223
timestamp 1712622712
transform 1 0 976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_224
timestamp 1712622712
transform 1 0 944 0 -1 3170
box -8 -3 16 105
use FILL  FILL_225
timestamp 1712622712
transform 1 0 936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_226
timestamp 1712622712
transform 1 0 928 0 -1 3170
box -8 -3 16 105
use FILL  FILL_227
timestamp 1712622712
transform 1 0 920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_228
timestamp 1712622712
transform 1 0 856 0 -1 3170
box -8 -3 16 105
use FILL  FILL_229
timestamp 1712622712
transform 1 0 848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_230
timestamp 1712622712
transform 1 0 784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_231
timestamp 1712622712
transform 1 0 776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_232
timestamp 1712622712
transform 1 0 728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_233
timestamp 1712622712
transform 1 0 720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_234
timestamp 1712622712
transform 1 0 632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_235
timestamp 1712622712
transform 1 0 624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_236
timestamp 1712622712
transform 1 0 616 0 -1 3170
box -8 -3 16 105
use FILL  FILL_237
timestamp 1712622712
transform 1 0 608 0 -1 3170
box -8 -3 16 105
use FILL  FILL_238
timestamp 1712622712
transform 1 0 528 0 -1 3170
box -8 -3 16 105
use FILL  FILL_239
timestamp 1712622712
transform 1 0 520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_240
timestamp 1712622712
transform 1 0 472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_241
timestamp 1712622712
transform 1 0 464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_242
timestamp 1712622712
transform 1 0 408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_243
timestamp 1712622712
transform 1 0 400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_244
timestamp 1712622712
transform 1 0 296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_245
timestamp 1712622712
transform 1 0 288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_246
timestamp 1712622712
transform 1 0 280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_247
timestamp 1712622712
transform 1 0 192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_248
timestamp 1712622712
transform 1 0 184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_249
timestamp 1712622712
transform 1 0 176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_250
timestamp 1712622712
transform 1 0 72 0 -1 3170
box -8 -3 16 105
use FILL  FILL_251
timestamp 1712622712
transform 1 0 3424 0 1 2970
box -8 -3 16 105
use FILL  FILL_252
timestamp 1712622712
transform 1 0 3416 0 1 2970
box -8 -3 16 105
use FILL  FILL_253
timestamp 1712622712
transform 1 0 3408 0 1 2970
box -8 -3 16 105
use FILL  FILL_254
timestamp 1712622712
transform 1 0 3400 0 1 2970
box -8 -3 16 105
use FILL  FILL_255
timestamp 1712622712
transform 1 0 3392 0 1 2970
box -8 -3 16 105
use FILL  FILL_256
timestamp 1712622712
transform 1 0 3384 0 1 2970
box -8 -3 16 105
use FILL  FILL_257
timestamp 1712622712
transform 1 0 3376 0 1 2970
box -8 -3 16 105
use FILL  FILL_258
timestamp 1712622712
transform 1 0 3336 0 1 2970
box -8 -3 16 105
use FILL  FILL_259
timestamp 1712622712
transform 1 0 3328 0 1 2970
box -8 -3 16 105
use FILL  FILL_260
timestamp 1712622712
transform 1 0 3320 0 1 2970
box -8 -3 16 105
use FILL  FILL_261
timestamp 1712622712
transform 1 0 3312 0 1 2970
box -8 -3 16 105
use FILL  FILL_262
timestamp 1712622712
transform 1 0 3304 0 1 2970
box -8 -3 16 105
use FILL  FILL_263
timestamp 1712622712
transform 1 0 3232 0 1 2970
box -8 -3 16 105
use FILL  FILL_264
timestamp 1712622712
transform 1 0 3224 0 1 2970
box -8 -3 16 105
use FILL  FILL_265
timestamp 1712622712
transform 1 0 3216 0 1 2970
box -8 -3 16 105
use FILL  FILL_266
timestamp 1712622712
transform 1 0 3208 0 1 2970
box -8 -3 16 105
use FILL  FILL_267
timestamp 1712622712
transform 1 0 3200 0 1 2970
box -8 -3 16 105
use FILL  FILL_268
timestamp 1712622712
transform 1 0 3096 0 1 2970
box -8 -3 16 105
use FILL  FILL_269
timestamp 1712622712
transform 1 0 3088 0 1 2970
box -8 -3 16 105
use FILL  FILL_270
timestamp 1712622712
transform 1 0 3080 0 1 2970
box -8 -3 16 105
use FILL  FILL_271
timestamp 1712622712
transform 1 0 3072 0 1 2970
box -8 -3 16 105
use FILL  FILL_272
timestamp 1712622712
transform 1 0 3008 0 1 2970
box -8 -3 16 105
use FILL  FILL_273
timestamp 1712622712
transform 1 0 3000 0 1 2970
box -8 -3 16 105
use FILL  FILL_274
timestamp 1712622712
transform 1 0 2992 0 1 2970
box -8 -3 16 105
use FILL  FILL_275
timestamp 1712622712
transform 1 0 2984 0 1 2970
box -8 -3 16 105
use FILL  FILL_276
timestamp 1712622712
transform 1 0 2976 0 1 2970
box -8 -3 16 105
use FILL  FILL_277
timestamp 1712622712
transform 1 0 2968 0 1 2970
box -8 -3 16 105
use FILL  FILL_278
timestamp 1712622712
transform 1 0 2920 0 1 2970
box -8 -3 16 105
use FILL  FILL_279
timestamp 1712622712
transform 1 0 2912 0 1 2970
box -8 -3 16 105
use FILL  FILL_280
timestamp 1712622712
transform 1 0 2904 0 1 2970
box -8 -3 16 105
use FILL  FILL_281
timestamp 1712622712
transform 1 0 2864 0 1 2970
box -8 -3 16 105
use FILL  FILL_282
timestamp 1712622712
transform 1 0 2856 0 1 2970
box -8 -3 16 105
use FILL  FILL_283
timestamp 1712622712
transform 1 0 2848 0 1 2970
box -8 -3 16 105
use FILL  FILL_284
timestamp 1712622712
transform 1 0 2824 0 1 2970
box -8 -3 16 105
use FILL  FILL_285
timestamp 1712622712
transform 1 0 2800 0 1 2970
box -8 -3 16 105
use FILL  FILL_286
timestamp 1712622712
transform 1 0 2792 0 1 2970
box -8 -3 16 105
use FILL  FILL_287
timestamp 1712622712
transform 1 0 2784 0 1 2970
box -8 -3 16 105
use FILL  FILL_288
timestamp 1712622712
transform 1 0 2736 0 1 2970
box -8 -3 16 105
use FILL  FILL_289
timestamp 1712622712
transform 1 0 2728 0 1 2970
box -8 -3 16 105
use FILL  FILL_290
timestamp 1712622712
transform 1 0 2720 0 1 2970
box -8 -3 16 105
use FILL  FILL_291
timestamp 1712622712
transform 1 0 2712 0 1 2970
box -8 -3 16 105
use FILL  FILL_292
timestamp 1712622712
transform 1 0 2704 0 1 2970
box -8 -3 16 105
use FILL  FILL_293
timestamp 1712622712
transform 1 0 2696 0 1 2970
box -8 -3 16 105
use FILL  FILL_294
timestamp 1712622712
transform 1 0 2624 0 1 2970
box -8 -3 16 105
use FILL  FILL_295
timestamp 1712622712
transform 1 0 2616 0 1 2970
box -8 -3 16 105
use FILL  FILL_296
timestamp 1712622712
transform 1 0 2608 0 1 2970
box -8 -3 16 105
use FILL  FILL_297
timestamp 1712622712
transform 1 0 2600 0 1 2970
box -8 -3 16 105
use FILL  FILL_298
timestamp 1712622712
transform 1 0 2592 0 1 2970
box -8 -3 16 105
use FILL  FILL_299
timestamp 1712622712
transform 1 0 2584 0 1 2970
box -8 -3 16 105
use FILL  FILL_300
timestamp 1712622712
transform 1 0 2512 0 1 2970
box -8 -3 16 105
use FILL  FILL_301
timestamp 1712622712
transform 1 0 2504 0 1 2970
box -8 -3 16 105
use FILL  FILL_302
timestamp 1712622712
transform 1 0 2496 0 1 2970
box -8 -3 16 105
use FILL  FILL_303
timestamp 1712622712
transform 1 0 2488 0 1 2970
box -8 -3 16 105
use FILL  FILL_304
timestamp 1712622712
transform 1 0 2456 0 1 2970
box -8 -3 16 105
use FILL  FILL_305
timestamp 1712622712
transform 1 0 2416 0 1 2970
box -8 -3 16 105
use FILL  FILL_306
timestamp 1712622712
transform 1 0 2408 0 1 2970
box -8 -3 16 105
use FILL  FILL_307
timestamp 1712622712
transform 1 0 2384 0 1 2970
box -8 -3 16 105
use FILL  FILL_308
timestamp 1712622712
transform 1 0 2376 0 1 2970
box -8 -3 16 105
use FILL  FILL_309
timestamp 1712622712
transform 1 0 2368 0 1 2970
box -8 -3 16 105
use FILL  FILL_310
timestamp 1712622712
transform 1 0 2360 0 1 2970
box -8 -3 16 105
use FILL  FILL_311
timestamp 1712622712
transform 1 0 2288 0 1 2970
box -8 -3 16 105
use FILL  FILL_312
timestamp 1712622712
transform 1 0 2280 0 1 2970
box -8 -3 16 105
use FILL  FILL_313
timestamp 1712622712
transform 1 0 2272 0 1 2970
box -8 -3 16 105
use FILL  FILL_314
timestamp 1712622712
transform 1 0 2240 0 1 2970
box -8 -3 16 105
use FILL  FILL_315
timestamp 1712622712
transform 1 0 2232 0 1 2970
box -8 -3 16 105
use FILL  FILL_316
timestamp 1712622712
transform 1 0 2168 0 1 2970
box -8 -3 16 105
use FILL  FILL_317
timestamp 1712622712
transform 1 0 2160 0 1 2970
box -8 -3 16 105
use FILL  FILL_318
timestamp 1712622712
transform 1 0 2152 0 1 2970
box -8 -3 16 105
use FILL  FILL_319
timestamp 1712622712
transform 1 0 2088 0 1 2970
box -8 -3 16 105
use FILL  FILL_320
timestamp 1712622712
transform 1 0 2080 0 1 2970
box -8 -3 16 105
use FILL  FILL_321
timestamp 1712622712
transform 1 0 2072 0 1 2970
box -8 -3 16 105
use FILL  FILL_322
timestamp 1712622712
transform 1 0 2032 0 1 2970
box -8 -3 16 105
use FILL  FILL_323
timestamp 1712622712
transform 1 0 1984 0 1 2970
box -8 -3 16 105
use FILL  FILL_324
timestamp 1712622712
transform 1 0 1976 0 1 2970
box -8 -3 16 105
use FILL  FILL_325
timestamp 1712622712
transform 1 0 1952 0 1 2970
box -8 -3 16 105
use FILL  FILL_326
timestamp 1712622712
transform 1 0 1912 0 1 2970
box -8 -3 16 105
use FILL  FILL_327
timestamp 1712622712
transform 1 0 1904 0 1 2970
box -8 -3 16 105
use FILL  FILL_328
timestamp 1712622712
transform 1 0 1856 0 1 2970
box -8 -3 16 105
use FILL  FILL_329
timestamp 1712622712
transform 1 0 1848 0 1 2970
box -8 -3 16 105
use FILL  FILL_330
timestamp 1712622712
transform 1 0 1800 0 1 2970
box -8 -3 16 105
use FILL  FILL_331
timestamp 1712622712
transform 1 0 1792 0 1 2970
box -8 -3 16 105
use FILL  FILL_332
timestamp 1712622712
transform 1 0 1784 0 1 2970
box -8 -3 16 105
use FILL  FILL_333
timestamp 1712622712
transform 1 0 1736 0 1 2970
box -8 -3 16 105
use FILL  FILL_334
timestamp 1712622712
transform 1 0 1728 0 1 2970
box -8 -3 16 105
use FILL  FILL_335
timestamp 1712622712
transform 1 0 1720 0 1 2970
box -8 -3 16 105
use FILL  FILL_336
timestamp 1712622712
transform 1 0 1680 0 1 2970
box -8 -3 16 105
use FILL  FILL_337
timestamp 1712622712
transform 1 0 1632 0 1 2970
box -8 -3 16 105
use FILL  FILL_338
timestamp 1712622712
transform 1 0 1624 0 1 2970
box -8 -3 16 105
use FILL  FILL_339
timestamp 1712622712
transform 1 0 1616 0 1 2970
box -8 -3 16 105
use FILL  FILL_340
timestamp 1712622712
transform 1 0 1608 0 1 2970
box -8 -3 16 105
use FILL  FILL_341
timestamp 1712622712
transform 1 0 1560 0 1 2970
box -8 -3 16 105
use FILL  FILL_342
timestamp 1712622712
transform 1 0 1552 0 1 2970
box -8 -3 16 105
use FILL  FILL_343
timestamp 1712622712
transform 1 0 1504 0 1 2970
box -8 -3 16 105
use FILL  FILL_344
timestamp 1712622712
transform 1 0 1496 0 1 2970
box -8 -3 16 105
use FILL  FILL_345
timestamp 1712622712
transform 1 0 1488 0 1 2970
box -8 -3 16 105
use FILL  FILL_346
timestamp 1712622712
transform 1 0 1440 0 1 2970
box -8 -3 16 105
use FILL  FILL_347
timestamp 1712622712
transform 1 0 1432 0 1 2970
box -8 -3 16 105
use FILL  FILL_348
timestamp 1712622712
transform 1 0 1392 0 1 2970
box -8 -3 16 105
use FILL  FILL_349
timestamp 1712622712
transform 1 0 1384 0 1 2970
box -8 -3 16 105
use FILL  FILL_350
timestamp 1712622712
transform 1 0 1376 0 1 2970
box -8 -3 16 105
use FILL  FILL_351
timestamp 1712622712
transform 1 0 1328 0 1 2970
box -8 -3 16 105
use FILL  FILL_352
timestamp 1712622712
transform 1 0 1320 0 1 2970
box -8 -3 16 105
use FILL  FILL_353
timestamp 1712622712
transform 1 0 1312 0 1 2970
box -8 -3 16 105
use FILL  FILL_354
timestamp 1712622712
transform 1 0 1272 0 1 2970
box -8 -3 16 105
use FILL  FILL_355
timestamp 1712622712
transform 1 0 1264 0 1 2970
box -8 -3 16 105
use FILL  FILL_356
timestamp 1712622712
transform 1 0 1224 0 1 2970
box -8 -3 16 105
use FILL  FILL_357
timestamp 1712622712
transform 1 0 1216 0 1 2970
box -8 -3 16 105
use FILL  FILL_358
timestamp 1712622712
transform 1 0 1168 0 1 2970
box -8 -3 16 105
use FILL  FILL_359
timestamp 1712622712
transform 1 0 1160 0 1 2970
box -8 -3 16 105
use FILL  FILL_360
timestamp 1712622712
transform 1 0 1112 0 1 2970
box -8 -3 16 105
use FILL  FILL_361
timestamp 1712622712
transform 1 0 1104 0 1 2970
box -8 -3 16 105
use FILL  FILL_362
timestamp 1712622712
transform 1 0 1096 0 1 2970
box -8 -3 16 105
use FILL  FILL_363
timestamp 1712622712
transform 1 0 1072 0 1 2970
box -8 -3 16 105
use FILL  FILL_364
timestamp 1712622712
transform 1 0 1064 0 1 2970
box -8 -3 16 105
use FILL  FILL_365
timestamp 1712622712
transform 1 0 1056 0 1 2970
box -8 -3 16 105
use FILL  FILL_366
timestamp 1712622712
transform 1 0 1000 0 1 2970
box -8 -3 16 105
use FILL  FILL_367
timestamp 1712622712
transform 1 0 992 0 1 2970
box -8 -3 16 105
use FILL  FILL_368
timestamp 1712622712
transform 1 0 984 0 1 2970
box -8 -3 16 105
use FILL  FILL_369
timestamp 1712622712
transform 1 0 936 0 1 2970
box -8 -3 16 105
use FILL  FILL_370
timestamp 1712622712
transform 1 0 928 0 1 2970
box -8 -3 16 105
use FILL  FILL_371
timestamp 1712622712
transform 1 0 920 0 1 2970
box -8 -3 16 105
use FILL  FILL_372
timestamp 1712622712
transform 1 0 864 0 1 2970
box -8 -3 16 105
use FILL  FILL_373
timestamp 1712622712
transform 1 0 856 0 1 2970
box -8 -3 16 105
use FILL  FILL_374
timestamp 1712622712
transform 1 0 816 0 1 2970
box -8 -3 16 105
use FILL  FILL_375
timestamp 1712622712
transform 1 0 808 0 1 2970
box -8 -3 16 105
use FILL  FILL_376
timestamp 1712622712
transform 1 0 776 0 1 2970
box -8 -3 16 105
use FILL  FILL_377
timestamp 1712622712
transform 1 0 752 0 1 2970
box -8 -3 16 105
use FILL  FILL_378
timestamp 1712622712
transform 1 0 744 0 1 2970
box -8 -3 16 105
use FILL  FILL_379
timestamp 1712622712
transform 1 0 696 0 1 2970
box -8 -3 16 105
use FILL  FILL_380
timestamp 1712622712
transform 1 0 688 0 1 2970
box -8 -3 16 105
use FILL  FILL_381
timestamp 1712622712
transform 1 0 680 0 1 2970
box -8 -3 16 105
use FILL  FILL_382
timestamp 1712622712
transform 1 0 624 0 1 2970
box -8 -3 16 105
use FILL  FILL_383
timestamp 1712622712
transform 1 0 616 0 1 2970
box -8 -3 16 105
use FILL  FILL_384
timestamp 1712622712
transform 1 0 608 0 1 2970
box -8 -3 16 105
use FILL  FILL_385
timestamp 1712622712
transform 1 0 552 0 1 2970
box -8 -3 16 105
use FILL  FILL_386
timestamp 1712622712
transform 1 0 504 0 1 2970
box -8 -3 16 105
use FILL  FILL_387
timestamp 1712622712
transform 1 0 496 0 1 2970
box -8 -3 16 105
use FILL  FILL_388
timestamp 1712622712
transform 1 0 488 0 1 2970
box -8 -3 16 105
use FILL  FILL_389
timestamp 1712622712
transform 1 0 440 0 1 2970
box -8 -3 16 105
use FILL  FILL_390
timestamp 1712622712
transform 1 0 432 0 1 2970
box -8 -3 16 105
use FILL  FILL_391
timestamp 1712622712
transform 1 0 376 0 1 2970
box -8 -3 16 105
use FILL  FILL_392
timestamp 1712622712
transform 1 0 368 0 1 2970
box -8 -3 16 105
use FILL  FILL_393
timestamp 1712622712
transform 1 0 360 0 1 2970
box -8 -3 16 105
use FILL  FILL_394
timestamp 1712622712
transform 1 0 256 0 1 2970
box -8 -3 16 105
use FILL  FILL_395
timestamp 1712622712
transform 1 0 248 0 1 2970
box -8 -3 16 105
use FILL  FILL_396
timestamp 1712622712
transform 1 0 240 0 1 2970
box -8 -3 16 105
use FILL  FILL_397
timestamp 1712622712
transform 1 0 184 0 1 2970
box -8 -3 16 105
use FILL  FILL_398
timestamp 1712622712
transform 1 0 176 0 1 2970
box -8 -3 16 105
use FILL  FILL_399
timestamp 1712622712
transform 1 0 72 0 1 2970
box -8 -3 16 105
use FILL  FILL_400
timestamp 1712622712
transform 1 0 3328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_401
timestamp 1712622712
transform 1 0 3224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_402
timestamp 1712622712
transform 1 0 3216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_403
timestamp 1712622712
transform 1 0 3192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_404
timestamp 1712622712
transform 1 0 3184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_405
timestamp 1712622712
transform 1 0 3176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_406
timestamp 1712622712
transform 1 0 3112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_407
timestamp 1712622712
transform 1 0 3104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_408
timestamp 1712622712
transform 1 0 3096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_409
timestamp 1712622712
transform 1 0 3088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_410
timestamp 1712622712
transform 1 0 3080 0 -1 2970
box -8 -3 16 105
use FILL  FILL_411
timestamp 1712622712
transform 1 0 2992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_412
timestamp 1712622712
transform 1 0 2984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_413
timestamp 1712622712
transform 1 0 2880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_414
timestamp 1712622712
transform 1 0 2872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_415
timestamp 1712622712
transform 1 0 2832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_416
timestamp 1712622712
transform 1 0 2824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_417
timestamp 1712622712
transform 1 0 2704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_418
timestamp 1712622712
transform 1 0 2696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_419
timestamp 1712622712
transform 1 0 2592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_420
timestamp 1712622712
transform 1 0 2584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_421
timestamp 1712622712
transform 1 0 2576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_422
timestamp 1712622712
transform 1 0 2504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_423
timestamp 1712622712
transform 1 0 2496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_424
timestamp 1712622712
transform 1 0 2488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_425
timestamp 1712622712
transform 1 0 2480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_426
timestamp 1712622712
transform 1 0 2472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_427
timestamp 1712622712
transform 1 0 2392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_428
timestamp 1712622712
transform 1 0 2384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_429
timestamp 1712622712
transform 1 0 2360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_430
timestamp 1712622712
transform 1 0 2352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_431
timestamp 1712622712
transform 1 0 2344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_432
timestamp 1712622712
transform 1 0 2264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_433
timestamp 1712622712
transform 1 0 2256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_434
timestamp 1712622712
transform 1 0 2248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_435
timestamp 1712622712
transform 1 0 2240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_436
timestamp 1712622712
transform 1 0 2168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_437
timestamp 1712622712
transform 1 0 2160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_438
timestamp 1712622712
transform 1 0 2152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_439
timestamp 1712622712
transform 1 0 2048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_440
timestamp 1712622712
transform 1 0 2040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_441
timestamp 1712622712
transform 1 0 2032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_442
timestamp 1712622712
transform 1 0 1976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_443
timestamp 1712622712
transform 1 0 1968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_444
timestamp 1712622712
transform 1 0 1960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_445
timestamp 1712622712
transform 1 0 1912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_446
timestamp 1712622712
transform 1 0 1872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_447
timestamp 1712622712
transform 1 0 1864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_448
timestamp 1712622712
transform 1 0 1856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_449
timestamp 1712622712
transform 1 0 1832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_450
timestamp 1712622712
transform 1 0 1784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_451
timestamp 1712622712
transform 1 0 1776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_452
timestamp 1712622712
transform 1 0 1736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_453
timestamp 1712622712
transform 1 0 1728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_454
timestamp 1712622712
transform 1 0 1680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_455
timestamp 1712622712
transform 1 0 1672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_456
timestamp 1712622712
transform 1 0 1664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_457
timestamp 1712622712
transform 1 0 1656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_458
timestamp 1712622712
transform 1 0 1576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_459
timestamp 1712622712
transform 1 0 1568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_460
timestamp 1712622712
transform 1 0 1344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_461
timestamp 1712622712
transform 1 0 1296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_462
timestamp 1712622712
transform 1 0 1288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_463
timestamp 1712622712
transform 1 0 1280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_464
timestamp 1712622712
transform 1 0 1200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_465
timestamp 1712622712
transform 1 0 1192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_466
timestamp 1712622712
transform 1 0 1184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_467
timestamp 1712622712
transform 1 0 1048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_468
timestamp 1712622712
transform 1 0 1040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_469
timestamp 1712622712
transform 1 0 1032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_470
timestamp 1712622712
transform 1 0 1008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_471
timestamp 1712622712
transform 1 0 944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_472
timestamp 1712622712
transform 1 0 936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_473
timestamp 1712622712
transform 1 0 928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_474
timestamp 1712622712
transform 1 0 888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_475
timestamp 1712622712
transform 1 0 824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_476
timestamp 1712622712
transform 1 0 816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_477
timestamp 1712622712
transform 1 0 808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_478
timestamp 1712622712
transform 1 0 728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_479
timestamp 1712622712
transform 1 0 720 0 -1 2970
box -8 -3 16 105
use FILL  FILL_480
timestamp 1712622712
transform 1 0 712 0 -1 2970
box -8 -3 16 105
use FILL  FILL_481
timestamp 1712622712
transform 1 0 664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_482
timestamp 1712622712
transform 1 0 616 0 -1 2970
box -8 -3 16 105
use FILL  FILL_483
timestamp 1712622712
transform 1 0 608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_484
timestamp 1712622712
transform 1 0 600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_485
timestamp 1712622712
transform 1 0 592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_486
timestamp 1712622712
transform 1 0 536 0 -1 2970
box -8 -3 16 105
use FILL  FILL_487
timestamp 1712622712
transform 1 0 528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_488
timestamp 1712622712
transform 1 0 520 0 -1 2970
box -8 -3 16 105
use FILL  FILL_489
timestamp 1712622712
transform 1 0 416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_490
timestamp 1712622712
transform 1 0 408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_491
timestamp 1712622712
transform 1 0 400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_492
timestamp 1712622712
transform 1 0 320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_493
timestamp 1712622712
transform 1 0 312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_494
timestamp 1712622712
transform 1 0 304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_495
timestamp 1712622712
transform 1 0 296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_496
timestamp 1712622712
transform 1 0 192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_497
timestamp 1712622712
transform 1 0 184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_498
timestamp 1712622712
transform 1 0 176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_499
timestamp 1712622712
transform 1 0 168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_500
timestamp 1712622712
transform 1 0 112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_501
timestamp 1712622712
transform 1 0 80 0 -1 2970
box -8 -3 16 105
use FILL  FILL_502
timestamp 1712622712
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_503
timestamp 1712622712
transform 1 0 3328 0 1 2770
box -8 -3 16 105
use FILL  FILL_504
timestamp 1712622712
transform 1 0 3320 0 1 2770
box -8 -3 16 105
use FILL  FILL_505
timestamp 1712622712
transform 1 0 3264 0 1 2770
box -8 -3 16 105
use FILL  FILL_506
timestamp 1712622712
transform 1 0 3256 0 1 2770
box -8 -3 16 105
use FILL  FILL_507
timestamp 1712622712
transform 1 0 3248 0 1 2770
box -8 -3 16 105
use FILL  FILL_508
timestamp 1712622712
transform 1 0 3208 0 1 2770
box -8 -3 16 105
use FILL  FILL_509
timestamp 1712622712
transform 1 0 3200 0 1 2770
box -8 -3 16 105
use FILL  FILL_510
timestamp 1712622712
transform 1 0 3192 0 1 2770
box -8 -3 16 105
use FILL  FILL_511
timestamp 1712622712
transform 1 0 3184 0 1 2770
box -8 -3 16 105
use FILL  FILL_512
timestamp 1712622712
transform 1 0 3176 0 1 2770
box -8 -3 16 105
use FILL  FILL_513
timestamp 1712622712
transform 1 0 3112 0 1 2770
box -8 -3 16 105
use FILL  FILL_514
timestamp 1712622712
transform 1 0 3104 0 1 2770
box -8 -3 16 105
use FILL  FILL_515
timestamp 1712622712
transform 1 0 3096 0 1 2770
box -8 -3 16 105
use FILL  FILL_516
timestamp 1712622712
transform 1 0 3088 0 1 2770
box -8 -3 16 105
use FILL  FILL_517
timestamp 1712622712
transform 1 0 3024 0 1 2770
box -8 -3 16 105
use FILL  FILL_518
timestamp 1712622712
transform 1 0 3016 0 1 2770
box -8 -3 16 105
use FILL  FILL_519
timestamp 1712622712
transform 1 0 3008 0 1 2770
box -8 -3 16 105
use FILL  FILL_520
timestamp 1712622712
transform 1 0 3000 0 1 2770
box -8 -3 16 105
use FILL  FILL_521
timestamp 1712622712
transform 1 0 2904 0 1 2770
box -8 -3 16 105
use FILL  FILL_522
timestamp 1712622712
transform 1 0 2800 0 1 2770
box -8 -3 16 105
use FILL  FILL_523
timestamp 1712622712
transform 1 0 2792 0 1 2770
box -8 -3 16 105
use FILL  FILL_524
timestamp 1712622712
transform 1 0 2784 0 1 2770
box -8 -3 16 105
use FILL  FILL_525
timestamp 1712622712
transform 1 0 2696 0 1 2770
box -8 -3 16 105
use FILL  FILL_526
timestamp 1712622712
transform 1 0 2688 0 1 2770
box -8 -3 16 105
use FILL  FILL_527
timestamp 1712622712
transform 1 0 2584 0 1 2770
box -8 -3 16 105
use FILL  FILL_528
timestamp 1712622712
transform 1 0 2576 0 1 2770
box -8 -3 16 105
use FILL  FILL_529
timestamp 1712622712
transform 1 0 2520 0 1 2770
box -8 -3 16 105
use FILL  FILL_530
timestamp 1712622712
transform 1 0 2512 0 1 2770
box -8 -3 16 105
use FILL  FILL_531
timestamp 1712622712
transform 1 0 2368 0 1 2770
box -8 -3 16 105
use FILL  FILL_532
timestamp 1712622712
transform 1 0 2360 0 1 2770
box -8 -3 16 105
use FILL  FILL_533
timestamp 1712622712
transform 1 0 2352 0 1 2770
box -8 -3 16 105
use FILL  FILL_534
timestamp 1712622712
transform 1 0 2120 0 1 2770
box -8 -3 16 105
use FILL  FILL_535
timestamp 1712622712
transform 1 0 1968 0 1 2770
box -8 -3 16 105
use FILL  FILL_536
timestamp 1712622712
transform 1 0 1960 0 1 2770
box -8 -3 16 105
use FILL  FILL_537
timestamp 1712622712
transform 1 0 1824 0 1 2770
box -8 -3 16 105
use FILL  FILL_538
timestamp 1712622712
transform 1 0 1816 0 1 2770
box -8 -3 16 105
use FILL  FILL_539
timestamp 1712622712
transform 1 0 1776 0 1 2770
box -8 -3 16 105
use FILL  FILL_540
timestamp 1712622712
transform 1 0 1672 0 1 2770
box -8 -3 16 105
use FILL  FILL_541
timestamp 1712622712
transform 1 0 1664 0 1 2770
box -8 -3 16 105
use FILL  FILL_542
timestamp 1712622712
transform 1 0 1624 0 1 2770
box -8 -3 16 105
use FILL  FILL_543
timestamp 1712622712
transform 1 0 1616 0 1 2770
box -8 -3 16 105
use FILL  FILL_544
timestamp 1712622712
transform 1 0 1512 0 1 2770
box -8 -3 16 105
use FILL  FILL_545
timestamp 1712622712
transform 1 0 1488 0 1 2770
box -8 -3 16 105
use FILL  FILL_546
timestamp 1712622712
transform 1 0 1480 0 1 2770
box -8 -3 16 105
use FILL  FILL_547
timestamp 1712622712
transform 1 0 1472 0 1 2770
box -8 -3 16 105
use FILL  FILL_548
timestamp 1712622712
transform 1 0 1368 0 1 2770
box -8 -3 16 105
use FILL  FILL_549
timestamp 1712622712
transform 1 0 1360 0 1 2770
box -8 -3 16 105
use FILL  FILL_550
timestamp 1712622712
transform 1 0 1304 0 1 2770
box -8 -3 16 105
use FILL  FILL_551
timestamp 1712622712
transform 1 0 1296 0 1 2770
box -8 -3 16 105
use FILL  FILL_552
timestamp 1712622712
transform 1 0 1192 0 1 2770
box -8 -3 16 105
use FILL  FILL_553
timestamp 1712622712
transform 1 0 1184 0 1 2770
box -8 -3 16 105
use FILL  FILL_554
timestamp 1712622712
transform 1 0 1176 0 1 2770
box -8 -3 16 105
use FILL  FILL_555
timestamp 1712622712
transform 1 0 1120 0 1 2770
box -8 -3 16 105
use FILL  FILL_556
timestamp 1712622712
transform 1 0 1112 0 1 2770
box -8 -3 16 105
use FILL  FILL_557
timestamp 1712622712
transform 1 0 1008 0 1 2770
box -8 -3 16 105
use FILL  FILL_558
timestamp 1712622712
transform 1 0 1000 0 1 2770
box -8 -3 16 105
use FILL  FILL_559
timestamp 1712622712
transform 1 0 992 0 1 2770
box -8 -3 16 105
use FILL  FILL_560
timestamp 1712622712
transform 1 0 984 0 1 2770
box -8 -3 16 105
use FILL  FILL_561
timestamp 1712622712
transform 1 0 920 0 1 2770
box -8 -3 16 105
use FILL  FILL_562
timestamp 1712622712
transform 1 0 912 0 1 2770
box -8 -3 16 105
use FILL  FILL_563
timestamp 1712622712
transform 1 0 904 0 1 2770
box -8 -3 16 105
use FILL  FILL_564
timestamp 1712622712
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_565
timestamp 1712622712
transform 1 0 888 0 1 2770
box -8 -3 16 105
use FILL  FILL_566
timestamp 1712622712
transform 1 0 848 0 1 2770
box -8 -3 16 105
use FILL  FILL_567
timestamp 1712622712
transform 1 0 816 0 1 2770
box -8 -3 16 105
use FILL  FILL_568
timestamp 1712622712
transform 1 0 808 0 1 2770
box -8 -3 16 105
use FILL  FILL_569
timestamp 1712622712
transform 1 0 800 0 1 2770
box -8 -3 16 105
use FILL  FILL_570
timestamp 1712622712
transform 1 0 792 0 1 2770
box -8 -3 16 105
use FILL  FILL_571
timestamp 1712622712
transform 1 0 752 0 1 2770
box -8 -3 16 105
use FILL  FILL_572
timestamp 1712622712
transform 1 0 744 0 1 2770
box -8 -3 16 105
use FILL  FILL_573
timestamp 1712622712
transform 1 0 704 0 1 2770
box -8 -3 16 105
use FILL  FILL_574
timestamp 1712622712
transform 1 0 696 0 1 2770
box -8 -3 16 105
use FILL  FILL_575
timestamp 1712622712
transform 1 0 688 0 1 2770
box -8 -3 16 105
use FILL  FILL_576
timestamp 1712622712
transform 1 0 640 0 1 2770
box -8 -3 16 105
use FILL  FILL_577
timestamp 1712622712
transform 1 0 632 0 1 2770
box -8 -3 16 105
use FILL  FILL_578
timestamp 1712622712
transform 1 0 624 0 1 2770
box -8 -3 16 105
use FILL  FILL_579
timestamp 1712622712
transform 1 0 576 0 1 2770
box -8 -3 16 105
use FILL  FILL_580
timestamp 1712622712
transform 1 0 568 0 1 2770
box -8 -3 16 105
use FILL  FILL_581
timestamp 1712622712
transform 1 0 528 0 1 2770
box -8 -3 16 105
use FILL  FILL_582
timestamp 1712622712
transform 1 0 520 0 1 2770
box -8 -3 16 105
use FILL  FILL_583
timestamp 1712622712
transform 1 0 512 0 1 2770
box -8 -3 16 105
use FILL  FILL_584
timestamp 1712622712
transform 1 0 504 0 1 2770
box -8 -3 16 105
use FILL  FILL_585
timestamp 1712622712
transform 1 0 496 0 1 2770
box -8 -3 16 105
use FILL  FILL_586
timestamp 1712622712
transform 1 0 416 0 1 2770
box -8 -3 16 105
use FILL  FILL_587
timestamp 1712622712
transform 1 0 408 0 1 2770
box -8 -3 16 105
use FILL  FILL_588
timestamp 1712622712
transform 1 0 400 0 1 2770
box -8 -3 16 105
use FILL  FILL_589
timestamp 1712622712
transform 1 0 296 0 1 2770
box -8 -3 16 105
use FILL  FILL_590
timestamp 1712622712
transform 1 0 288 0 1 2770
box -8 -3 16 105
use FILL  FILL_591
timestamp 1712622712
transform 1 0 184 0 1 2770
box -8 -3 16 105
use FILL  FILL_592
timestamp 1712622712
transform 1 0 176 0 1 2770
box -8 -3 16 105
use FILL  FILL_593
timestamp 1712622712
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_594
timestamp 1712622712
transform 1 0 3424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_595
timestamp 1712622712
transform 1 0 3320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_596
timestamp 1712622712
transform 1 0 3312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_597
timestamp 1712622712
transform 1 0 3304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_598
timestamp 1712622712
transform 1 0 3240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_599
timestamp 1712622712
transform 1 0 3232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_600
timestamp 1712622712
transform 1 0 3224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_601
timestamp 1712622712
transform 1 0 3216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_602
timestamp 1712622712
transform 1 0 3208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_603
timestamp 1712622712
transform 1 0 3200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_604
timestamp 1712622712
transform 1 0 3192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_605
timestamp 1712622712
transform 1 0 3120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_606
timestamp 1712622712
transform 1 0 3112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_607
timestamp 1712622712
transform 1 0 3104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_608
timestamp 1712622712
transform 1 0 3096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_609
timestamp 1712622712
transform 1 0 3088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_610
timestamp 1712622712
transform 1 0 2984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_611
timestamp 1712622712
transform 1 0 2976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_612
timestamp 1712622712
transform 1 0 2872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_613
timestamp 1712622712
transform 1 0 2864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_614
timestamp 1712622712
transform 1 0 2856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_615
timestamp 1712622712
transform 1 0 2848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_616
timestamp 1712622712
transform 1 0 2840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_617
timestamp 1712622712
transform 1 0 2792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_618
timestamp 1712622712
transform 1 0 2784 0 -1 2770
box -8 -3 16 105
use FILL  FILL_619
timestamp 1712622712
transform 1 0 2776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_620
timestamp 1712622712
transform 1 0 2744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_621
timestamp 1712622712
transform 1 0 2736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_622
timestamp 1712622712
transform 1 0 2728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_623
timestamp 1712622712
transform 1 0 2680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_624
timestamp 1712622712
transform 1 0 2672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_625
timestamp 1712622712
transform 1 0 2664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_626
timestamp 1712622712
transform 1 0 2560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_627
timestamp 1712622712
transform 1 0 2552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_628
timestamp 1712622712
transform 1 0 2448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_629
timestamp 1712622712
transform 1 0 2440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_630
timestamp 1712622712
transform 1 0 2336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_631
timestamp 1712622712
transform 1 0 2304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_632
timestamp 1712622712
transform 1 0 2200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_633
timestamp 1712622712
transform 1 0 2192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_634
timestamp 1712622712
transform 1 0 2184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_635
timestamp 1712622712
transform 1 0 2128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_636
timestamp 1712622712
transform 1 0 2120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_637
timestamp 1712622712
transform 1 0 2112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_638
timestamp 1712622712
transform 1 0 2056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_639
timestamp 1712622712
transform 1 0 2048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_640
timestamp 1712622712
transform 1 0 2040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_641
timestamp 1712622712
transform 1 0 2008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_642
timestamp 1712622712
transform 1 0 2000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_643
timestamp 1712622712
transform 1 0 1992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_644
timestamp 1712622712
transform 1 0 1888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_645
timestamp 1712622712
transform 1 0 1880 0 -1 2770
box -8 -3 16 105
use FILL  FILL_646
timestamp 1712622712
transform 1 0 1872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_647
timestamp 1712622712
transform 1 0 1864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_648
timestamp 1712622712
transform 1 0 1816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_649
timestamp 1712622712
transform 1 0 1808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_650
timestamp 1712622712
transform 1 0 1800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_651
timestamp 1712622712
transform 1 0 1752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_652
timestamp 1712622712
transform 1 0 1744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_653
timestamp 1712622712
transform 1 0 1736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_654
timestamp 1712622712
transform 1 0 1712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_655
timestamp 1712622712
transform 1 0 1704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_656
timestamp 1712622712
transform 1 0 1696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_657
timestamp 1712622712
transform 1 0 1688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_658
timestamp 1712622712
transform 1 0 1640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_659
timestamp 1712622712
transform 1 0 1632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_660
timestamp 1712622712
transform 1 0 1624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_661
timestamp 1712622712
transform 1 0 1600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_662
timestamp 1712622712
transform 1 0 1592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_663
timestamp 1712622712
transform 1 0 1584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_664
timestamp 1712622712
transform 1 0 1536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_665
timestamp 1712622712
transform 1 0 1528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_666
timestamp 1712622712
transform 1 0 1520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_667
timestamp 1712622712
transform 1 0 1512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_668
timestamp 1712622712
transform 1 0 1408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_669
timestamp 1712622712
transform 1 0 1400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_670
timestamp 1712622712
transform 1 0 1392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_671
timestamp 1712622712
transform 1 0 1384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_672
timestamp 1712622712
transform 1 0 1376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_673
timestamp 1712622712
transform 1 0 1368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_674
timestamp 1712622712
transform 1 0 1312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_675
timestamp 1712622712
transform 1 0 1304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_676
timestamp 1712622712
transform 1 0 1296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_677
timestamp 1712622712
transform 1 0 1288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_678
timestamp 1712622712
transform 1 0 1280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_679
timestamp 1712622712
transform 1 0 1272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_680
timestamp 1712622712
transform 1 0 1264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_681
timestamp 1712622712
transform 1 0 1216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_682
timestamp 1712622712
transform 1 0 1208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_683
timestamp 1712622712
transform 1 0 1200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_684
timestamp 1712622712
transform 1 0 1192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_685
timestamp 1712622712
transform 1 0 1184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_686
timestamp 1712622712
transform 1 0 1176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_687
timestamp 1712622712
transform 1 0 1168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_688
timestamp 1712622712
transform 1 0 1160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_689
timestamp 1712622712
transform 1 0 1104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_690
timestamp 1712622712
transform 1 0 1080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_691
timestamp 1712622712
transform 1 0 1072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_692
timestamp 1712622712
transform 1 0 1064 0 -1 2770
box -8 -3 16 105
use FILL  FILL_693
timestamp 1712622712
transform 1 0 1056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_694
timestamp 1712622712
transform 1 0 1048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_695
timestamp 1712622712
transform 1 0 944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_696
timestamp 1712622712
transform 1 0 936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_697
timestamp 1712622712
transform 1 0 928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_698
timestamp 1712622712
transform 1 0 920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_699
timestamp 1712622712
transform 1 0 872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_700
timestamp 1712622712
transform 1 0 864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_701
timestamp 1712622712
transform 1 0 760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_702
timestamp 1712622712
transform 1 0 752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_703
timestamp 1712622712
transform 1 0 744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_704
timestamp 1712622712
transform 1 0 736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_705
timestamp 1712622712
transform 1 0 728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_706
timestamp 1712622712
transform 1 0 680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_707
timestamp 1712622712
transform 1 0 672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_708
timestamp 1712622712
transform 1 0 664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_709
timestamp 1712622712
transform 1 0 640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_710
timestamp 1712622712
transform 1 0 632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_711
timestamp 1712622712
transform 1 0 624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_712
timestamp 1712622712
transform 1 0 576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_713
timestamp 1712622712
transform 1 0 568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_714
timestamp 1712622712
transform 1 0 560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_715
timestamp 1712622712
transform 1 0 456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_716
timestamp 1712622712
transform 1 0 448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_717
timestamp 1712622712
transform 1 0 344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_718
timestamp 1712622712
transform 1 0 336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_719
timestamp 1712622712
transform 1 0 328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_720
timestamp 1712622712
transform 1 0 224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_721
timestamp 1712622712
transform 1 0 216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_722
timestamp 1712622712
transform 1 0 208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_723
timestamp 1712622712
transform 1 0 104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_724
timestamp 1712622712
transform 1 0 96 0 -1 2770
box -8 -3 16 105
use FILL  FILL_725
timestamp 1712622712
transform 1 0 88 0 -1 2770
box -8 -3 16 105
use FILL  FILL_726
timestamp 1712622712
transform 1 0 80 0 -1 2770
box -8 -3 16 105
use FILL  FILL_727
timestamp 1712622712
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_728
timestamp 1712622712
transform 1 0 3424 0 1 2570
box -8 -3 16 105
use FILL  FILL_729
timestamp 1712622712
transform 1 0 3392 0 1 2570
box -8 -3 16 105
use FILL  FILL_730
timestamp 1712622712
transform 1 0 3384 0 1 2570
box -8 -3 16 105
use FILL  FILL_731
timestamp 1712622712
transform 1 0 3376 0 1 2570
box -8 -3 16 105
use FILL  FILL_732
timestamp 1712622712
transform 1 0 3368 0 1 2570
box -8 -3 16 105
use FILL  FILL_733
timestamp 1712622712
transform 1 0 3320 0 1 2570
box -8 -3 16 105
use FILL  FILL_734
timestamp 1712622712
transform 1 0 3312 0 1 2570
box -8 -3 16 105
use FILL  FILL_735
timestamp 1712622712
transform 1 0 3304 0 1 2570
box -8 -3 16 105
use FILL  FILL_736
timestamp 1712622712
transform 1 0 3272 0 1 2570
box -8 -3 16 105
use FILL  FILL_737
timestamp 1712622712
transform 1 0 3264 0 1 2570
box -8 -3 16 105
use FILL  FILL_738
timestamp 1712622712
transform 1 0 3256 0 1 2570
box -8 -3 16 105
use FILL  FILL_739
timestamp 1712622712
transform 1 0 3248 0 1 2570
box -8 -3 16 105
use FILL  FILL_740
timestamp 1712622712
transform 1 0 3200 0 1 2570
box -8 -3 16 105
use FILL  FILL_741
timestamp 1712622712
transform 1 0 3192 0 1 2570
box -8 -3 16 105
use FILL  FILL_742
timestamp 1712622712
transform 1 0 3184 0 1 2570
box -8 -3 16 105
use FILL  FILL_743
timestamp 1712622712
transform 1 0 3176 0 1 2570
box -8 -3 16 105
use FILL  FILL_744
timestamp 1712622712
transform 1 0 3168 0 1 2570
box -8 -3 16 105
use FILL  FILL_745
timestamp 1712622712
transform 1 0 3160 0 1 2570
box -8 -3 16 105
use FILL  FILL_746
timestamp 1712622712
transform 1 0 3120 0 1 2570
box -8 -3 16 105
use FILL  FILL_747
timestamp 1712622712
transform 1 0 3112 0 1 2570
box -8 -3 16 105
use FILL  FILL_748
timestamp 1712622712
transform 1 0 3104 0 1 2570
box -8 -3 16 105
use FILL  FILL_749
timestamp 1712622712
transform 1 0 3064 0 1 2570
box -8 -3 16 105
use FILL  FILL_750
timestamp 1712622712
transform 1 0 3056 0 1 2570
box -8 -3 16 105
use FILL  FILL_751
timestamp 1712622712
transform 1 0 3048 0 1 2570
box -8 -3 16 105
use FILL  FILL_752
timestamp 1712622712
transform 1 0 3040 0 1 2570
box -8 -3 16 105
use FILL  FILL_753
timestamp 1712622712
transform 1 0 2936 0 1 2570
box -8 -3 16 105
use FILL  FILL_754
timestamp 1712622712
transform 1 0 2928 0 1 2570
box -8 -3 16 105
use FILL  FILL_755
timestamp 1712622712
transform 1 0 2920 0 1 2570
box -8 -3 16 105
use FILL  FILL_756
timestamp 1712622712
transform 1 0 2872 0 1 2570
box -8 -3 16 105
use FILL  FILL_757
timestamp 1712622712
transform 1 0 2864 0 1 2570
box -8 -3 16 105
use FILL  FILL_758
timestamp 1712622712
transform 1 0 2856 0 1 2570
box -8 -3 16 105
use FILL  FILL_759
timestamp 1712622712
transform 1 0 2848 0 1 2570
box -8 -3 16 105
use FILL  FILL_760
timestamp 1712622712
transform 1 0 2744 0 1 2570
box -8 -3 16 105
use FILL  FILL_761
timestamp 1712622712
transform 1 0 2736 0 1 2570
box -8 -3 16 105
use FILL  FILL_762
timestamp 1712622712
transform 1 0 2632 0 1 2570
box -8 -3 16 105
use FILL  FILL_763
timestamp 1712622712
transform 1 0 2624 0 1 2570
box -8 -3 16 105
use FILL  FILL_764
timestamp 1712622712
transform 1 0 2616 0 1 2570
box -8 -3 16 105
use FILL  FILL_765
timestamp 1712622712
transform 1 0 2512 0 1 2570
box -8 -3 16 105
use FILL  FILL_766
timestamp 1712622712
transform 1 0 2504 0 1 2570
box -8 -3 16 105
use FILL  FILL_767
timestamp 1712622712
transform 1 0 2496 0 1 2570
box -8 -3 16 105
use FILL  FILL_768
timestamp 1712622712
transform 1 0 2488 0 1 2570
box -8 -3 16 105
use FILL  FILL_769
timestamp 1712622712
transform 1 0 2440 0 1 2570
box -8 -3 16 105
use FILL  FILL_770
timestamp 1712622712
transform 1 0 2432 0 1 2570
box -8 -3 16 105
use FILL  FILL_771
timestamp 1712622712
transform 1 0 2424 0 1 2570
box -8 -3 16 105
use FILL  FILL_772
timestamp 1712622712
transform 1 0 2376 0 1 2570
box -8 -3 16 105
use FILL  FILL_773
timestamp 1712622712
transform 1 0 2368 0 1 2570
box -8 -3 16 105
use FILL  FILL_774
timestamp 1712622712
transform 1 0 2360 0 1 2570
box -8 -3 16 105
use FILL  FILL_775
timestamp 1712622712
transform 1 0 2352 0 1 2570
box -8 -3 16 105
use FILL  FILL_776
timestamp 1712622712
transform 1 0 2344 0 1 2570
box -8 -3 16 105
use FILL  FILL_777
timestamp 1712622712
transform 1 0 2264 0 1 2570
box -8 -3 16 105
use FILL  FILL_778
timestamp 1712622712
transform 1 0 2256 0 1 2570
box -8 -3 16 105
use FILL  FILL_779
timestamp 1712622712
transform 1 0 2248 0 1 2570
box -8 -3 16 105
use FILL  FILL_780
timestamp 1712622712
transform 1 0 2240 0 1 2570
box -8 -3 16 105
use FILL  FILL_781
timestamp 1712622712
transform 1 0 2136 0 1 2570
box -8 -3 16 105
use FILL  FILL_782
timestamp 1712622712
transform 1 0 2128 0 1 2570
box -8 -3 16 105
use FILL  FILL_783
timestamp 1712622712
transform 1 0 2120 0 1 2570
box -8 -3 16 105
use FILL  FILL_784
timestamp 1712622712
transform 1 0 2016 0 1 2570
box -8 -3 16 105
use FILL  FILL_785
timestamp 1712622712
transform 1 0 2008 0 1 2570
box -8 -3 16 105
use FILL  FILL_786
timestamp 1712622712
transform 1 0 2000 0 1 2570
box -8 -3 16 105
use FILL  FILL_787
timestamp 1712622712
transform 1 0 1896 0 1 2570
box -8 -3 16 105
use FILL  FILL_788
timestamp 1712622712
transform 1 0 1888 0 1 2570
box -8 -3 16 105
use FILL  FILL_789
timestamp 1712622712
transform 1 0 1784 0 1 2570
box -8 -3 16 105
use FILL  FILL_790
timestamp 1712622712
transform 1 0 1776 0 1 2570
box -8 -3 16 105
use FILL  FILL_791
timestamp 1712622712
transform 1 0 1672 0 1 2570
box -8 -3 16 105
use FILL  FILL_792
timestamp 1712622712
transform 1 0 1664 0 1 2570
box -8 -3 16 105
use FILL  FILL_793
timestamp 1712622712
transform 1 0 1560 0 1 2570
box -8 -3 16 105
use FILL  FILL_794
timestamp 1712622712
transform 1 0 1552 0 1 2570
box -8 -3 16 105
use FILL  FILL_795
timestamp 1712622712
transform 1 0 1544 0 1 2570
box -8 -3 16 105
use FILL  FILL_796
timestamp 1712622712
transform 1 0 1536 0 1 2570
box -8 -3 16 105
use FILL  FILL_797
timestamp 1712622712
transform 1 0 1488 0 1 2570
box -8 -3 16 105
use FILL  FILL_798
timestamp 1712622712
transform 1 0 1480 0 1 2570
box -8 -3 16 105
use FILL  FILL_799
timestamp 1712622712
transform 1 0 1432 0 1 2570
box -8 -3 16 105
use FILL  FILL_800
timestamp 1712622712
transform 1 0 1424 0 1 2570
box -8 -3 16 105
use FILL  FILL_801
timestamp 1712622712
transform 1 0 1416 0 1 2570
box -8 -3 16 105
use FILL  FILL_802
timestamp 1712622712
transform 1 0 1312 0 1 2570
box -8 -3 16 105
use FILL  FILL_803
timestamp 1712622712
transform 1 0 1304 0 1 2570
box -8 -3 16 105
use FILL  FILL_804
timestamp 1712622712
transform 1 0 1200 0 1 2570
box -8 -3 16 105
use FILL  FILL_805
timestamp 1712622712
transform 1 0 1096 0 1 2570
box -8 -3 16 105
use FILL  FILL_806
timestamp 1712622712
transform 1 0 1088 0 1 2570
box -8 -3 16 105
use FILL  FILL_807
timestamp 1712622712
transform 1 0 984 0 1 2570
box -8 -3 16 105
use FILL  FILL_808
timestamp 1712622712
transform 1 0 880 0 1 2570
box -8 -3 16 105
use FILL  FILL_809
timestamp 1712622712
transform 1 0 776 0 1 2570
box -8 -3 16 105
use FILL  FILL_810
timestamp 1712622712
transform 1 0 768 0 1 2570
box -8 -3 16 105
use FILL  FILL_811
timestamp 1712622712
transform 1 0 664 0 1 2570
box -8 -3 16 105
use FILL  FILL_812
timestamp 1712622712
transform 1 0 560 0 1 2570
box -8 -3 16 105
use FILL  FILL_813
timestamp 1712622712
transform 1 0 552 0 1 2570
box -8 -3 16 105
use FILL  FILL_814
timestamp 1712622712
transform 1 0 544 0 1 2570
box -8 -3 16 105
use FILL  FILL_815
timestamp 1712622712
transform 1 0 488 0 1 2570
box -8 -3 16 105
use FILL  FILL_816
timestamp 1712622712
transform 1 0 480 0 1 2570
box -8 -3 16 105
use FILL  FILL_817
timestamp 1712622712
transform 1 0 472 0 1 2570
box -8 -3 16 105
use FILL  FILL_818
timestamp 1712622712
transform 1 0 464 0 1 2570
box -8 -3 16 105
use FILL  FILL_819
timestamp 1712622712
transform 1 0 360 0 1 2570
box -8 -3 16 105
use FILL  FILL_820
timestamp 1712622712
transform 1 0 352 0 1 2570
box -8 -3 16 105
use FILL  FILL_821
timestamp 1712622712
transform 1 0 344 0 1 2570
box -8 -3 16 105
use FILL  FILL_822
timestamp 1712622712
transform 1 0 336 0 1 2570
box -8 -3 16 105
use FILL  FILL_823
timestamp 1712622712
transform 1 0 288 0 1 2570
box -8 -3 16 105
use FILL  FILL_824
timestamp 1712622712
transform 1 0 280 0 1 2570
box -8 -3 16 105
use FILL  FILL_825
timestamp 1712622712
transform 1 0 272 0 1 2570
box -8 -3 16 105
use FILL  FILL_826
timestamp 1712622712
transform 1 0 224 0 1 2570
box -8 -3 16 105
use FILL  FILL_827
timestamp 1712622712
transform 1 0 216 0 1 2570
box -8 -3 16 105
use FILL  FILL_828
timestamp 1712622712
transform 1 0 208 0 1 2570
box -8 -3 16 105
use FILL  FILL_829
timestamp 1712622712
transform 1 0 200 0 1 2570
box -8 -3 16 105
use FILL  FILL_830
timestamp 1712622712
transform 1 0 192 0 1 2570
box -8 -3 16 105
use FILL  FILL_831
timestamp 1712622712
transform 1 0 144 0 1 2570
box -8 -3 16 105
use FILL  FILL_832
timestamp 1712622712
transform 1 0 136 0 1 2570
box -8 -3 16 105
use FILL  FILL_833
timestamp 1712622712
transform 1 0 128 0 1 2570
box -8 -3 16 105
use FILL  FILL_834
timestamp 1712622712
transform 1 0 80 0 1 2570
box -8 -3 16 105
use FILL  FILL_835
timestamp 1712622712
transform 1 0 72 0 1 2570
box -8 -3 16 105
use FILL  FILL_836
timestamp 1712622712
transform 1 0 3328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_837
timestamp 1712622712
transform 1 0 3224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_838
timestamp 1712622712
transform 1 0 3216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_839
timestamp 1712622712
transform 1 0 3208 0 -1 2570
box -8 -3 16 105
use FILL  FILL_840
timestamp 1712622712
transform 1 0 3200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_841
timestamp 1712622712
transform 1 0 3128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_842
timestamp 1712622712
transform 1 0 3120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_843
timestamp 1712622712
transform 1 0 3112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_844
timestamp 1712622712
transform 1 0 3104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_845
timestamp 1712622712
transform 1 0 3096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_846
timestamp 1712622712
transform 1 0 3088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_847
timestamp 1712622712
transform 1 0 3016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_848
timestamp 1712622712
transform 1 0 3008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_849
timestamp 1712622712
transform 1 0 3000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_850
timestamp 1712622712
transform 1 0 2992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_851
timestamp 1712622712
transform 1 0 2888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_852
timestamp 1712622712
transform 1 0 2880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_853
timestamp 1712622712
transform 1 0 2872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_854
timestamp 1712622712
transform 1 0 2864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_855
timestamp 1712622712
transform 1 0 2816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_856
timestamp 1712622712
transform 1 0 2808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_857
timestamp 1712622712
transform 1 0 2800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_858
timestamp 1712622712
transform 1 0 2792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_859
timestamp 1712622712
transform 1 0 2784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_860
timestamp 1712622712
transform 1 0 2736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_861
timestamp 1712622712
transform 1 0 2728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_862
timestamp 1712622712
transform 1 0 2720 0 -1 2570
box -8 -3 16 105
use FILL  FILL_863
timestamp 1712622712
transform 1 0 2712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_864
timestamp 1712622712
transform 1 0 2704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_865
timestamp 1712622712
transform 1 0 2656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_866
timestamp 1712622712
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_867
timestamp 1712622712
transform 1 0 2640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_868
timestamp 1712622712
transform 1 0 2632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_869
timestamp 1712622712
transform 1 0 2584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_870
timestamp 1712622712
transform 1 0 2576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_871
timestamp 1712622712
transform 1 0 2568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_872
timestamp 1712622712
transform 1 0 2560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_873
timestamp 1712622712
transform 1 0 2552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_874
timestamp 1712622712
transform 1 0 2544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_875
timestamp 1712622712
transform 1 0 2496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_876
timestamp 1712622712
transform 1 0 2488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_877
timestamp 1712622712
transform 1 0 2480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_878
timestamp 1712622712
transform 1 0 2472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_879
timestamp 1712622712
transform 1 0 2376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_880
timestamp 1712622712
transform 1 0 2368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_881
timestamp 1712622712
transform 1 0 2360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_882
timestamp 1712622712
transform 1 0 2352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_883
timestamp 1712622712
transform 1 0 2304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_884
timestamp 1712622712
transform 1 0 2296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_885
timestamp 1712622712
transform 1 0 2288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_886
timestamp 1712622712
transform 1 0 2256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_887
timestamp 1712622712
transform 1 0 2208 0 -1 2570
box -8 -3 16 105
use FILL  FILL_888
timestamp 1712622712
transform 1 0 2200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_889
timestamp 1712622712
transform 1 0 2192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_890
timestamp 1712622712
transform 1 0 2184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_891
timestamp 1712622712
transform 1 0 2176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_892
timestamp 1712622712
transform 1 0 2104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_893
timestamp 1712622712
transform 1 0 2096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_894
timestamp 1712622712
transform 1 0 2088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_895
timestamp 1712622712
transform 1 0 2080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_896
timestamp 1712622712
transform 1 0 2072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_897
timestamp 1712622712
transform 1 0 2024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_898
timestamp 1712622712
transform 1 0 2016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_899
timestamp 1712622712
transform 1 0 2008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_900
timestamp 1712622712
transform 1 0 2000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_901
timestamp 1712622712
transform 1 0 1952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_902
timestamp 1712622712
transform 1 0 1944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_903
timestamp 1712622712
transform 1 0 1936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_904
timestamp 1712622712
transform 1 0 1880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_905
timestamp 1712622712
transform 1 0 1872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_906
timestamp 1712622712
transform 1 0 1824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_907
timestamp 1712622712
transform 1 0 1816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_908
timestamp 1712622712
transform 1 0 1808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_909
timestamp 1712622712
transform 1 0 1800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_910
timestamp 1712622712
transform 1 0 1792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_911
timestamp 1712622712
transform 1 0 1744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_912
timestamp 1712622712
transform 1 0 1712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_913
timestamp 1712622712
transform 1 0 1704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_914
timestamp 1712622712
transform 1 0 1696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_915
timestamp 1712622712
transform 1 0 1648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_916
timestamp 1712622712
transform 1 0 1640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_917
timestamp 1712622712
transform 1 0 1632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_918
timestamp 1712622712
transform 1 0 1624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_919
timestamp 1712622712
transform 1 0 1576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_920
timestamp 1712622712
transform 1 0 1568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_921
timestamp 1712622712
transform 1 0 1560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_922
timestamp 1712622712
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_923
timestamp 1712622712
transform 1 0 1352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_924
timestamp 1712622712
transform 1 0 1248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_925
timestamp 1712622712
transform 1 0 1240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_926
timestamp 1712622712
transform 1 0 1192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_927
timestamp 1712622712
transform 1 0 1184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_928
timestamp 1712622712
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_929
timestamp 1712622712
transform 1 0 1128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_930
timestamp 1712622712
transform 1 0 1120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_931
timestamp 1712622712
transform 1 0 1016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_932
timestamp 1712622712
transform 1 0 1008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_933
timestamp 1712622712
transform 1 0 1000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_934
timestamp 1712622712
transform 1 0 992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_935
timestamp 1712622712
transform 1 0 944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_936
timestamp 1712622712
transform 1 0 936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_937
timestamp 1712622712
transform 1 0 928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_938
timestamp 1712622712
transform 1 0 920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_939
timestamp 1712622712
transform 1 0 912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_940
timestamp 1712622712
transform 1 0 864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_941
timestamp 1712622712
transform 1 0 856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_942
timestamp 1712622712
transform 1 0 848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_943
timestamp 1712622712
transform 1 0 840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_944
timestamp 1712622712
transform 1 0 792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_945
timestamp 1712622712
transform 1 0 784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_946
timestamp 1712622712
transform 1 0 776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_947
timestamp 1712622712
transform 1 0 768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_948
timestamp 1712622712
transform 1 0 760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_949
timestamp 1712622712
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_950
timestamp 1712622712
transform 1 0 704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_951
timestamp 1712622712
transform 1 0 696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_952
timestamp 1712622712
transform 1 0 688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_953
timestamp 1712622712
transform 1 0 680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_954
timestamp 1712622712
transform 1 0 672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_955
timestamp 1712622712
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_956
timestamp 1712622712
transform 1 0 656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_957
timestamp 1712622712
transform 1 0 608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_958
timestamp 1712622712
transform 1 0 600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_959
timestamp 1712622712
transform 1 0 592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_960
timestamp 1712622712
transform 1 0 584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_961
timestamp 1712622712
transform 1 0 560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_962
timestamp 1712622712
transform 1 0 552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_963
timestamp 1712622712
transform 1 0 544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_964
timestamp 1712622712
transform 1 0 536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_965
timestamp 1712622712
transform 1 0 488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_966
timestamp 1712622712
transform 1 0 480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_967
timestamp 1712622712
transform 1 0 472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_968
timestamp 1712622712
transform 1 0 464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_969
timestamp 1712622712
transform 1 0 456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_970
timestamp 1712622712
transform 1 0 448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_971
timestamp 1712622712
transform 1 0 400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_972
timestamp 1712622712
transform 1 0 392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_973
timestamp 1712622712
transform 1 0 384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_974
timestamp 1712622712
transform 1 0 376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_975
timestamp 1712622712
transform 1 0 368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_976
timestamp 1712622712
transform 1 0 320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_977
timestamp 1712622712
transform 1 0 312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_978
timestamp 1712622712
transform 1 0 304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_979
timestamp 1712622712
transform 1 0 296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_980
timestamp 1712622712
transform 1 0 192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_981
timestamp 1712622712
transform 1 0 184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_982
timestamp 1712622712
transform 1 0 80 0 -1 2570
box -8 -3 16 105
use FILL  FILL_983
timestamp 1712622712
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_984
timestamp 1712622712
transform 1 0 3424 0 1 2370
box -8 -3 16 105
use FILL  FILL_985
timestamp 1712622712
transform 1 0 3384 0 1 2370
box -8 -3 16 105
use FILL  FILL_986
timestamp 1712622712
transform 1 0 3376 0 1 2370
box -8 -3 16 105
use FILL  FILL_987
timestamp 1712622712
transform 1 0 3368 0 1 2370
box -8 -3 16 105
use FILL  FILL_988
timestamp 1712622712
transform 1 0 3360 0 1 2370
box -8 -3 16 105
use FILL  FILL_989
timestamp 1712622712
transform 1 0 3320 0 1 2370
box -8 -3 16 105
use FILL  FILL_990
timestamp 1712622712
transform 1 0 3272 0 1 2370
box -8 -3 16 105
use FILL  FILL_991
timestamp 1712622712
transform 1 0 3264 0 1 2370
box -8 -3 16 105
use FILL  FILL_992
timestamp 1712622712
transform 1 0 3256 0 1 2370
box -8 -3 16 105
use FILL  FILL_993
timestamp 1712622712
transform 1 0 3152 0 1 2370
box -8 -3 16 105
use FILL  FILL_994
timestamp 1712622712
transform 1 0 2952 0 1 2370
box -8 -3 16 105
use FILL  FILL_995
timestamp 1712622712
transform 1 0 2656 0 1 2370
box -8 -3 16 105
use FILL  FILL_996
timestamp 1712622712
transform 1 0 2360 0 1 2370
box -8 -3 16 105
use FILL  FILL_997
timestamp 1712622712
transform 1 0 2064 0 1 2370
box -8 -3 16 105
use FILL  FILL_998
timestamp 1712622712
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use FILL  FILL_999
timestamp 1712622712
transform 1 0 1760 0 1 2370
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1712622712
transform 1 0 1728 0 1 2370
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1712622712
transform 1 0 1624 0 1 2370
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1712622712
transform 1 0 1616 0 1 2370
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1712622712
transform 1 0 1512 0 1 2370
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1712622712
transform 1 0 1504 0 1 2370
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1712622712
transform 1 0 1496 0 1 2370
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1712622712
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1712622712
transform 1 0 1448 0 1 2370
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1712622712
transform 1 0 1440 0 1 2370
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1712622712
transform 1 0 1400 0 1 2370
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1712622712
transform 1 0 1392 0 1 2370
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1712622712
transform 1 0 1384 0 1 2370
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1712622712
transform 1 0 1376 0 1 2370
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1712622712
transform 1 0 1368 0 1 2370
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1712622712
transform 1 0 1328 0 1 2370
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1712622712
transform 1 0 1320 0 1 2370
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1712622712
transform 1 0 1280 0 1 2370
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1712622712
transform 1 0 1272 0 1 2370
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1712622712
transform 1 0 1264 0 1 2370
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1712622712
transform 1 0 1256 0 1 2370
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1712622712
transform 1 0 1248 0 1 2370
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1712622712
transform 1 0 1144 0 1 2370
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1712622712
transform 1 0 1136 0 1 2370
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1712622712
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1712622712
transform 1 0 1088 0 1 2370
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1712622712
transform 1 0 1080 0 1 2370
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1712622712
transform 1 0 1072 0 1 2370
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1712622712
transform 1 0 1064 0 1 2370
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1712622712
transform 1 0 960 0 1 2370
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1712622712
transform 1 0 952 0 1 2370
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1712622712
transform 1 0 848 0 1 2370
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1712622712
transform 1 0 840 0 1 2370
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1712622712
transform 1 0 736 0 1 2370
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1712622712
transform 1 0 728 0 1 2370
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1712622712
transform 1 0 624 0 1 2370
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1712622712
transform 1 0 520 0 1 2370
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1712622712
transform 1 0 512 0 1 2370
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1712622712
transform 1 0 408 0 1 2370
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1712622712
transform 1 0 400 0 1 2370
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1712622712
transform 1 0 296 0 1 2370
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1712622712
transform 1 0 288 0 1 2370
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1712622712
transform 1 0 184 0 1 2370
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1712622712
transform 1 0 176 0 1 2370
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1712622712
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1712622712
transform 1 0 3424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1712622712
transform 1 0 3416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1712622712
transform 1 0 3408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1712622712
transform 1 0 3352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1712622712
transform 1 0 3344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1712622712
transform 1 0 3336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1712622712
transform 1 0 3328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1712622712
transform 1 0 3320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1712622712
transform 1 0 3264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1712622712
transform 1 0 3232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1712622712
transform 1 0 3224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1712622712
transform 1 0 3216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1712622712
transform 1 0 3208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1712622712
transform 1 0 3200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1712622712
transform 1 0 3192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1712622712
transform 1 0 3136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1712622712
transform 1 0 3128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1712622712
transform 1 0 3120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1712622712
transform 1 0 3112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1712622712
transform 1 0 3080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1712622712
transform 1 0 3040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1712622712
transform 1 0 3032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1712622712
transform 1 0 3024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1712622712
transform 1 0 3016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1712622712
transform 1 0 2976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1712622712
transform 1 0 2968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1712622712
transform 1 0 2960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1712622712
transform 1 0 2952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1712622712
transform 1 0 2928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1712622712
transform 1 0 2888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1712622712
transform 1 0 2880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1712622712
transform 1 0 2872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1712622712
transform 1 0 2864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1712622712
transform 1 0 2856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1712622712
transform 1 0 2816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1712622712
transform 1 0 2808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1712622712
transform 1 0 2800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1712622712
transform 1 0 2792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1712622712
transform 1 0 2752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1712622712
transform 1 0 2744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1712622712
transform 1 0 2736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1712622712
transform 1 0 2728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1712622712
transform 1 0 2688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1712622712
transform 1 0 2680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1712622712
transform 1 0 2648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1712622712
transform 1 0 2640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1712622712
transform 1 0 2632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1712622712
transform 1 0 2592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1712622712
transform 1 0 2584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1712622712
transform 1 0 2576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1712622712
transform 1 0 2536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1712622712
transform 1 0 2528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1712622712
transform 1 0 2520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1712622712
transform 1 0 2512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1712622712
transform 1 0 2472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1712622712
transform 1 0 2464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1712622712
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1712622712
transform 1 0 2416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1712622712
transform 1 0 2408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1712622712
transform 1 0 2400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1712622712
transform 1 0 2392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1712622712
transform 1 0 2352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1712622712
transform 1 0 2344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1712622712
transform 1 0 2336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1712622712
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1712622712
transform 1 0 2288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1712622712
transform 1 0 2280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1712622712
transform 1 0 2272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1712622712
transform 1 0 2264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1712622712
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1712622712
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1712622712
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1712622712
transform 1 0 2168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1712622712
transform 1 0 2160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1712622712
transform 1 0 2152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1712622712
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1712622712
transform 1 0 2136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1712622712
transform 1 0 2096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1712622712
transform 1 0 2088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1712622712
transform 1 0 2080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1712622712
transform 1 0 2072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1712622712
transform 1 0 2032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1712622712
transform 1 0 2024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1712622712
transform 1 0 2016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1712622712
transform 1 0 2008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1712622712
transform 1 0 1968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1712622712
transform 1 0 1960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1712622712
transform 1 0 1952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1712622712
transform 1 0 1944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1712622712
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1712622712
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1712622712
transform 1 0 1888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1712622712
transform 1 0 1880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1712622712
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1712622712
transform 1 0 1832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1712622712
transform 1 0 1824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1712622712
transform 1 0 1816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1712622712
transform 1 0 1776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1712622712
transform 1 0 1768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1712622712
transform 1 0 1736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1712622712
transform 1 0 1704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1712622712
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1712622712
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1712622712
transform 1 0 1648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1712622712
transform 1 0 1640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1712622712
transform 1 0 1608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1712622712
transform 1 0 1600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1712622712
transform 1 0 1560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1712622712
transform 1 0 1552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1712622712
transform 1 0 1544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1712622712
transform 1 0 1536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1712622712
transform 1 0 1528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1712622712
transform 1 0 1488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1712622712
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1712622712
transform 1 0 1440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1712622712
transform 1 0 1432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1712622712
transform 1 0 1424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1712622712
transform 1 0 1416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1712622712
transform 1 0 1376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1712622712
transform 1 0 1368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1712622712
transform 1 0 1360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1712622712
transform 1 0 1320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1712622712
transform 1 0 1312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1712622712
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1712622712
transform 1 0 1296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1712622712
transform 1 0 1288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1712622712
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1712622712
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1712622712
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1712622712
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1712622712
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1712622712
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1712622712
transform 1 0 1168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1712622712
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1712622712
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1712622712
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1712622712
transform 1 0 1056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1712622712
transform 1 0 1048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1712622712
transform 1 0 1040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1712622712
transform 1 0 1032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1712622712
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1712622712
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1712622712
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1712622712
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1712622712
transform 1 0 944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1712622712
transform 1 0 936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1712622712
transform 1 0 928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1712622712
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1712622712
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1712622712
transform 1 0 872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1712622712
transform 1 0 832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1712622712
transform 1 0 824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1712622712
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1712622712
transform 1 0 776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1712622712
transform 1 0 768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1712622712
transform 1 0 760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1712622712
transform 1 0 752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1712622712
transform 1 0 712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1712622712
transform 1 0 704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1712622712
transform 1 0 696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1712622712
transform 1 0 688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1712622712
transform 1 0 648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1712622712
transform 1 0 640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1712622712
transform 1 0 632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1712622712
transform 1 0 624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1712622712
transform 1 0 616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1712622712
transform 1 0 576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1712622712
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1712622712
transform 1 0 560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1712622712
transform 1 0 552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1712622712
transform 1 0 512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1712622712
transform 1 0 504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1712622712
transform 1 0 496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1712622712
transform 1 0 488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1712622712
transform 1 0 448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1712622712
transform 1 0 440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1712622712
transform 1 0 432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1712622712
transform 1 0 424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1712622712
transform 1 0 384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1712622712
transform 1 0 376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1712622712
transform 1 0 368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1712622712
transform 1 0 360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1712622712
transform 1 0 352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1712622712
transform 1 0 344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1712622712
transform 1 0 304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1712622712
transform 1 0 296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1712622712
transform 1 0 256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1712622712
transform 1 0 248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1712622712
transform 1 0 240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1712622712
transform 1 0 232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1712622712
transform 1 0 224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1712622712
transform 1 0 120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1712622712
transform 1 0 112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1712622712
transform 1 0 104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1712622712
transform 1 0 96 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1712622712
transform 1 0 88 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1712622712
transform 1 0 80 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1712622712
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1712622712
transform 1 0 3424 0 1 2170
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1712622712
transform 1 0 3416 0 1 2170
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1712622712
transform 1 0 3384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1712622712
transform 1 0 3376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1712622712
transform 1 0 3368 0 1 2170
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1712622712
transform 1 0 3304 0 1 2170
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1712622712
transform 1 0 3296 0 1 2170
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1712622712
transform 1 0 3288 0 1 2170
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1712622712
transform 1 0 3280 0 1 2170
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1712622712
transform 1 0 3208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1712622712
transform 1 0 3200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1712622712
transform 1 0 3176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1712622712
transform 1 0 3168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1712622712
transform 1 0 3160 0 1 2170
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1712622712
transform 1 0 3152 0 1 2170
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1712622712
transform 1 0 3088 0 1 2170
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1712622712
transform 1 0 3080 0 1 2170
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1712622712
transform 1 0 3072 0 1 2170
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1712622712
transform 1 0 3064 0 1 2170
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1712622712
transform 1 0 3056 0 1 2170
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1712622712
transform 1 0 3016 0 1 2170
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1712622712
transform 1 0 3008 0 1 2170
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1712622712
transform 1 0 2968 0 1 2170
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1712622712
transform 1 0 2960 0 1 2170
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1712622712
transform 1 0 2952 0 1 2170
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1712622712
transform 1 0 2944 0 1 2170
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1712622712
transform 1 0 2936 0 1 2170
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1712622712
transform 1 0 2896 0 1 2170
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1712622712
transform 1 0 2888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1712622712
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1712622712
transform 1 0 2840 0 1 2170
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1712622712
transform 1 0 2832 0 1 2170
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1712622712
transform 1 0 2824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1712622712
transform 1 0 2816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1712622712
transform 1 0 2752 0 1 2170
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1712622712
transform 1 0 2744 0 1 2170
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1712622712
transform 1 0 2712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1712622712
transform 1 0 2704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1712622712
transform 1 0 2696 0 1 2170
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1712622712
transform 1 0 2688 0 1 2170
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1712622712
transform 1 0 2632 0 1 2170
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1712622712
transform 1 0 2624 0 1 2170
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1712622712
transform 1 0 2616 0 1 2170
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1712622712
transform 1 0 2608 0 1 2170
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1712622712
transform 1 0 2600 0 1 2170
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1712622712
transform 1 0 2536 0 1 2170
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1712622712
transform 1 0 2528 0 1 2170
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1712622712
transform 1 0 2520 0 1 2170
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1712622712
transform 1 0 2512 0 1 2170
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1712622712
transform 1 0 2504 0 1 2170
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1712622712
transform 1 0 2496 0 1 2170
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1712622712
transform 1 0 2448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1712622712
transform 1 0 2440 0 1 2170
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1712622712
transform 1 0 2432 0 1 2170
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1712622712
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1712622712
transform 1 0 2392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1712622712
transform 1 0 2384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1712622712
transform 1 0 2376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1712622712
transform 1 0 2328 0 1 2170
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1712622712
transform 1 0 2320 0 1 2170
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1712622712
transform 1 0 2312 0 1 2170
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1712622712
transform 1 0 2304 0 1 2170
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1712622712
transform 1 0 2272 0 1 2170
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1712622712
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1712622712
transform 1 0 2216 0 1 2170
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1712622712
transform 1 0 2208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1712622712
transform 1 0 2200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1712622712
transform 1 0 2192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1712622712
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1712622712
transform 1 0 2136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1712622712
transform 1 0 2128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1712622712
transform 1 0 2120 0 1 2170
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1712622712
transform 1 0 2088 0 1 2170
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1712622712
transform 1 0 2080 0 1 2170
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1712622712
transform 1 0 2072 0 1 2170
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1712622712
transform 1 0 2024 0 1 2170
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1712622712
transform 1 0 2016 0 1 2170
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1712622712
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1712622712
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1712622712
transform 1 0 1992 0 1 2170
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1712622712
transform 1 0 1960 0 1 2170
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1712622712
transform 1 0 1952 0 1 2170
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1712622712
transform 1 0 1904 0 1 2170
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1712622712
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1712622712
transform 1 0 1888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1712622712
transform 1 0 1880 0 1 2170
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1712622712
transform 1 0 1872 0 1 2170
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1712622712
transform 1 0 1832 0 1 2170
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1712622712
transform 1 0 1824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1712622712
transform 1 0 1792 0 1 2170
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1712622712
transform 1 0 1784 0 1 2170
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1712622712
transform 1 0 1776 0 1 2170
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1712622712
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1712622712
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1712622712
transform 1 0 1712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1712622712
transform 1 0 1688 0 1 2170
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1712622712
transform 1 0 1680 0 1 2170
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1712622712
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1712622712
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1712622712
transform 1 0 1656 0 1 2170
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1712622712
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1712622712
transform 1 0 1584 0 1 2170
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1712622712
transform 1 0 1576 0 1 2170
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1712622712
transform 1 0 1568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1712622712
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1712622712
transform 1 0 1504 0 1 2170
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1712622712
transform 1 0 1496 0 1 2170
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1712622712
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1712622712
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1712622712
transform 1 0 1472 0 1 2170
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1712622712
transform 1 0 1448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1712622712
transform 1 0 1400 0 1 2170
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1712622712
transform 1 0 1392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1712622712
transform 1 0 1384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1712622712
transform 1 0 1376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1712622712
transform 1 0 1344 0 1 2170
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1712622712
transform 1 0 1304 0 1 2170
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1712622712
transform 1 0 1296 0 1 2170
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1712622712
transform 1 0 1288 0 1 2170
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1712622712
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1712622712
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1712622712
transform 1 0 1240 0 1 2170
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1712622712
transform 1 0 1192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1712622712
transform 1 0 1184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1712622712
transform 1 0 1176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1712622712
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1712622712
transform 1 0 1128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1712622712
transform 1 0 1120 0 1 2170
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1712622712
transform 1 0 1088 0 1 2170
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1712622712
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1712622712
transform 1 0 1072 0 1 2170
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1712622712
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1712622712
transform 1 0 1024 0 1 2170
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1712622712
transform 1 0 984 0 1 2170
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1712622712
transform 1 0 976 0 1 2170
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1712622712
transform 1 0 968 0 1 2170
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1712622712
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1712622712
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1712622712
transform 1 0 904 0 1 2170
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1712622712
transform 1 0 896 0 1 2170
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1712622712
transform 1 0 856 0 1 2170
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1712622712
transform 1 0 832 0 1 2170
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1712622712
transform 1 0 824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1712622712
transform 1 0 816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1712622712
transform 1 0 808 0 1 2170
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1712622712
transform 1 0 776 0 1 2170
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1712622712
transform 1 0 768 0 1 2170
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1712622712
transform 1 0 760 0 1 2170
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1712622712
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1712622712
transform 1 0 704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1712622712
transform 1 0 696 0 1 2170
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1712622712
transform 1 0 688 0 1 2170
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1712622712
transform 1 0 680 0 1 2170
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1712622712
transform 1 0 632 0 1 2170
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1712622712
transform 1 0 624 0 1 2170
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1712622712
transform 1 0 616 0 1 2170
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1712622712
transform 1 0 608 0 1 2170
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1712622712
transform 1 0 576 0 1 2170
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1712622712
transform 1 0 568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1712622712
transform 1 0 560 0 1 2170
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1712622712
transform 1 0 552 0 1 2170
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1712622712
transform 1 0 504 0 1 2170
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1712622712
transform 1 0 496 0 1 2170
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1712622712
transform 1 0 488 0 1 2170
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1712622712
transform 1 0 480 0 1 2170
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1712622712
transform 1 0 448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1712622712
transform 1 0 440 0 1 2170
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1712622712
transform 1 0 432 0 1 2170
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1712622712
transform 1 0 424 0 1 2170
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1712622712
transform 1 0 384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1712622712
transform 1 0 376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1712622712
transform 1 0 368 0 1 2170
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1712622712
transform 1 0 336 0 1 2170
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1712622712
transform 1 0 328 0 1 2170
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1712622712
transform 1 0 320 0 1 2170
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1712622712
transform 1 0 312 0 1 2170
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1712622712
transform 1 0 272 0 1 2170
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1712622712
transform 1 0 264 0 1 2170
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1712622712
transform 1 0 256 0 1 2170
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1712622712
transform 1 0 248 0 1 2170
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1712622712
transform 1 0 208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1712622712
transform 1 0 200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1712622712
transform 1 0 192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1712622712
transform 1 0 184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1712622712
transform 1 0 176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1712622712
transform 1 0 136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1712622712
transform 1 0 128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1712622712
transform 1 0 120 0 1 2170
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1712622712
transform 1 0 80 0 1 2170
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1712622712
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1712622712
transform 1 0 3424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1712622712
transform 1 0 3416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1712622712
transform 1 0 3344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1712622712
transform 1 0 3336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1712622712
transform 1 0 3272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1712622712
transform 1 0 3264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1712622712
transform 1 0 3240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1712622712
transform 1 0 3232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1712622712
transform 1 0 3224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1712622712
transform 1 0 3200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1712622712
transform 1 0 3136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1712622712
transform 1 0 3128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1712622712
transform 1 0 3120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1712622712
transform 1 0 3072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1712622712
transform 1 0 3064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1712622712
transform 1 0 3024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1712622712
transform 1 0 3016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1712622712
transform 1 0 3008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1712622712
transform 1 0 3000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1712622712
transform 1 0 2928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1712622712
transform 1 0 2920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1712622712
transform 1 0 2912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1712622712
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1712622712
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1712622712
transform 1 0 2816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1712622712
transform 1 0 2808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1712622712
transform 1 0 2800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1712622712
transform 1 0 2760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1712622712
transform 1 0 2752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1712622712
transform 1 0 2744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1712622712
transform 1 0 2680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1712622712
transform 1 0 2672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1712622712
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1712622712
transform 1 0 2656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1712622712
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1712622712
transform 1 0 2584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1712622712
transform 1 0 2576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1712622712
transform 1 0 2568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1712622712
transform 1 0 2512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1712622712
transform 1 0 2504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1712622712
transform 1 0 2496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1712622712
transform 1 0 2488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1712622712
transform 1 0 2440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1712622712
transform 1 0 2432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1712622712
transform 1 0 2392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1712622712
transform 1 0 2384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1712622712
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1712622712
transform 1 0 2352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1712622712
transform 1 0 2304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1712622712
transform 1 0 2296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1712622712
transform 1 0 2288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1712622712
transform 1 0 2280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1712622712
transform 1 0 2232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1712622712
transform 1 0 2224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1712622712
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1712622712
transform 1 0 2168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1712622712
transform 1 0 2160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1712622712
transform 1 0 2152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1712622712
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1712622712
transform 1 0 2112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1712622712
transform 1 0 2072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1712622712
transform 1 0 2064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1712622712
transform 1 0 2056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1712622712
transform 1 0 2048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1712622712
transform 1 0 2000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1712622712
transform 1 0 1992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1712622712
transform 1 0 1984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1712622712
transform 1 0 1952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1712622712
transform 1 0 1944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1712622712
transform 1 0 1936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1712622712
transform 1 0 1928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1712622712
transform 1 0 1896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1712622712
transform 1 0 1848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1712622712
transform 1 0 1840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1712622712
transform 1 0 1832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1712622712
transform 1 0 1824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1712622712
transform 1 0 1816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1712622712
transform 1 0 1808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1712622712
transform 1 0 1736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1712622712
transform 1 0 1728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1712622712
transform 1 0 1720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1712622712
transform 1 0 1712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1712622712
transform 1 0 1704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1712622712
transform 1 0 1656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1712622712
transform 1 0 1616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1712622712
transform 1 0 1608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1712622712
transform 1 0 1600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1712622712
transform 1 0 1592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1712622712
transform 1 0 1544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1712622712
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1712622712
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1712622712
transform 1 0 1480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1712622712
transform 1 0 1472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1712622712
transform 1 0 1464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1712622712
transform 1 0 1416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1712622712
transform 1 0 1408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1712622712
transform 1 0 1400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1712622712
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1712622712
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1712622712
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1712622712
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1712622712
transform 1 0 1304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1712622712
transform 1 0 1296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1712622712
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1712622712
transform 1 0 1224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1712622712
transform 1 0 1216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1712622712
transform 1 0 1168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1712622712
transform 1 0 1160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1712622712
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1712622712
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1712622712
transform 1 0 1096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1712622712
transform 1 0 1088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1712622712
transform 1 0 1040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1712622712
transform 1 0 1016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1712622712
transform 1 0 1008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1712622712
transform 1 0 1000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1712622712
transform 1 0 992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1712622712
transform 1 0 968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1712622712
transform 1 0 912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1712622712
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1712622712
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1712622712
transform 1 0 888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1712622712
transform 1 0 880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1712622712
transform 1 0 872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1712622712
transform 1 0 800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1712622712
transform 1 0 792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1712622712
transform 1 0 784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1712622712
transform 1 0 776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1712622712
transform 1 0 768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1712622712
transform 1 0 760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1712622712
transform 1 0 704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1712622712
transform 1 0 696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1712622712
transform 1 0 688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1712622712
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1712622712
transform 1 0 632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1712622712
transform 1 0 624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1712622712
transform 1 0 616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1712622712
transform 1 0 608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1712622712
transform 1 0 560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1712622712
transform 1 0 552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1712622712
transform 1 0 544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1712622712
transform 1 0 504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1712622712
transform 1 0 496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1712622712
transform 1 0 488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1712622712
transform 1 0 440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1712622712
transform 1 0 432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1712622712
transform 1 0 424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1712622712
transform 1 0 416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1712622712
transform 1 0 368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1712622712
transform 1 0 360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1712622712
transform 1 0 352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1712622712
transform 1 0 344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1712622712
transform 1 0 312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1712622712
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1712622712
transform 1 0 256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1712622712
transform 1 0 248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1712622712
transform 1 0 240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1712622712
transform 1 0 232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1712622712
transform 1 0 224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1712622712
transform 1 0 216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1712622712
transform 1 0 160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1712622712
transform 1 0 152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1712622712
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1712622712
transform 1 0 136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1712622712
transform 1 0 128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1712622712
transform 1 0 80 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1712622712
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1712622712
transform 1 0 3424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1712622712
transform 1 0 3416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1712622712
transform 1 0 3408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1712622712
transform 1 0 3400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1712622712
transform 1 0 3392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1712622712
transform 1 0 3384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1712622712
transform 1 0 3376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1712622712
transform 1 0 3368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1712622712
transform 1 0 3360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1712622712
transform 1 0 3320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1712622712
transform 1 0 3312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1712622712
transform 1 0 3304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1712622712
transform 1 0 3296 0 1 1970
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1712622712
transform 1 0 3288 0 1 1970
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1712622712
transform 1 0 3280 0 1 1970
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1712622712
transform 1 0 3272 0 1 1970
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1712622712
transform 1 0 3224 0 1 1970
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1712622712
transform 1 0 3216 0 1 1970
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1712622712
transform 1 0 3208 0 1 1970
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1712622712
transform 1 0 3200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1712622712
transform 1 0 3160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1712622712
transform 1 0 3152 0 1 1970
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1712622712
transform 1 0 3144 0 1 1970
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1712622712
transform 1 0 3136 0 1 1970
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1712622712
transform 1 0 3128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1712622712
transform 1 0 3080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1712622712
transform 1 0 3072 0 1 1970
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1712622712
transform 1 0 3064 0 1 1970
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1712622712
transform 1 0 3056 0 1 1970
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1712622712
transform 1 0 3016 0 1 1970
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1712622712
transform 1 0 3008 0 1 1970
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1712622712
transform 1 0 3000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1712622712
transform 1 0 2952 0 1 1970
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1712622712
transform 1 0 2944 0 1 1970
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1712622712
transform 1 0 2936 0 1 1970
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1712622712
transform 1 0 2928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1712622712
transform 1 0 2920 0 1 1970
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1712622712
transform 1 0 2880 0 1 1970
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1712622712
transform 1 0 2872 0 1 1970
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1712622712
transform 1 0 2832 0 1 1970
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1712622712
transform 1 0 2824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1712622712
transform 1 0 2816 0 1 1970
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1712622712
transform 1 0 2808 0 1 1970
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1712622712
transform 1 0 2760 0 1 1970
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1712622712
transform 1 0 2752 0 1 1970
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1712622712
transform 1 0 2744 0 1 1970
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1712622712
transform 1 0 2704 0 1 1970
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1712622712
transform 1 0 2696 0 1 1970
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1712622712
transform 1 0 2688 0 1 1970
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1712622712
transform 1 0 2656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1712622712
transform 1 0 2648 0 1 1970
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1712622712
transform 1 0 2640 0 1 1970
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1712622712
transform 1 0 2600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1712622712
transform 1 0 2592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1712622712
transform 1 0 2544 0 1 1970
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1712622712
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1712622712
transform 1 0 2528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1712622712
transform 1 0 2520 0 1 1970
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1712622712
transform 1 0 2512 0 1 1970
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1712622712
transform 1 0 2456 0 1 1970
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1712622712
transform 1 0 2448 0 1 1970
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1712622712
transform 1 0 2440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1712622712
transform 1 0 2432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1712622712
transform 1 0 2424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1712622712
transform 1 0 2416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1712622712
transform 1 0 2360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1712622712
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1712622712
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1712622712
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1712622712
transform 1 0 2304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1712622712
transform 1 0 2224 0 1 1970
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1712622712
transform 1 0 2216 0 1 1970
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1712622712
transform 1 0 2208 0 1 1970
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1712622712
transform 1 0 2200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1712622712
transform 1 0 2192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1712622712
transform 1 0 2128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1712622712
transform 1 0 2120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1712622712
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1712622712
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1712622712
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1712622712
transform 1 0 2048 0 1 1970
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1712622712
transform 1 0 2040 0 1 1970
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1712622712
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1712622712
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1712622712
transform 1 0 1984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1712622712
transform 1 0 1976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1712622712
transform 1 0 1968 0 1 1970
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1712622712
transform 1 0 1904 0 1 1970
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1712622712
transform 1 0 1896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1712622712
transform 1 0 1888 0 1 1970
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1712622712
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1712622712
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1712622712
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1712622712
transform 1 0 1800 0 1 1970
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1712622712
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1712622712
transform 1 0 1752 0 1 1970
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1712622712
transform 1 0 1744 0 1 1970
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1712622712
transform 1 0 1736 0 1 1970
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1712622712
transform 1 0 1688 0 1 1970
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1712622712
transform 1 0 1680 0 1 1970
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1712622712
transform 1 0 1672 0 1 1970
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1712622712
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1712622712
transform 1 0 1624 0 1 1970
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1712622712
transform 1 0 1616 0 1 1970
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1712622712
transform 1 0 1608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1712622712
transform 1 0 1600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1712622712
transform 1 0 1536 0 1 1970
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1712622712
transform 1 0 1528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1712622712
transform 1 0 1520 0 1 1970
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1712622712
transform 1 0 1512 0 1 1970
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1712622712
transform 1 0 1504 0 1 1970
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1712622712
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1712622712
transform 1 0 1488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1712622712
transform 1 0 1424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1712622712
transform 1 0 1416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1712622712
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1712622712
transform 1 0 1376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1712622712
transform 1 0 1368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1712622712
transform 1 0 1360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1712622712
transform 1 0 1304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1712622712
transform 1 0 1296 0 1 1970
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1712622712
transform 1 0 1288 0 1 1970
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1712622712
transform 1 0 1280 0 1 1970
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1712622712
transform 1 0 1272 0 1 1970
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1712622712
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1712622712
transform 1 0 1192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1712622712
transform 1 0 1184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1712622712
transform 1 0 1144 0 1 1970
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1712622712
transform 1 0 1136 0 1 1970
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1712622712
transform 1 0 1128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1712622712
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1712622712
transform 1 0 1056 0 1 1970
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1712622712
transform 1 0 1048 0 1 1970
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1712622712
transform 1 0 1040 0 1 1970
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1712622712
transform 1 0 1032 0 1 1970
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1712622712
transform 1 0 1024 0 1 1970
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1712622712
transform 1 0 1016 0 1 1970
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1712622712
transform 1 0 952 0 1 1970
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1712622712
transform 1 0 944 0 1 1970
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1712622712
transform 1 0 936 0 1 1970
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1712622712
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1712622712
transform 1 0 848 0 1 1970
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1712622712
transform 1 0 840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1712622712
transform 1 0 832 0 1 1970
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1712622712
transform 1 0 824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1712622712
transform 1 0 816 0 1 1970
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1712622712
transform 1 0 768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1712622712
transform 1 0 760 0 1 1970
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1712622712
transform 1 0 728 0 1 1970
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1712622712
transform 1 0 720 0 1 1970
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1712622712
transform 1 0 712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1712622712
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1712622712
transform 1 0 656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1712622712
transform 1 0 648 0 1 1970
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1712622712
transform 1 0 640 0 1 1970
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1712622712
transform 1 0 608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1712622712
transform 1 0 584 0 1 1970
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1712622712
transform 1 0 576 0 1 1970
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1712622712
transform 1 0 568 0 1 1970
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1712622712
transform 1 0 536 0 1 1970
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1712622712
transform 1 0 528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1712622712
transform 1 0 488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1712622712
transform 1 0 480 0 1 1970
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1712622712
transform 1 0 472 0 1 1970
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1712622712
transform 1 0 440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1712622712
transform 1 0 432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1712622712
transform 1 0 392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1712622712
transform 1 0 384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1712622712
transform 1 0 376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1712622712
transform 1 0 344 0 1 1970
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1712622712
transform 1 0 336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1712622712
transform 1 0 328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1712622712
transform 1 0 280 0 1 1970
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1712622712
transform 1 0 272 0 1 1970
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1712622712
transform 1 0 264 0 1 1970
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1712622712
transform 1 0 256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1712622712
transform 1 0 208 0 1 1970
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1712622712
transform 1 0 200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1712622712
transform 1 0 192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1712622712
transform 1 0 160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1712622712
transform 1 0 152 0 1 1970
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1712622712
transform 1 0 144 0 1 1970
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1712622712
transform 1 0 80 0 1 1970
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1712622712
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1712622712
transform 1 0 3304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1712622712
transform 1 0 3248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1712622712
transform 1 0 3240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1712622712
transform 1 0 3232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1712622712
transform 1 0 3136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1712622712
transform 1 0 3128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1712622712
transform 1 0 3120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1712622712
transform 1 0 3112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1712622712
transform 1 0 3072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1712622712
transform 1 0 3064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1712622712
transform 1 0 3056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1712622712
transform 1 0 3016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1712622712
transform 1 0 3008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1712622712
transform 1 0 3000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1712622712
transform 1 0 2960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1712622712
transform 1 0 2952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1712622712
transform 1 0 2944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1712622712
transform 1 0 2920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1712622712
transform 1 0 2880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1712622712
transform 1 0 2872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1712622712
transform 1 0 2864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1712622712
transform 1 0 2856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1712622712
transform 1 0 2824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1712622712
transform 1 0 2816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1712622712
transform 1 0 2760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1712622712
transform 1 0 2736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1712622712
transform 1 0 2728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1712622712
transform 1 0 2720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1712622712
transform 1 0 2712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1712622712
transform 1 0 2704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1712622712
transform 1 0 2696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1712622712
transform 1 0 2632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1712622712
transform 1 0 2624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1712622712
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1712622712
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1712622712
transform 1 0 2536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1712622712
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1712622712
transform 1 0 2520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1712622712
transform 1 0 2512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1712622712
transform 1 0 2480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1712622712
transform 1 0 2472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1712622712
transform 1 0 2432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1712622712
transform 1 0 2424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1712622712
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1712622712
transform 1 0 2376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1712622712
transform 1 0 2368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1712622712
transform 1 0 2320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1712622712
transform 1 0 2312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1712622712
transform 1 0 2304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1712622712
transform 1 0 2296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1712622712
transform 1 0 2272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1712622712
transform 1 0 2232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1712622712
transform 1 0 2224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1712622712
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1712622712
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1712622712
transform 1 0 2160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1712622712
transform 1 0 2152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1712622712
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1712622712
transform 1 0 2112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1712622712
transform 1 0 2104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1712622712
transform 1 0 2096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1712622712
transform 1 0 2056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1712622712
transform 1 0 2016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1712622712
transform 1 0 2008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1712622712
transform 1 0 2000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1712622712
transform 1 0 1992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1712622712
transform 1 0 1984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1712622712
transform 1 0 1952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1712622712
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1712622712
transform 1 0 1896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1712622712
transform 1 0 1888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1712622712
transform 1 0 1880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1712622712
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1712622712
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1712622712
transform 1 0 1856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1712622712
transform 1 0 1784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1712622712
transform 1 0 1776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1712622712
transform 1 0 1768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1712622712
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1712622712
transform 1 0 1752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1712622712
transform 1 0 1704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1712622712
transform 1 0 1696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1712622712
transform 1 0 1672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1712622712
transform 1 0 1664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1712622712
transform 1 0 1656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1712622712
transform 1 0 1616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1712622712
transform 1 0 1576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1712622712
transform 1 0 1568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1712622712
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1712622712
transform 1 0 1552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1712622712
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1712622712
transform 1 0 1480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1712622712
transform 1 0 1472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1712622712
transform 1 0 1464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1712622712
transform 1 0 1456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1712622712
transform 1 0 1400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1712622712
transform 1 0 1392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1712622712
transform 1 0 1384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1712622712
transform 1 0 1376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1712622712
transform 1 0 1344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1712622712
transform 1 0 1296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1712622712
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1712622712
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1712622712
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1712622712
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1712622712
transform 1 0 1216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1712622712
transform 1 0 1184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1712622712
transform 1 0 1176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1712622712
transform 1 0 1168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1712622712
transform 1 0 1160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1712622712
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1712622712
transform 1 0 1120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1712622712
transform 1 0 1072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1712622712
transform 1 0 1064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1712622712
transform 1 0 1056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1712622712
transform 1 0 1048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1712622712
transform 1 0 1000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1712622712
transform 1 0 992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1712622712
transform 1 0 952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1712622712
transform 1 0 944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1712622712
transform 1 0 936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1712622712
transform 1 0 928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1712622712
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1712622712
transform 1 0 848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1712622712
transform 1 0 840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1712622712
transform 1 0 832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1712622712
transform 1 0 824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1712622712
transform 1 0 768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1712622712
transform 1 0 760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1712622712
transform 1 0 752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1712622712
transform 1 0 712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1712622712
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1712622712
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1712622712
transform 1 0 648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1712622712
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1712622712
transform 1 0 632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1712622712
transform 1 0 600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1712622712
transform 1 0 592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1712622712
transform 1 0 584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1712622712
transform 1 0 544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1712622712
transform 1 0 536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1712622712
transform 1 0 488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1712622712
transform 1 0 480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1712622712
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1712622712
transform 1 0 424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1712622712
transform 1 0 416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1712622712
transform 1 0 408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1712622712
transform 1 0 360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1712622712
transform 1 0 352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1712622712
transform 1 0 312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1712622712
transform 1 0 304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1712622712
transform 1 0 264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1712622712
transform 1 0 256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1712622712
transform 1 0 248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1712622712
transform 1 0 200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1712622712
transform 1 0 192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1712622712
transform 1 0 184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1712622712
transform 1 0 152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1712622712
transform 1 0 144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1712622712
transform 1 0 104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1712622712
transform 1 0 96 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1712622712
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1712622712
transform 1 0 3424 0 1 1770
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1712622712
transform 1 0 3416 0 1 1770
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1712622712
transform 1 0 3408 0 1 1770
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1712622712
transform 1 0 3400 0 1 1770
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1712622712
transform 1 0 3392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1712622712
transform 1 0 3384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1712622712
transform 1 0 3376 0 1 1770
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1712622712
transform 1 0 3368 0 1 1770
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1712622712
transform 1 0 3320 0 1 1770
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1712622712
transform 1 0 3312 0 1 1770
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1712622712
transform 1 0 3304 0 1 1770
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1712622712
transform 1 0 3272 0 1 1770
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1712622712
transform 1 0 3264 0 1 1770
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1712622712
transform 1 0 3256 0 1 1770
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1712622712
transform 1 0 3248 0 1 1770
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1712622712
transform 1 0 3240 0 1 1770
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1712622712
transform 1 0 3208 0 1 1770
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1712622712
transform 1 0 3168 0 1 1770
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1712622712
transform 1 0 3160 0 1 1770
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1712622712
transform 1 0 3152 0 1 1770
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1712622712
transform 1 0 3128 0 1 1770
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1712622712
transform 1 0 3120 0 1 1770
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1712622712
transform 1 0 3112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1712622712
transform 1 0 3072 0 1 1770
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1712622712
transform 1 0 3064 0 1 1770
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1712622712
transform 1 0 3056 0 1 1770
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1712622712
transform 1 0 3048 0 1 1770
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1712622712
transform 1 0 3008 0 1 1770
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1712622712
transform 1 0 3000 0 1 1770
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1712622712
transform 1 0 2992 0 1 1770
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1712622712
transform 1 0 2944 0 1 1770
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1712622712
transform 1 0 2936 0 1 1770
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1712622712
transform 1 0 2928 0 1 1770
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1712622712
transform 1 0 2920 0 1 1770
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1712622712
transform 1 0 2912 0 1 1770
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1712622712
transform 1 0 2888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1712622712
transform 1 0 2840 0 1 1770
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1712622712
transform 1 0 2832 0 1 1770
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1712622712
transform 1 0 2824 0 1 1770
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1712622712
transform 1 0 2816 0 1 1770
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1712622712
transform 1 0 2768 0 1 1770
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1712622712
transform 1 0 2760 0 1 1770
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1712622712
transform 1 0 2752 0 1 1770
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1712622712
transform 1 0 2744 0 1 1770
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1712622712
transform 1 0 2696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1712622712
transform 1 0 2688 0 1 1770
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1712622712
transform 1 0 2680 0 1 1770
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1712622712
transform 1 0 2640 0 1 1770
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1712622712
transform 1 0 2632 0 1 1770
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1712622712
transform 1 0 2624 0 1 1770
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1712622712
transform 1 0 2616 0 1 1770
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1712622712
transform 1 0 2576 0 1 1770
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1712622712
transform 1 0 2536 0 1 1770
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1712622712
transform 1 0 2528 0 1 1770
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1712622712
transform 1 0 2520 0 1 1770
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1712622712
transform 1 0 2512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1712622712
transform 1 0 2488 0 1 1770
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1712622712
transform 1 0 2448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1712622712
transform 1 0 2440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1712622712
transform 1 0 2432 0 1 1770
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1712622712
transform 1 0 2424 0 1 1770
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1712622712
transform 1 0 2368 0 1 1770
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1712622712
transform 1 0 2360 0 1 1770
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1712622712
transform 1 0 2352 0 1 1770
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1712622712
transform 1 0 2344 0 1 1770
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1712622712
transform 1 0 2312 0 1 1770
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1712622712
transform 1 0 2264 0 1 1770
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1712622712
transform 1 0 2256 0 1 1770
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1712622712
transform 1 0 2248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1712622712
transform 1 0 2240 0 1 1770
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1712622712
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1712622712
transform 1 0 2184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1712622712
transform 1 0 2176 0 1 1770
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1712622712
transform 1 0 2128 0 1 1770
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1712622712
transform 1 0 2120 0 1 1770
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1712622712
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1712622712
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1712622712
transform 1 0 2056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1712622712
transform 1 0 2048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1712622712
transform 1 0 2008 0 1 1770
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1712622712
transform 1 0 2000 0 1 1770
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1712622712
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1712622712
transform 1 0 1968 0 1 1770
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1712622712
transform 1 0 1960 0 1 1770
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1712622712
transform 1 0 1952 0 1 1770
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1712622712
transform 1 0 1888 0 1 1770
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1712622712
transform 1 0 1880 0 1 1770
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1712622712
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1712622712
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1712622712
transform 1 0 1792 0 1 1770
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1712622712
transform 1 0 1784 0 1 1770
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1712622712
transform 1 0 1776 0 1 1770
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1712622712
transform 1 0 1768 0 1 1770
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1712622712
transform 1 0 1760 0 1 1770
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1712622712
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1712622712
transform 1 0 1688 0 1 1770
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1712622712
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1712622712
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1712622712
transform 1 0 1632 0 1 1770
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1712622712
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1712622712
transform 1 0 1576 0 1 1770
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1712622712
transform 1 0 1568 0 1 1770
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1712622712
transform 1 0 1560 0 1 1770
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1712622712
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1712622712
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1712622712
transform 1 0 1456 0 1 1770
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1712622712
transform 1 0 1448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1712622712
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1712622712
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1712622712
transform 1 0 1368 0 1 1770
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1712622712
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1712622712
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1712622712
transform 1 0 1344 0 1 1770
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1712622712
transform 1 0 1280 0 1 1770
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1712622712
transform 1 0 1272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1712622712
transform 1 0 1232 0 1 1770
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1712622712
transform 1 0 1224 0 1 1770
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1712622712
transform 1 0 1216 0 1 1770
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1712622712
transform 1 0 1208 0 1 1770
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1712622712
transform 1 0 1160 0 1 1770
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1712622712
transform 1 0 1152 0 1 1770
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1712622712
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1712622712
transform 1 0 1104 0 1 1770
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1712622712
transform 1 0 1096 0 1 1770
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1712622712
transform 1 0 1088 0 1 1770
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1712622712
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1712622712
transform 1 0 1032 0 1 1770
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1712622712
transform 1 0 1024 0 1 1770
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1712622712
transform 1 0 976 0 1 1770
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1712622712
transform 1 0 968 0 1 1770
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1712622712
transform 1 0 960 0 1 1770
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1712622712
transform 1 0 952 0 1 1770
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1712622712
transform 1 0 904 0 1 1770
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1712622712
transform 1 0 896 0 1 1770
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1712622712
transform 1 0 888 0 1 1770
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1712622712
transform 1 0 848 0 1 1770
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1712622712
transform 1 0 840 0 1 1770
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1712622712
transform 1 0 832 0 1 1770
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1712622712
transform 1 0 808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1712622712
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1712622712
transform 1 0 768 0 1 1770
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1712622712
transform 1 0 760 0 1 1770
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1712622712
transform 1 0 736 0 1 1770
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1712622712
transform 1 0 728 0 1 1770
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1712622712
transform 1 0 688 0 1 1770
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1712622712
transform 1 0 680 0 1 1770
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1712622712
transform 1 0 672 0 1 1770
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1712622712
transform 1 0 664 0 1 1770
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1712622712
transform 1 0 624 0 1 1770
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1712622712
transform 1 0 616 0 1 1770
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1712622712
transform 1 0 608 0 1 1770
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1712622712
transform 1 0 600 0 1 1770
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1712622712
transform 1 0 552 0 1 1770
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1712622712
transform 1 0 544 0 1 1770
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1712622712
transform 1 0 536 0 1 1770
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1712622712
transform 1 0 528 0 1 1770
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1712622712
transform 1 0 480 0 1 1770
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1712622712
transform 1 0 472 0 1 1770
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1712622712
transform 1 0 464 0 1 1770
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1712622712
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1712622712
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1712622712
transform 1 0 400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1712622712
transform 1 0 392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1712622712
transform 1 0 384 0 1 1770
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1712622712
transform 1 0 376 0 1 1770
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1712622712
transform 1 0 320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1712622712
transform 1 0 312 0 1 1770
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1712622712
transform 1 0 304 0 1 1770
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1712622712
transform 1 0 296 0 1 1770
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1712622712
transform 1 0 288 0 1 1770
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1712622712
transform 1 0 280 0 1 1770
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1712622712
transform 1 0 272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1712622712
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1712622712
transform 1 0 200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1712622712
transform 1 0 192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1712622712
transform 1 0 184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1712622712
transform 1 0 176 0 1 1770
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1712622712
transform 1 0 168 0 1 1770
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1712622712
transform 1 0 136 0 1 1770
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1712622712
transform 1 0 88 0 1 1770
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1712622712
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1712622712
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1712622712
transform 1 0 3424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1712622712
transform 1 0 3320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1712622712
transform 1 0 3312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1712622712
transform 1 0 3240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1712622712
transform 1 0 3232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1712622712
transform 1 0 3224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1712622712
transform 1 0 3192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1712622712
transform 1 0 3152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1712622712
transform 1 0 3144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1712622712
transform 1 0 3136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1712622712
transform 1 0 3088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1712622712
transform 1 0 3080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1712622712
transform 1 0 3072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1712622712
transform 1 0 3064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1712622712
transform 1 0 3016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1712622712
transform 1 0 3008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1712622712
transform 1 0 3000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1712622712
transform 1 0 2952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1712622712
transform 1 0 2944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1712622712
transform 1 0 2936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1712622712
transform 1 0 2888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1712622712
transform 1 0 2880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1712622712
transform 1 0 2872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1712622712
transform 1 0 2864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1712622712
transform 1 0 2856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1712622712
transform 1 0 2784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1712622712
transform 1 0 2776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1712622712
transform 1 0 2768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1712622712
transform 1 0 2760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1712622712
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1712622712
transform 1 0 2712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1712622712
transform 1 0 2704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1712622712
transform 1 0 2696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1712622712
transform 1 0 2640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1712622712
transform 1 0 2632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1712622712
transform 1 0 2624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1712622712
transform 1 0 2616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1712622712
transform 1 0 2576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1712622712
transform 1 0 2552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1712622712
transform 1 0 2544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1712622712
transform 1 0 2536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1712622712
transform 1 0 2528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1712622712
transform 1 0 2480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1712622712
transform 1 0 2472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1712622712
transform 1 0 2464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1712622712
transform 1 0 2456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1712622712
transform 1 0 2408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1712622712
transform 1 0 2400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1712622712
transform 1 0 2392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1712622712
transform 1 0 2384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1712622712
transform 1 0 2336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1712622712
transform 1 0 2328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1712622712
transform 1 0 2320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1712622712
transform 1 0 2288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1712622712
transform 1 0 2280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1712622712
transform 1 0 2272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1712622712
transform 1 0 2264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1712622712
transform 1 0 2216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1712622712
transform 1 0 2208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1712622712
transform 1 0 2176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1712622712
transform 1 0 2168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1712622712
transform 1 0 2160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1712622712
transform 1 0 2152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1712622712
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1712622712
transform 1 0 2088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1712622712
transform 1 0 2080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1712622712
transform 1 0 2072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1712622712
transform 1 0 2064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1712622712
transform 1 0 2016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1712622712
transform 1 0 2008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1712622712
transform 1 0 1968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1712622712
transform 1 0 1960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1712622712
transform 1 0 1952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1712622712
transform 1 0 1920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1712622712
transform 1 0 1912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1712622712
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1712622712
transform 1 0 1856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1712622712
transform 1 0 1848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1712622712
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1712622712
transform 1 0 1808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1712622712
transform 1 0 1800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1712622712
transform 1 0 1768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1712622712
transform 1 0 1760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1712622712
transform 1 0 1720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1712622712
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1712622712
transform 1 0 1656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1712622712
transform 1 0 1648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1712622712
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1712622712
transform 1 0 1576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1712622712
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1712622712
transform 1 0 1560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1712622712
transform 1 0 1552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1712622712
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1712622712
transform 1 0 1504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1712622712
transform 1 0 1464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1712622712
transform 1 0 1456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1712622712
transform 1 0 1448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1712622712
transform 1 0 1440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1712622712
transform 1 0 1400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1712622712
transform 1 0 1392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1712622712
transform 1 0 1384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1712622712
transform 1 0 1376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1712622712
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1712622712
transform 1 0 1328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1712622712
transform 1 0 1320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1712622712
transform 1 0 1312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1712622712
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1712622712
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1712622712
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1712622712
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1712622712
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1712622712
transform 1 0 1224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1712622712
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1712622712
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1712622712
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1712622712
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1712622712
transform 1 0 1104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1712622712
transform 1 0 1096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1712622712
transform 1 0 1088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1712622712
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1712622712
transform 1 0 1040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1712622712
transform 1 0 1032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1712622712
transform 1 0 1024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1712622712
transform 1 0 984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1712622712
transform 1 0 976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1712622712
transform 1 0 968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1712622712
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1712622712
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1712622712
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1712622712
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1712622712
transform 1 0 864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1712622712
transform 1 0 856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1712622712
transform 1 0 824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1712622712
transform 1 0 816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1712622712
transform 1 0 808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1712622712
transform 1 0 776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1712622712
transform 1 0 768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1712622712
transform 1 0 760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1712622712
transform 1 0 752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1712622712
transform 1 0 704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1712622712
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1712622712
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1712622712
transform 1 0 656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1712622712
transform 1 0 648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1712622712
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1712622712
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1712622712
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1712622712
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1712622712
transform 1 0 552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1712622712
transform 1 0 544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1712622712
transform 1 0 536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1712622712
transform 1 0 528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1712622712
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1712622712
transform 1 0 472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1712622712
transform 1 0 464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1712622712
transform 1 0 456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1712622712
transform 1 0 448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1712622712
transform 1 0 440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1712622712
transform 1 0 376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1712622712
transform 1 0 368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1712622712
transform 1 0 360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1712622712
transform 1 0 352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1712622712
transform 1 0 344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1712622712
transform 1 0 336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1712622712
transform 1 0 328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1712622712
transform 1 0 280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1712622712
transform 1 0 272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1712622712
transform 1 0 264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1712622712
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1712622712
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1712622712
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1712622712
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1712622712
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1712622712
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1712622712
transform 1 0 160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1712622712
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1712622712
transform 1 0 144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1712622712
transform 1 0 136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1712622712
transform 1 0 104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1712622712
transform 1 0 96 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1712622712
transform 1 0 88 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1712622712
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1712622712
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1712622712
transform 1 0 3328 0 1 1570
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1712622712
transform 1 0 3320 0 1 1570
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1712622712
transform 1 0 3232 0 1 1570
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1712622712
transform 1 0 3224 0 1 1570
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1712622712
transform 1 0 3216 0 1 1570
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1712622712
transform 1 0 3208 0 1 1570
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1712622712
transform 1 0 3104 0 1 1570
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1712622712
transform 1 0 3096 0 1 1570
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1712622712
transform 1 0 3064 0 1 1570
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1712622712
transform 1 0 3016 0 1 1570
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1712622712
transform 1 0 3008 0 1 1570
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1712622712
transform 1 0 3000 0 1 1570
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1712622712
transform 1 0 2992 0 1 1570
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1712622712
transform 1 0 2936 0 1 1570
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1712622712
transform 1 0 2928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1712622712
transform 1 0 2920 0 1 1570
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1712622712
transform 1 0 2912 0 1 1570
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1712622712
transform 1 0 2904 0 1 1570
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1712622712
transform 1 0 2896 0 1 1570
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1712622712
transform 1 0 2832 0 1 1570
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1712622712
transform 1 0 2824 0 1 1570
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1712622712
transform 1 0 2816 0 1 1570
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1712622712
transform 1 0 2776 0 1 1570
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1712622712
transform 1 0 2768 0 1 1570
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1712622712
transform 1 0 2760 0 1 1570
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1712622712
transform 1 0 2728 0 1 1570
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1712622712
transform 1 0 2720 0 1 1570
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1712622712
transform 1 0 2712 0 1 1570
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1712622712
transform 1 0 2680 0 1 1570
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1712622712
transform 1 0 2672 0 1 1570
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1712622712
transform 1 0 2632 0 1 1570
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1712622712
transform 1 0 2624 0 1 1570
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1712622712
transform 1 0 2616 0 1 1570
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1712622712
transform 1 0 2608 0 1 1570
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1712622712
transform 1 0 2600 0 1 1570
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1712622712
transform 1 0 2536 0 1 1570
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1712622712
transform 1 0 2528 0 1 1570
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1712622712
transform 1 0 2520 0 1 1570
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1712622712
transform 1 0 2512 0 1 1570
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1712622712
transform 1 0 2504 0 1 1570
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1712622712
transform 1 0 2480 0 1 1570
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1712622712
transform 1 0 2440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1712622712
transform 1 0 2432 0 1 1570
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1712622712
transform 1 0 2424 0 1 1570
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1712622712
transform 1 0 2416 0 1 1570
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1712622712
transform 1 0 2376 0 1 1570
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1712622712
transform 1 0 2368 0 1 1570
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1712622712
transform 1 0 2328 0 1 1570
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1712622712
transform 1 0 2320 0 1 1570
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1712622712
transform 1 0 2312 0 1 1570
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1712622712
transform 1 0 2304 0 1 1570
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1712622712
transform 1 0 2264 0 1 1570
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1712622712
transform 1 0 2256 0 1 1570
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1712622712
transform 1 0 2232 0 1 1570
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1712622712
transform 1 0 2224 0 1 1570
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1712622712
transform 1 0 2216 0 1 1570
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1712622712
transform 1 0 2176 0 1 1570
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1712622712
transform 1 0 2168 0 1 1570
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1712622712
transform 1 0 2160 0 1 1570
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1712622712
transform 1 0 2136 0 1 1570
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1712622712
transform 1 0 2104 0 1 1570
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1712622712
transform 1 0 2096 0 1 1570
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1712622712
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1712622712
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1712622712
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1712622712
transform 1 0 2064 0 1 1570
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1712622712
transform 1 0 2000 0 1 1570
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1712622712
transform 1 0 1992 0 1 1570
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1712622712
transform 1 0 1984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1712622712
transform 1 0 1976 0 1 1570
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1712622712
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1712622712
transform 1 0 1904 0 1 1570
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1712622712
transform 1 0 1896 0 1 1570
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1712622712
transform 1 0 1888 0 1 1570
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1712622712
transform 1 0 1880 0 1 1570
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1712622712
transform 1 0 1872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1712622712
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1712622712
transform 1 0 1792 0 1 1570
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1712622712
transform 1 0 1784 0 1 1570
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1712622712
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1712622712
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1712622712
transform 1 0 1760 0 1 1570
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1712622712
transform 1 0 1696 0 1 1570
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1712622712
transform 1 0 1688 0 1 1570
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1712622712
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1712622712
transform 1 0 1672 0 1 1570
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1712622712
transform 1 0 1632 0 1 1570
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1712622712
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1712622712
transform 1 0 1576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1712622712
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1712622712
transform 1 0 1560 0 1 1570
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1712622712
transform 1 0 1552 0 1 1570
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1712622712
transform 1 0 1512 0 1 1570
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1712622712
transform 1 0 1504 0 1 1570
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1712622712
transform 1 0 1456 0 1 1570
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1712622712
transform 1 0 1448 0 1 1570
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1712622712
transform 1 0 1440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1712622712
transform 1 0 1432 0 1 1570
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1712622712
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1712622712
transform 1 0 1352 0 1 1570
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1712622712
transform 1 0 1344 0 1 1570
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1712622712
transform 1 0 1336 0 1 1570
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1712622712
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1712622712
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1712622712
transform 1 0 1256 0 1 1570
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1712622712
transform 1 0 1248 0 1 1570
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1712622712
transform 1 0 1240 0 1 1570
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1712622712
transform 1 0 1232 0 1 1570
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1712622712
transform 1 0 1168 0 1 1570
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1712622712
transform 1 0 1160 0 1 1570
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1712622712
transform 1 0 1152 0 1 1570
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1712622712
transform 1 0 1144 0 1 1570
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1712622712
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1712622712
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1712622712
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1712622712
transform 1 0 1072 0 1 1570
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1712622712
transform 1 0 1000 0 1 1570
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1712622712
transform 1 0 992 0 1 1570
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1712622712
transform 1 0 984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1712622712
transform 1 0 944 0 1 1570
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1712622712
transform 1 0 936 0 1 1570
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1712622712
transform 1 0 928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1712622712
transform 1 0 920 0 1 1570
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1712622712
transform 1 0 848 0 1 1570
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1712622712
transform 1 0 840 0 1 1570
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1712622712
transform 1 0 832 0 1 1570
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1712622712
transform 1 0 824 0 1 1570
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1712622712
transform 1 0 816 0 1 1570
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1712622712
transform 1 0 808 0 1 1570
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1712622712
transform 1 0 744 0 1 1570
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1712622712
transform 1 0 736 0 1 1570
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1712622712
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1712622712
transform 1 0 704 0 1 1570
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1712622712
transform 1 0 696 0 1 1570
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1712622712
transform 1 0 656 0 1 1570
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1712622712
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1712622712
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1712622712
transform 1 0 600 0 1 1570
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1712622712
transform 1 0 592 0 1 1570
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1712622712
transform 1 0 544 0 1 1570
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1712622712
transform 1 0 536 0 1 1570
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1712622712
transform 1 0 528 0 1 1570
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1712622712
transform 1 0 472 0 1 1570
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1712622712
transform 1 0 464 0 1 1570
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1712622712
transform 1 0 456 0 1 1570
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1712622712
transform 1 0 408 0 1 1570
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1712622712
transform 1 0 400 0 1 1570
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1712622712
transform 1 0 392 0 1 1570
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1712622712
transform 1 0 352 0 1 1570
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1712622712
transform 1 0 320 0 1 1570
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1712622712
transform 1 0 312 0 1 1570
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1712622712
transform 1 0 304 0 1 1570
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1712622712
transform 1 0 256 0 1 1570
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1712622712
transform 1 0 248 0 1 1570
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1712622712
transform 1 0 240 0 1 1570
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1712622712
transform 1 0 192 0 1 1570
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1712622712
transform 1 0 184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1712622712
transform 1 0 176 0 1 1570
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1712622712
transform 1 0 168 0 1 1570
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1712622712
transform 1 0 120 0 1 1570
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1712622712
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1712622712
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1712622712
transform 1 0 3424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1712622712
transform 1 0 3416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1712622712
transform 1 0 3360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1712622712
transform 1 0 3352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1712622712
transform 1 0 3344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1712622712
transform 1 0 3336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1712622712
transform 1 0 3328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1712622712
transform 1 0 3272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1712622712
transform 1 0 3264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1712622712
transform 1 0 3256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1712622712
transform 1 0 3248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1712622712
transform 1 0 3144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1712622712
transform 1 0 3136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1712622712
transform 1 0 3128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1712622712
transform 1 0 3120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1712622712
transform 1 0 3056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1712622712
transform 1 0 3048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1712622712
transform 1 0 3040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1712622712
transform 1 0 3032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1712622712
transform 1 0 2992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1712622712
transform 1 0 2984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1712622712
transform 1 0 2944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1712622712
transform 1 0 2936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1712622712
transform 1 0 2928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1712622712
transform 1 0 2888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1712622712
transform 1 0 2880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1712622712
transform 1 0 2872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1712622712
transform 1 0 2840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1712622712
transform 1 0 2832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1712622712
transform 1 0 2792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1712622712
transform 1 0 2784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1712622712
transform 1 0 2776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1712622712
transform 1 0 2744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1712622712
transform 1 0 2736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1712622712
transform 1 0 2696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1712622712
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1712622712
transform 1 0 2680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1712622712
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1712622712
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1712622712
transform 1 0 2624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1712622712
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1712622712
transform 1 0 2584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1712622712
transform 1 0 2552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1712622712
transform 1 0 2544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1712622712
transform 1 0 2536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1712622712
transform 1 0 2480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1712622712
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1712622712
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1712622712
transform 1 0 2456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1712622712
transform 1 0 2448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1712622712
transform 1 0 2392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1712622712
transform 1 0 2384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1712622712
transform 1 0 2376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1712622712
transform 1 0 2368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1712622712
transform 1 0 2304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1712622712
transform 1 0 2296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1712622712
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1712622712
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1712622712
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1712622712
transform 1 0 2224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1712622712
transform 1 0 2216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1712622712
transform 1 0 2176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1712622712
transform 1 0 2168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1712622712
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1712622712
transform 1 0 2152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1712622712
transform 1 0 2104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1712622712
transform 1 0 2096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1712622712
transform 1 0 2088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1712622712
transform 1 0 2056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1712622712
transform 1 0 2048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1712622712
transform 1 0 2008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1712622712
transform 1 0 2000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1712622712
transform 1 0 1992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1712622712
transform 1 0 1944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1712622712
transform 1 0 1936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1712622712
transform 1 0 1928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1712622712
transform 1 0 1888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1712622712
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1712622712
transform 1 0 1872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1712622712
transform 1 0 1840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1712622712
transform 1 0 1808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1712622712
transform 1 0 1800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1712622712
transform 1 0 1792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1712622712
transform 1 0 1784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1712622712
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1712622712
transform 1 0 1736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1712622712
transform 1 0 1696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1712622712
transform 1 0 1688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1712622712
transform 1 0 1680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1712622712
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1712622712
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1712622712
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1712622712
transform 1 0 1584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1712622712
transform 1 0 1576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1712622712
transform 1 0 1568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1712622712
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1712622712
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1712622712
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1712622712
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1712622712
transform 1 0 1472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1712622712
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1712622712
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1712622712
transform 1 0 1384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1712622712
transform 1 0 1376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1712622712
transform 1 0 1368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1712622712
transform 1 0 1360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1712622712
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1712622712
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1712622712
transform 1 0 1288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1712622712
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1712622712
transform 1 0 1272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1712622712
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1712622712
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1712622712
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1712622712
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1712622712
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1712622712
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1712622712
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1712622712
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1712622712
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1712622712
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1712622712
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1712622712
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1712622712
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1712622712
transform 1 0 960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1712622712
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1712622712
transform 1 0 944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1712622712
transform 1 0 936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1712622712
transform 1 0 928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1712622712
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1712622712
transform 1 0 856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1712622712
transform 1 0 848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1712622712
transform 1 0 840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1712622712
transform 1 0 808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1712622712
transform 1 0 800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1712622712
transform 1 0 792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1712622712
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1712622712
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1712622712
transform 1 0 736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1712622712
transform 1 0 696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1712622712
transform 1 0 688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1712622712
transform 1 0 680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1712622712
transform 1 0 672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1712622712
transform 1 0 632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1712622712
transform 1 0 624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1712622712
transform 1 0 584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1712622712
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1712622712
transform 1 0 568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1712622712
transform 1 0 560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1712622712
transform 1 0 512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1712622712
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1712622712
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1712622712
transform 1 0 456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1712622712
transform 1 0 448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1712622712
transform 1 0 400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1712622712
transform 1 0 392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1712622712
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1712622712
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1712622712
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1712622712
transform 1 0 336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1712622712
transform 1 0 328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1712622712
transform 1 0 288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1712622712
transform 1 0 280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1712622712
transform 1 0 272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1712622712
transform 1 0 264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1712622712
transform 1 0 256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1712622712
transform 1 0 200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1712622712
transform 1 0 192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1712622712
transform 1 0 184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1712622712
transform 1 0 176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1712622712
transform 1 0 168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1712622712
transform 1 0 160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1712622712
transform 1 0 128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1712622712
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1712622712
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1712622712
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1712622712
transform 1 0 3424 0 1 1370
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1712622712
transform 1 0 3416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1712622712
transform 1 0 3408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1712622712
transform 1 0 3360 0 1 1370
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1712622712
transform 1 0 3352 0 1 1370
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1712622712
transform 1 0 3312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1712622712
transform 1 0 3304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1712622712
transform 1 0 3296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1712622712
transform 1 0 3288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1712622712
transform 1 0 3280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1712622712
transform 1 0 3224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1712622712
transform 1 0 3216 0 1 1370
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1712622712
transform 1 0 3208 0 1 1370
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1712622712
transform 1 0 3200 0 1 1370
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1712622712
transform 1 0 3192 0 1 1370
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1712622712
transform 1 0 3184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1712622712
transform 1 0 3152 0 1 1370
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1712622712
transform 1 0 3144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1712622712
transform 1 0 3136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1712622712
transform 1 0 3128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1712622712
transform 1 0 3120 0 1 1370
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1712622712
transform 1 0 3112 0 1 1370
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1712622712
transform 1 0 3104 0 1 1370
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1712622712
transform 1 0 3072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1712622712
transform 1 0 3064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1712622712
transform 1 0 3056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1712622712
transform 1 0 3016 0 1 1370
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1712622712
transform 1 0 3008 0 1 1370
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1712622712
transform 1 0 3000 0 1 1370
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1712622712
transform 1 0 2992 0 1 1370
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1712622712
transform 1 0 2984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1712622712
transform 1 0 2976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1712622712
transform 1 0 2936 0 1 1370
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1712622712
transform 1 0 2928 0 1 1370
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1712622712
transform 1 0 2920 0 1 1370
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1712622712
transform 1 0 2912 0 1 1370
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1712622712
transform 1 0 2872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1712622712
transform 1 0 2864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1712622712
transform 1 0 2840 0 1 1370
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1712622712
transform 1 0 2832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1712622712
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1712622712
transform 1 0 2792 0 1 1370
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1712622712
transform 1 0 2784 0 1 1370
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1712622712
transform 1 0 2760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1712622712
transform 1 0 2752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1712622712
transform 1 0 2744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1712622712
transform 1 0 2736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1712622712
transform 1 0 2688 0 1 1370
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1712622712
transform 1 0 2680 0 1 1370
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1712622712
transform 1 0 2672 0 1 1370
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1712622712
transform 1 0 2664 0 1 1370
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1712622712
transform 1 0 2656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1712622712
transform 1 0 2616 0 1 1370
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1712622712
transform 1 0 2608 0 1 1370
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1712622712
transform 1 0 2600 0 1 1370
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1712622712
transform 1 0 2560 0 1 1370
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1712622712
transform 1 0 2552 0 1 1370
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1712622712
transform 1 0 2544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1712622712
transform 1 0 2536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1712622712
transform 1 0 2528 0 1 1370
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1712622712
transform 1 0 2480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1712622712
transform 1 0 2472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1712622712
transform 1 0 2464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1712622712
transform 1 0 2456 0 1 1370
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1712622712
transform 1 0 2416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1712622712
transform 1 0 2408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1712622712
transform 1 0 2400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1712622712
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1712622712
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1712622712
transform 1 0 2328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1712622712
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1712622712
transform 1 0 2296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1712622712
transform 1 0 2288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1712622712
transform 1 0 2280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1712622712
transform 1 0 2240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1712622712
transform 1 0 2232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1712622712
transform 1 0 2224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1712622712
transform 1 0 2184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1712622712
transform 1 0 2176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1712622712
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1712622712
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1712622712
transform 1 0 2120 0 1 1370
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1712622712
transform 1 0 2112 0 1 1370
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1712622712
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1712622712
transform 1 0 2064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1712622712
transform 1 0 2056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1712622712
transform 1 0 2016 0 1 1370
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1712622712
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1712622712
transform 1 0 2000 0 1 1370
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1712622712
transform 1 0 1952 0 1 1370
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1712622712
transform 1 0 1944 0 1 1370
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1712622712
transform 1 0 1936 0 1 1370
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1712622712
transform 1 0 1896 0 1 1370
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1712622712
transform 1 0 1888 0 1 1370
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1712622712
transform 1 0 1880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1712622712
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1712622712
transform 1 0 1864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1712622712
transform 1 0 1808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1712622712
transform 1 0 1800 0 1 1370
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1712622712
transform 1 0 1792 0 1 1370
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1712622712
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1712622712
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1712622712
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1712622712
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1712622712
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1712622712
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1712622712
transform 1 0 1656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1712622712
transform 1 0 1648 0 1 1370
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1712622712
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1712622712
transform 1 0 1632 0 1 1370
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1712622712
transform 1 0 1592 0 1 1370
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1712622712
transform 1 0 1584 0 1 1370
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1712622712
transform 1 0 1576 0 1 1370
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1712622712
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1712622712
transform 1 0 1520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1712622712
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1712622712
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1712622712
transform 1 0 1496 0 1 1370
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1712622712
transform 1 0 1488 0 1 1370
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1712622712
transform 1 0 1480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1712622712
transform 1 0 1416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1712622712
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1712622712
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1712622712
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1712622712
transform 1 0 1384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1712622712
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1712622712
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1712622712
transform 1 0 1304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1712622712
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1712622712
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1712622712
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1712622712
transform 1 0 1224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1712622712
transform 1 0 1216 0 1 1370
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1712622712
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1712622712
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1712622712
transform 1 0 1168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1712622712
transform 1 0 1136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1712622712
transform 1 0 1128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1712622712
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1712622712
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1712622712
transform 1 0 1072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1712622712
transform 1 0 1064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1712622712
transform 1 0 1016 0 1 1370
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1712622712
transform 1 0 1008 0 1 1370
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1712622712
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1712622712
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1712622712
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1712622712
transform 1 0 944 0 1 1370
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1712622712
transform 1 0 920 0 1 1370
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1712622712
transform 1 0 880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1712622712
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1712622712
transform 1 0 864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1712622712
transform 1 0 856 0 1 1370
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1712622712
transform 1 0 848 0 1 1370
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1712622712
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1712622712
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1712622712
transform 1 0 768 0 1 1370
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1712622712
transform 1 0 760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1712622712
transform 1 0 752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1712622712
transform 1 0 712 0 1 1370
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1712622712
transform 1 0 672 0 1 1370
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1712622712
transform 1 0 664 0 1 1370
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1712622712
transform 1 0 656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1712622712
transform 1 0 648 0 1 1370
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1712622712
transform 1 0 640 0 1 1370
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1712622712
transform 1 0 600 0 1 1370
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1712622712
transform 1 0 592 0 1 1370
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1712622712
transform 1 0 544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1712622712
transform 1 0 536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1712622712
transform 1 0 528 0 1 1370
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1712622712
transform 1 0 520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1712622712
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1712622712
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1712622712
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1712622712
transform 1 0 456 0 1 1370
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1712622712
transform 1 0 408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1712622712
transform 1 0 400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1712622712
transform 1 0 392 0 1 1370
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1712622712
transform 1 0 384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1712622712
transform 1 0 352 0 1 1370
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1712622712
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1712622712
transform 1 0 304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1712622712
transform 1 0 296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1712622712
transform 1 0 288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1712622712
transform 1 0 280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1712622712
transform 1 0 232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1712622712
transform 1 0 200 0 1 1370
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1712622712
transform 1 0 192 0 1 1370
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1712622712
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1712622712
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1712622712
transform 1 0 168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1712622712
transform 1 0 136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1712622712
transform 1 0 88 0 1 1370
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1712622712
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1712622712
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1712622712
transform 1 0 3424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1712622712
transform 1 0 3416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1712622712
transform 1 0 3376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1712622712
transform 1 0 3368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1712622712
transform 1 0 3328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1712622712
transform 1 0 3320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1712622712
transform 1 0 3312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1712622712
transform 1 0 3280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1712622712
transform 1 0 3272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1712622712
transform 1 0 3208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1712622712
transform 1 0 3200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1712622712
transform 1 0 3192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1712622712
transform 1 0 3088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1712622712
transform 1 0 3080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1712622712
transform 1 0 3072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1712622712
transform 1 0 3064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1712622712
transform 1 0 3008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1712622712
transform 1 0 3000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1712622712
transform 1 0 2992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1712622712
transform 1 0 2952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1712622712
transform 1 0 2944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1712622712
transform 1 0 2936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1712622712
transform 1 0 2928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1712622712
transform 1 0 2880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1712622712
transform 1 0 2872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1712622712
transform 1 0 2864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1712622712
transform 1 0 2856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1712622712
transform 1 0 2848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1712622712
transform 1 0 2800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1712622712
transform 1 0 2792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1712622712
transform 1 0 2784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1712622712
transform 1 0 2752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1712622712
transform 1 0 2744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1712622712
transform 1 0 2736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1712622712
transform 1 0 2704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1712622712
transform 1 0 2696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1712622712
transform 1 0 2688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1712622712
transform 1 0 2680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1712622712
transform 1 0 2624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1712622712
transform 1 0 2616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1712622712
transform 1 0 2608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1712622712
transform 1 0 2600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1712622712
transform 1 0 2576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1712622712
transform 1 0 2568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1712622712
transform 1 0 2520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1712622712
transform 1 0 2512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1712622712
transform 1 0 2504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1712622712
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1712622712
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1712622712
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1712622712
transform 1 0 2448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1712622712
transform 1 0 2440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1712622712
transform 1 0 2432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1712622712
transform 1 0 2384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1712622712
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1712622712
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1712622712
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1712622712
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1712622712
transform 1 0 2312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1712622712
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1712622712
transform 1 0 2296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1712622712
transform 1 0 2288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1712622712
transform 1 0 2248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1712622712
transform 1 0 2240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1712622712
transform 1 0 2232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1712622712
transform 1 0 2224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1712622712
transform 1 0 2184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1712622712
transform 1 0 2176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1712622712
transform 1 0 2168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1712622712
transform 1 0 2160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1712622712
transform 1 0 2152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1712622712
transform 1 0 2104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1712622712
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1712622712
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1712622712
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1712622712
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1712622712
transform 1 0 2064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1712622712
transform 1 0 2056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1712622712
transform 1 0 2008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1712622712
transform 1 0 2000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1712622712
transform 1 0 1992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1712622712
transform 1 0 1984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1712622712
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1712622712
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1712622712
transform 1 0 1936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1712622712
transform 1 0 1928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1712622712
transform 1 0 1920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1712622712
transform 1 0 1912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1712622712
transform 1 0 1904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1712622712
transform 1 0 1856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1712622712
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1712622712
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1712622712
transform 1 0 1832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1712622712
transform 1 0 1824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1712622712
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1712622712
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1712622712
transform 1 0 1768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1712622712
transform 1 0 1760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1712622712
transform 1 0 1752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1712622712
transform 1 0 1712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1712622712
transform 1 0 1704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1712622712
transform 1 0 1696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1712622712
transform 1 0 1688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1712622712
transform 1 0 1680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1712622712
transform 1 0 1640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1712622712
transform 1 0 1632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1712622712
transform 1 0 1624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1712622712
transform 1 0 1616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1712622712
transform 1 0 1608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1712622712
transform 1 0 1600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1712622712
transform 1 0 1552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1712622712
transform 1 0 1544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1712622712
transform 1 0 1536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1712622712
transform 1 0 1528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1712622712
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1712622712
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1712622712
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1712622712
transform 1 0 1456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1712622712
transform 1 0 1448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1712622712
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1712622712
transform 1 0 1432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1712622712
transform 1 0 1424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1712622712
transform 1 0 1392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1712622712
transform 1 0 1384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1712622712
transform 1 0 1376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1712622712
transform 1 0 1336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1712622712
transform 1 0 1328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1712622712
transform 1 0 1320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1712622712
transform 1 0 1312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1712622712
transform 1 0 1304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1712622712
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1712622712
transform 1 0 1248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1712622712
transform 1 0 1240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1712622712
transform 1 0 1232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1712622712
transform 1 0 1224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1712622712
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1712622712
transform 1 0 1168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1712622712
transform 1 0 1160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1712622712
transform 1 0 1152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1712622712
transform 1 0 1144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1712622712
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1712622712
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1712622712
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1712622712
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1712622712
transform 1 0 1064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1712622712
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1712622712
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1712622712
transform 1 0 1000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1712622712
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1712622712
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1712622712
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1712622712
transform 1 0 968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1712622712
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1712622712
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1712622712
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1712622712
transform 1 0 880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1712622712
transform 1 0 872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1712622712
transform 1 0 864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1712622712
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1712622712
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1712622712
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1712622712
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1712622712
transform 1 0 768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1712622712
transform 1 0 760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1712622712
transform 1 0 752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1712622712
transform 1 0 744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1712622712
transform 1 0 688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1712622712
transform 1 0 680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1712622712
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1712622712
transform 1 0 664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1712622712
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1712622712
transform 1 0 616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1712622712
transform 1 0 608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1712622712
transform 1 0 600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1712622712
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1712622712
transform 1 0 544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1712622712
transform 1 0 536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1712622712
transform 1 0 528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1712622712
transform 1 0 520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1712622712
transform 1 0 512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1712622712
transform 1 0 464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1712622712
transform 1 0 456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1712622712
transform 1 0 448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1712622712
transform 1 0 440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1712622712
transform 1 0 432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1712622712
transform 1 0 424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1712622712
transform 1 0 384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1712622712
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1712622712
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1712622712
transform 1 0 344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1712622712
transform 1 0 336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1712622712
transform 1 0 328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1712622712
transform 1 0 320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1712622712
transform 1 0 280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1712622712
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1712622712
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1712622712
transform 1 0 256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1712622712
transform 1 0 216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1712622712
transform 1 0 208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1712622712
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1712622712
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1712622712
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1712622712
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1712622712
transform 1 0 128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1712622712
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1712622712
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1712622712
transform 1 0 104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1712622712
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1712622712
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1712622712
transform 1 0 3424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1712622712
transform 1 0 3416 0 1 1170
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1712622712
transform 1 0 3408 0 1 1170
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1712622712
transform 1 0 3400 0 1 1170
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1712622712
transform 1 0 3360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1712622712
transform 1 0 3352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1712622712
transform 1 0 3344 0 1 1170
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1712622712
transform 1 0 3336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1712622712
transform 1 0 3304 0 1 1170
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1712622712
transform 1 0 3296 0 1 1170
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1712622712
transform 1 0 3288 0 1 1170
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1712622712
transform 1 0 3248 0 1 1170
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1712622712
transform 1 0 3240 0 1 1170
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1712622712
transform 1 0 3232 0 1 1170
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1712622712
transform 1 0 3224 0 1 1170
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1712622712
transform 1 0 3216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1712622712
transform 1 0 3208 0 1 1170
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1712622712
transform 1 0 3152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1712622712
transform 1 0 3144 0 1 1170
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1712622712
transform 1 0 3136 0 1 1170
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1712622712
transform 1 0 3128 0 1 1170
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1712622712
transform 1 0 3120 0 1 1170
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1712622712
transform 1 0 3112 0 1 1170
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1712622712
transform 1 0 3072 0 1 1170
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1712622712
transform 1 0 3064 0 1 1170
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1712622712
transform 1 0 3024 0 1 1170
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1712622712
transform 1 0 3016 0 1 1170
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1712622712
transform 1 0 3008 0 1 1170
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1712622712
transform 1 0 3000 0 1 1170
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1712622712
transform 1 0 2992 0 1 1170
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1712622712
transform 1 0 2944 0 1 1170
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1712622712
transform 1 0 2936 0 1 1170
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1712622712
transform 1 0 2904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1712622712
transform 1 0 2896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1712622712
transform 1 0 2888 0 1 1170
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1712622712
transform 1 0 2880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1712622712
transform 1 0 2872 0 1 1170
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1712622712
transform 1 0 2816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1712622712
transform 1 0 2808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1712622712
transform 1 0 2800 0 1 1170
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1712622712
transform 1 0 2792 0 1 1170
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1712622712
transform 1 0 2784 0 1 1170
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1712622712
transform 1 0 2728 0 1 1170
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1712622712
transform 1 0 2720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1712622712
transform 1 0 2712 0 1 1170
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1712622712
transform 1 0 2704 0 1 1170
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1712622712
transform 1 0 2696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1712622712
transform 1 0 2688 0 1 1170
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1712622712
transform 1 0 2656 0 1 1170
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1712622712
transform 1 0 2632 0 1 1170
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1712622712
transform 1 0 2608 0 1 1170
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1712622712
transform 1 0 2600 0 1 1170
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1712622712
transform 1 0 2576 0 1 1170
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1712622712
transform 1 0 2568 0 1 1170
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1712622712
transform 1 0 2560 0 1 1170
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1712622712
transform 1 0 2552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1712622712
transform 1 0 2544 0 1 1170
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1712622712
transform 1 0 2488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1712622712
transform 1 0 2480 0 1 1170
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1712622712
transform 1 0 2472 0 1 1170
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1712622712
transform 1 0 2464 0 1 1170
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1712622712
transform 1 0 2456 0 1 1170
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1712622712
transform 1 0 2424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1712622712
transform 1 0 2392 0 1 1170
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1712622712
transform 1 0 2384 0 1 1170
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1712622712
transform 1 0 2376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1712622712
transform 1 0 2368 0 1 1170
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1712622712
transform 1 0 2360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1712622712
transform 1 0 2336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1712622712
transform 1 0 2296 0 1 1170
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1712622712
transform 1 0 2288 0 1 1170
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1712622712
transform 1 0 2280 0 1 1170
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1712622712
transform 1 0 2272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1712622712
transform 1 0 2264 0 1 1170
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1712622712
transform 1 0 2216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1712622712
transform 1 0 2208 0 1 1170
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1712622712
transform 1 0 2200 0 1 1170
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1712622712
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3130
timestamp 1712622712
transform 1 0 2160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1712622712
transform 1 0 2152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1712622712
transform 1 0 2144 0 1 1170
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1712622712
transform 1 0 2136 0 1 1170
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1712622712
transform 1 0 2088 0 1 1170
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1712622712
transform 1 0 2080 0 1 1170
box -8 -3 16 105
use FILL  FILL_3136
timestamp 1712622712
transform 1 0 2072 0 1 1170
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1712622712
transform 1 0 2064 0 1 1170
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1712622712
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1712622712
transform 1 0 2024 0 1 1170
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1712622712
transform 1 0 2016 0 1 1170
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1712622712
transform 1 0 1976 0 1 1170
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1712622712
transform 1 0 1968 0 1 1170
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1712622712
transform 1 0 1960 0 1 1170
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1712622712
transform 1 0 1952 0 1 1170
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1712622712
transform 1 0 1912 0 1 1170
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1712622712
transform 1 0 1904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1712622712
transform 1 0 1896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1712622712
transform 1 0 1856 0 1 1170
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1712622712
transform 1 0 1848 0 1 1170
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1712622712
transform 1 0 1840 0 1 1170
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1712622712
transform 1 0 1832 0 1 1170
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1712622712
transform 1 0 1792 0 1 1170
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1712622712
transform 1 0 1784 0 1 1170
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1712622712
transform 1 0 1776 0 1 1170
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1712622712
transform 1 0 1768 0 1 1170
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1712622712
transform 1 0 1760 0 1 1170
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1712622712
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1712622712
transform 1 0 1712 0 1 1170
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1712622712
transform 1 0 1704 0 1 1170
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1712622712
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1712622712
transform 1 0 1656 0 1 1170
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1712622712
transform 1 0 1648 0 1 1170
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1712622712
transform 1 0 1640 0 1 1170
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1712622712
transform 1 0 1632 0 1 1170
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1712622712
transform 1 0 1584 0 1 1170
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1712622712
transform 1 0 1576 0 1 1170
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1712622712
transform 1 0 1568 0 1 1170
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1712622712
transform 1 0 1560 0 1 1170
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1712622712
transform 1 0 1552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1712622712
transform 1 0 1544 0 1 1170
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1712622712
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1712622712
transform 1 0 1488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1712622712
transform 1 0 1480 0 1 1170
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1712622712
transform 1 0 1472 0 1 1170
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1712622712
transform 1 0 1464 0 1 1170
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1712622712
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1712622712
transform 1 0 1416 0 1 1170
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1712622712
transform 1 0 1408 0 1 1170
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1712622712
transform 1 0 1400 0 1 1170
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1712622712
transform 1 0 1360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1712622712
transform 1 0 1352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1712622712
transform 1 0 1344 0 1 1170
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1712622712
transform 1 0 1336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1712622712
transform 1 0 1328 0 1 1170
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1712622712
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1712622712
transform 1 0 1288 0 1 1170
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1712622712
transform 1 0 1280 0 1 1170
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1712622712
transform 1 0 1272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1712622712
transform 1 0 1224 0 1 1170
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1712622712
transform 1 0 1216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1712622712
transform 1 0 1208 0 1 1170
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1712622712
transform 1 0 1200 0 1 1170
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1712622712
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1712622712
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1712622712
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1712622712
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1712622712
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1712622712
transform 1 0 1104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1712622712
transform 1 0 1096 0 1 1170
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1712622712
transform 1 0 1088 0 1 1170
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1712622712
transform 1 0 1080 0 1 1170
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1712622712
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1712622712
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1712622712
transform 1 0 1000 0 1 1170
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1712622712
transform 1 0 992 0 1 1170
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1712622712
transform 1 0 984 0 1 1170
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1712622712
transform 1 0 976 0 1 1170
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1712622712
transform 1 0 968 0 1 1170
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1712622712
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1712622712
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1712622712
transform 1 0 904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1712622712
transform 1 0 896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1712622712
transform 1 0 888 0 1 1170
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1712622712
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1712622712
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1712622712
transform 1 0 832 0 1 1170
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1712622712
transform 1 0 824 0 1 1170
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1712622712
transform 1 0 816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1712622712
transform 1 0 776 0 1 1170
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1712622712
transform 1 0 768 0 1 1170
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1712622712
transform 1 0 760 0 1 1170
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1712622712
transform 1 0 752 0 1 1170
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1712622712
transform 1 0 744 0 1 1170
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1712622712
transform 1 0 696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1712622712
transform 1 0 688 0 1 1170
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1712622712
transform 1 0 680 0 1 1170
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1712622712
transform 1 0 672 0 1 1170
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1712622712
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1712622712
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1712622712
transform 1 0 616 0 1 1170
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1712622712
transform 1 0 608 0 1 1170
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1712622712
transform 1 0 600 0 1 1170
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1712622712
transform 1 0 592 0 1 1170
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1712622712
transform 1 0 584 0 1 1170
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1712622712
transform 1 0 536 0 1 1170
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1712622712
transform 1 0 528 0 1 1170
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1712622712
transform 1 0 520 0 1 1170
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1712622712
transform 1 0 512 0 1 1170
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1712622712
transform 1 0 504 0 1 1170
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1712622712
transform 1 0 496 0 1 1170
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1712622712
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1712622712
transform 1 0 440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1712622712
transform 1 0 432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1712622712
transform 1 0 424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1712622712
transform 1 0 416 0 1 1170
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1712622712
transform 1 0 408 0 1 1170
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1712622712
transform 1 0 360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1712622712
transform 1 0 352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1712622712
transform 1 0 344 0 1 1170
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1712622712
transform 1 0 336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1712622712
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1712622712
transform 1 0 320 0 1 1170
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1712622712
transform 1 0 280 0 1 1170
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1712622712
transform 1 0 272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1712622712
transform 1 0 264 0 1 1170
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1712622712
transform 1 0 256 0 1 1170
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1712622712
transform 1 0 216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1712622712
transform 1 0 208 0 1 1170
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1712622712
transform 1 0 200 0 1 1170
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1712622712
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1712622712
transform 1 0 184 0 1 1170
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1712622712
transform 1 0 176 0 1 1170
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1712622712
transform 1 0 136 0 1 1170
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1712622712
transform 1 0 128 0 1 1170
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1712622712
transform 1 0 120 0 1 1170
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1712622712
transform 1 0 88 0 1 1170
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1712622712
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1712622712
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1712622712
transform 1 0 3424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1712622712
transform 1 0 3416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1712622712
transform 1 0 3408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1712622712
transform 1 0 3336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1712622712
transform 1 0 3328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1712622712
transform 1 0 3320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1712622712
transform 1 0 3312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1712622712
transform 1 0 3304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1712622712
transform 1 0 3240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1712622712
transform 1 0 3232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1712622712
transform 1 0 3224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1712622712
transform 1 0 3216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1712622712
transform 1 0 3208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1712622712
transform 1 0 3160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1712622712
transform 1 0 3120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1712622712
transform 1 0 3112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1712622712
transform 1 0 3104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1712622712
transform 1 0 3096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1712622712
transform 1 0 3056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1712622712
transform 1 0 3048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1712622712
transform 1 0 3024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1712622712
transform 1 0 3016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1712622712
transform 1 0 3008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1712622712
transform 1 0 3000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1712622712
transform 1 0 2960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1712622712
transform 1 0 2952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1712622712
transform 1 0 2920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1712622712
transform 1 0 2912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1712622712
transform 1 0 2904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1712622712
transform 1 0 2896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1712622712
transform 1 0 2856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1712622712
transform 1 0 2848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1712622712
transform 1 0 2840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1712622712
transform 1 0 2816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1712622712
transform 1 0 2808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1712622712
transform 1 0 2800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1712622712
transform 1 0 2792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1712622712
transform 1 0 2760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1712622712
transform 1 0 2728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1712622712
transform 1 0 2720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1712622712
transform 1 0 2712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1712622712
transform 1 0 2704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1712622712
transform 1 0 2696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1712622712
transform 1 0 2688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1712622712
transform 1 0 2624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1712622712
transform 1 0 2616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1712622712
transform 1 0 2608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1712622712
transform 1 0 2600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1712622712
transform 1 0 2592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1712622712
transform 1 0 2584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1712622712
transform 1 0 2528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1712622712
transform 1 0 2520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1712622712
transform 1 0 2512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1712622712
transform 1 0 2504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1712622712
transform 1 0 2496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1712622712
transform 1 0 2488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1712622712
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1712622712
transform 1 0 2432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1712622712
transform 1 0 2424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1712622712
transform 1 0 2416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3329
timestamp 1712622712
transform 1 0 2408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1712622712
transform 1 0 2368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1712622712
transform 1 0 2360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1712622712
transform 1 0 2352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1712622712
transform 1 0 2344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1712622712
transform 1 0 2336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1712622712
transform 1 0 2328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1712622712
transform 1 0 2272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1712622712
transform 1 0 2264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1712622712
transform 1 0 2256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1712622712
transform 1 0 2248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1712622712
transform 1 0 2240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1712622712
transform 1 0 2232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1712622712
transform 1 0 2224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1712622712
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1712622712
transform 1 0 2160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1712622712
transform 1 0 2152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1712622712
transform 1 0 2144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1712622712
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1712622712
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1712622712
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1712622712
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1712622712
transform 1 0 2056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1712622712
transform 1 0 2048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1712622712
transform 1 0 2040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1712622712
transform 1 0 2032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1712622712
transform 1 0 2024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1712622712
transform 1 0 2016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1712622712
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1712622712
transform 1 0 1976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1712622712
transform 1 0 1944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1712622712
transform 1 0 1936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1712622712
transform 1 0 1928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1712622712
transform 1 0 1920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1712622712
transform 1 0 1912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1712622712
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1712622712
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1712622712
transform 1 0 1840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1712622712
transform 1 0 1832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1712622712
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1712622712
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1712622712
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1712622712
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1712622712
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1712622712
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1712622712
transform 1 0 1736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1712622712
transform 1 0 1728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1712622712
transform 1 0 1720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1712622712
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1712622712
transform 1 0 1688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1712622712
transform 1 0 1664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3380
timestamp 1712622712
transform 1 0 1656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1712622712
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1712622712
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1712622712
transform 1 0 1600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1712622712
transform 1 0 1592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1712622712
transform 1 0 1584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1712622712
transform 1 0 1576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1712622712
transform 1 0 1568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1712622712
transform 1 0 1528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1712622712
transform 1 0 1520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1712622712
transform 1 0 1512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1712622712
transform 1 0 1504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1712622712
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1712622712
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1712622712
transform 1 0 1432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1712622712
transform 1 0 1424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1712622712
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1712622712
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1712622712
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3399
timestamp 1712622712
transform 1 0 1360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1712622712
transform 1 0 1352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1712622712
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1712622712
transform 1 0 1304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1712622712
transform 1 0 1296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1712622712
transform 1 0 1288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1712622712
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1712622712
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1712622712
transform 1 0 1248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1712622712
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1712622712
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1712622712
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1712622712
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1712622712
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1712622712
transform 1 0 1152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1712622712
transform 1 0 1144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1712622712
transform 1 0 1112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1712622712
transform 1 0 1104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1712622712
transform 1 0 1096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1712622712
transform 1 0 1088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1712622712
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1712622712
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1712622712
transform 1 0 1024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1712622712
transform 1 0 1016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1712622712
transform 1 0 1008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1712622712
transform 1 0 1000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1712622712
transform 1 0 968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1712622712
transform 1 0 960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1712622712
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1712622712
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1712622712
transform 1 0 912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1712622712
transform 1 0 904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1712622712
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1712622712
transform 1 0 864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1712622712
transform 1 0 856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1712622712
transform 1 0 848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1712622712
transform 1 0 808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1712622712
transform 1 0 800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1712622712
transform 1 0 792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1712622712
transform 1 0 784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1712622712
transform 1 0 760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1712622712
transform 1 0 752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1712622712
transform 1 0 712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1712622712
transform 1 0 704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1712622712
transform 1 0 696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1712622712
transform 1 0 688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1712622712
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1712622712
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1712622712
transform 1 0 616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3448
timestamp 1712622712
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1712622712
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1712622712
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1712622712
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1712622712
transform 1 0 560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1712622712
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1712622712
transform 1 0 512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1712622712
transform 1 0 504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1712622712
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1712622712
transform 1 0 488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3458
timestamp 1712622712
transform 1 0 440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1712622712
transform 1 0 432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1712622712
transform 1 0 424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1712622712
transform 1 0 416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1712622712
transform 1 0 368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1712622712
transform 1 0 360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3464
timestamp 1712622712
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1712622712
transform 1 0 344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1712622712
transform 1 0 336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1712622712
transform 1 0 296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1712622712
transform 1 0 288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3469
timestamp 1712622712
transform 1 0 280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1712622712
transform 1 0 232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1712622712
transform 1 0 224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1712622712
transform 1 0 216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1712622712
transform 1 0 208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1712622712
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1712622712
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1712622712
transform 1 0 144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1712622712
transform 1 0 136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1712622712
transform 1 0 128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1712622712
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1712622712
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1712622712
transform 1 0 3424 0 1 970
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1712622712
transform 1 0 3392 0 1 970
box -8 -3 16 105
use FILL  FILL_3483
timestamp 1712622712
transform 1 0 3384 0 1 970
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1712622712
transform 1 0 3376 0 1 970
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1712622712
transform 1 0 3368 0 1 970
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1712622712
transform 1 0 3320 0 1 970
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1712622712
transform 1 0 3312 0 1 970
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1712622712
transform 1 0 3304 0 1 970
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1712622712
transform 1 0 3256 0 1 970
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1712622712
transform 1 0 3248 0 1 970
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1712622712
transform 1 0 3240 0 1 970
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1712622712
transform 1 0 3232 0 1 970
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1712622712
transform 1 0 3224 0 1 970
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1712622712
transform 1 0 3160 0 1 970
box -8 -3 16 105
use FILL  FILL_3495
timestamp 1712622712
transform 1 0 3152 0 1 970
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1712622712
transform 1 0 3144 0 1 970
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1712622712
transform 1 0 3040 0 1 970
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1712622712
transform 1 0 3032 0 1 970
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1712622712
transform 1 0 3024 0 1 970
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1712622712
transform 1 0 3016 0 1 970
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1712622712
transform 1 0 3008 0 1 970
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1712622712
transform 1 0 2952 0 1 970
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1712622712
transform 1 0 2944 0 1 970
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1712622712
transform 1 0 2936 0 1 970
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1712622712
transform 1 0 2896 0 1 970
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1712622712
transform 1 0 2888 0 1 970
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1712622712
transform 1 0 2880 0 1 970
box -8 -3 16 105
use FILL  FILL_3508
timestamp 1712622712
transform 1 0 2872 0 1 970
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1712622712
transform 1 0 2832 0 1 970
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1712622712
transform 1 0 2824 0 1 970
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1712622712
transform 1 0 2784 0 1 970
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1712622712
transform 1 0 2776 0 1 970
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1712622712
transform 1 0 2768 0 1 970
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1712622712
transform 1 0 2760 0 1 970
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1712622712
transform 1 0 2752 0 1 970
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1712622712
transform 1 0 2744 0 1 970
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1712622712
transform 1 0 2688 0 1 970
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1712622712
transform 1 0 2680 0 1 970
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1712622712
transform 1 0 2672 0 1 970
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1712622712
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1712622712
transform 1 0 2624 0 1 970
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1712622712
transform 1 0 2616 0 1 970
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1712622712
transform 1 0 2608 0 1 970
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1712622712
transform 1 0 2600 0 1 970
box -8 -3 16 105
use FILL  FILL_3525
timestamp 1712622712
transform 1 0 2552 0 1 970
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1712622712
transform 1 0 2544 0 1 970
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1712622712
transform 1 0 2536 0 1 970
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1712622712
transform 1 0 2528 0 1 970
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1712622712
transform 1 0 2496 0 1 970
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1712622712
transform 1 0 2488 0 1 970
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1712622712
transform 1 0 2480 0 1 970
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1712622712
transform 1 0 2432 0 1 970
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1712622712
transform 1 0 2424 0 1 970
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1712622712
transform 1 0 2416 0 1 970
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1712622712
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1712622712
transform 1 0 2360 0 1 970
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1712622712
transform 1 0 2352 0 1 970
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1712622712
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1712622712
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1712622712
transform 1 0 2296 0 1 970
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1712622712
transform 1 0 2288 0 1 970
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1712622712
transform 1 0 2280 0 1 970
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1712622712
transform 1 0 2272 0 1 970
box -8 -3 16 105
use FILL  FILL_3544
timestamp 1712622712
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1712622712
transform 1 0 2224 0 1 970
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1712622712
transform 1 0 2216 0 1 970
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1712622712
transform 1 0 2176 0 1 970
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1712622712
transform 1 0 2168 0 1 970
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1712622712
transform 1 0 2160 0 1 970
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1712622712
transform 1 0 2152 0 1 970
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1712622712
transform 1 0 2112 0 1 970
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1712622712
transform 1 0 2104 0 1 970
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1712622712
transform 1 0 2096 0 1 970
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1712622712
transform 1 0 2088 0 1 970
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1712622712
transform 1 0 2048 0 1 970
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1712622712
transform 1 0 2040 0 1 970
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1712622712
transform 1 0 2032 0 1 970
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1712622712
transform 1 0 2024 0 1 970
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1712622712
transform 1 0 2016 0 1 970
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1712622712
transform 1 0 1976 0 1 970
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1712622712
transform 1 0 1952 0 1 970
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1712622712
transform 1 0 1944 0 1 970
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1712622712
transform 1 0 1936 0 1 970
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1712622712
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1712622712
transform 1 0 1904 0 1 970
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1712622712
transform 1 0 1896 0 1 970
box -8 -3 16 105
use FILL  FILL_3567
timestamp 1712622712
transform 1 0 1856 0 1 970
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1712622712
transform 1 0 1848 0 1 970
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1712622712
transform 1 0 1840 0 1 970
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1712622712
transform 1 0 1832 0 1 970
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1712622712
transform 1 0 1800 0 1 970
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1712622712
transform 1 0 1792 0 1 970
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1712622712
transform 1 0 1784 0 1 970
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1712622712
transform 1 0 1744 0 1 970
box -8 -3 16 105
use FILL  FILL_3575
timestamp 1712622712
transform 1 0 1736 0 1 970
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1712622712
transform 1 0 1728 0 1 970
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1712622712
transform 1 0 1720 0 1 970
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1712622712
transform 1 0 1680 0 1 970
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1712622712
transform 1 0 1672 0 1 970
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1712622712
transform 1 0 1664 0 1 970
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1712622712
transform 1 0 1632 0 1 970
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1712622712
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1712622712
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1712622712
transform 1 0 1608 0 1 970
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1712622712
transform 1 0 1600 0 1 970
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1712622712
transform 1 0 1552 0 1 970
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1712622712
transform 1 0 1544 0 1 970
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1712622712
transform 1 0 1536 0 1 970
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1712622712
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1712622712
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1712622712
transform 1 0 1472 0 1 970
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1712622712
transform 1 0 1464 0 1 970
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1712622712
transform 1 0 1456 0 1 970
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1712622712
transform 1 0 1448 0 1 970
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1712622712
transform 1 0 1408 0 1 970
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1712622712
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1712622712
transform 1 0 1368 0 1 970
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1712622712
transform 1 0 1360 0 1 970
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1712622712
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1712622712
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1712622712
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1712622712
transform 1 0 1304 0 1 970
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1712622712
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1712622712
transform 1 0 1248 0 1 970
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1712622712
transform 1 0 1240 0 1 970
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1712622712
transform 1 0 1232 0 1 970
box -8 -3 16 105
use FILL  FILL_3607
timestamp 1712622712
transform 1 0 1224 0 1 970
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1712622712
transform 1 0 1192 0 1 970
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1712622712
transform 1 0 1184 0 1 970
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1712622712
transform 1 0 1176 0 1 970
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1712622712
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1712622712
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1712622712
transform 1 0 1120 0 1 970
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1712622712
transform 1 0 1080 0 1 970
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1712622712
transform 1 0 1072 0 1 970
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1712622712
transform 1 0 1064 0 1 970
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1712622712
transform 1 0 1056 0 1 970
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1712622712
transform 1 0 1016 0 1 970
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1712622712
transform 1 0 1008 0 1 970
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1712622712
transform 1 0 1000 0 1 970
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1712622712
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1712622712
transform 1 0 952 0 1 970
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1712622712
transform 1 0 944 0 1 970
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1712622712
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1712622712
transform 1 0 928 0 1 970
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1712622712
transform 1 0 904 0 1 970
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1712622712
transform 1 0 896 0 1 970
box -8 -3 16 105
use FILL  FILL_3628
timestamp 1712622712
transform 1 0 864 0 1 970
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1712622712
transform 1 0 856 0 1 970
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1712622712
transform 1 0 848 0 1 970
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1712622712
transform 1 0 808 0 1 970
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1712622712
transform 1 0 800 0 1 970
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1712622712
transform 1 0 792 0 1 970
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1712622712
transform 1 0 784 0 1 970
box -8 -3 16 105
use FILL  FILL_3635
timestamp 1712622712
transform 1 0 744 0 1 970
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1712622712
transform 1 0 736 0 1 970
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1712622712
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1712622712
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1712622712
transform 1 0 680 0 1 970
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1712622712
transform 1 0 672 0 1 970
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1712622712
transform 1 0 664 0 1 970
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1712622712
transform 1 0 656 0 1 970
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1712622712
transform 1 0 616 0 1 970
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1712622712
transform 1 0 608 0 1 970
box -8 -3 16 105
use FILL  FILL_3645
timestamp 1712622712
transform 1 0 600 0 1 970
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1712622712
transform 1 0 568 0 1 970
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1712622712
transform 1 0 560 0 1 970
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1712622712
transform 1 0 552 0 1 970
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1712622712
transform 1 0 544 0 1 970
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1712622712
transform 1 0 536 0 1 970
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1712622712
transform 1 0 480 0 1 970
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1712622712
transform 1 0 472 0 1 970
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1712622712
transform 1 0 464 0 1 970
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1712622712
transform 1 0 416 0 1 970
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1712622712
transform 1 0 408 0 1 970
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1712622712
transform 1 0 400 0 1 970
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1712622712
transform 1 0 392 0 1 970
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1712622712
transform 1 0 384 0 1 970
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1712622712
transform 1 0 376 0 1 970
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1712622712
transform 1 0 344 0 1 970
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1712622712
transform 1 0 304 0 1 970
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1712622712
transform 1 0 296 0 1 970
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1712622712
transform 1 0 288 0 1 970
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1712622712
transform 1 0 280 0 1 970
box -8 -3 16 105
use FILL  FILL_3665
timestamp 1712622712
transform 1 0 272 0 1 970
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1712622712
transform 1 0 240 0 1 970
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1712622712
transform 1 0 232 0 1 970
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1712622712
transform 1 0 224 0 1 970
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1712622712
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1712622712
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1712622712
transform 1 0 160 0 1 970
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1712622712
transform 1 0 152 0 1 970
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1712622712
transform 1 0 144 0 1 970
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1712622712
transform 1 0 136 0 1 970
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1712622712
transform 1 0 88 0 1 970
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1712622712
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_3677
timestamp 1712622712
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1712622712
transform 1 0 3424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1712622712
transform 1 0 3384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1712622712
transform 1 0 3376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1712622712
transform 1 0 3368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1712622712
transform 1 0 3360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1712622712
transform 1 0 3304 0 -1 970
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1712622712
transform 1 0 3296 0 -1 970
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1712622712
transform 1 0 3288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1712622712
transform 1 0 3264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1712622712
transform 1 0 3256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1712622712
transform 1 0 3248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1712622712
transform 1 0 3208 0 -1 970
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1712622712
transform 1 0 3160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1712622712
transform 1 0 3152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1712622712
transform 1 0 3144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1712622712
transform 1 0 3040 0 -1 970
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1712622712
transform 1 0 3032 0 -1 970
box -8 -3 16 105
use FILL  FILL_3695
timestamp 1712622712
transform 1 0 3024 0 -1 970
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1712622712
transform 1 0 3000 0 -1 970
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1712622712
transform 1 0 2976 0 -1 970
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1712622712
transform 1 0 2952 0 -1 970
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1712622712
transform 1 0 2944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1712622712
transform 1 0 2936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1712622712
transform 1 0 2896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1712622712
transform 1 0 2888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1712622712
transform 1 0 2880 0 -1 970
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1712622712
transform 1 0 2840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1712622712
transform 1 0 2832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1712622712
transform 1 0 2824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1712622712
transform 1 0 2784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1712622712
transform 1 0 2776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1712622712
transform 1 0 2768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1712622712
transform 1 0 2760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1712622712
transform 1 0 2752 0 -1 970
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1712622712
transform 1 0 2744 0 -1 970
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1712622712
transform 1 0 2688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1712622712
transform 1 0 2680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3715
timestamp 1712622712
transform 1 0 2672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1712622712
transform 1 0 2624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1712622712
transform 1 0 2616 0 -1 970
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1712622712
transform 1 0 2608 0 -1 970
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1712622712
transform 1 0 2600 0 -1 970
box -8 -3 16 105
use FILL  FILL_3720
timestamp 1712622712
transform 1 0 2552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1712622712
transform 1 0 2544 0 -1 970
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1712622712
transform 1 0 2536 0 -1 970
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1712622712
transform 1 0 2488 0 -1 970
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1712622712
transform 1 0 2480 0 -1 970
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1712622712
transform 1 0 2472 0 -1 970
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1712622712
transform 1 0 2464 0 -1 970
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1712622712
transform 1 0 2432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1712622712
transform 1 0 2424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1712622712
transform 1 0 2416 0 -1 970
box -8 -3 16 105
use FILL  FILL_3730
timestamp 1712622712
transform 1 0 2368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1712622712
transform 1 0 2360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1712622712
transform 1 0 2352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1712622712
transform 1 0 2344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1712622712
transform 1 0 2336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1712622712
transform 1 0 2328 0 -1 970
box -8 -3 16 105
use FILL  FILL_3736
timestamp 1712622712
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1712622712
transform 1 0 2256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1712622712
transform 1 0 2248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1712622712
transform 1 0 2240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1712622712
transform 1 0 2232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1712622712
transform 1 0 2224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1712622712
transform 1 0 2176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1712622712
transform 1 0 2144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1712622712
transform 1 0 2136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1712622712
transform 1 0 2128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1712622712
transform 1 0 2120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1712622712
transform 1 0 2112 0 -1 970
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1712622712
transform 1 0 2064 0 -1 970
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1712622712
transform 1 0 2056 0 -1 970
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1712622712
transform 1 0 2048 0 -1 970
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1712622712
transform 1 0 2016 0 -1 970
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1712622712
transform 1 0 2008 0 -1 970
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1712622712
transform 1 0 2000 0 -1 970
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1712622712
transform 1 0 1960 0 -1 970
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1712622712
transform 1 0 1952 0 -1 970
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1712622712
transform 1 0 1944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3757
timestamp 1712622712
transform 1 0 1936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1712622712
transform 1 0 1904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1712622712
transform 1 0 1896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1712622712
transform 1 0 1888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1712622712
transform 1 0 1848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1712622712
transform 1 0 1840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1712622712
transform 1 0 1832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1712622712
transform 1 0 1824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1712622712
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1712622712
transform 1 0 1776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1712622712
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3768
timestamp 1712622712
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1712622712
transform 1 0 1752 0 -1 970
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1712622712
transform 1 0 1744 0 -1 970
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1712622712
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1712622712
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1712622712
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1712622712
transform 1 0 1672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1712622712
transform 1 0 1664 0 -1 970
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1712622712
transform 1 0 1632 0 -1 970
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1712622712
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1712622712
transform 1 0 1616 0 -1 970
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1712622712
transform 1 0 1576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3780
timestamp 1712622712
transform 1 0 1568 0 -1 970
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1712622712
transform 1 0 1560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1712622712
transform 1 0 1552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1712622712
transform 1 0 1544 0 -1 970
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1712622712
transform 1 0 1536 0 -1 970
box -8 -3 16 105
use FILL  FILL_3785
timestamp 1712622712
transform 1 0 1496 0 -1 970
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1712622712
transform 1 0 1488 0 -1 970
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1712622712
transform 1 0 1480 0 -1 970
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1712622712
transform 1 0 1440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3789
timestamp 1712622712
transform 1 0 1432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1712622712
transform 1 0 1424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1712622712
transform 1 0 1416 0 -1 970
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1712622712
transform 1 0 1408 0 -1 970
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1712622712
transform 1 0 1360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1712622712
transform 1 0 1352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1712622712
transform 1 0 1344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1712622712
transform 1 0 1336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1712622712
transform 1 0 1328 0 -1 970
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1712622712
transform 1 0 1320 0 -1 970
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1712622712
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1712622712
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1712622712
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1712622712
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1712622712
transform 1 0 1232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1712622712
transform 1 0 1224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1712622712
transform 1 0 1184 0 -1 970
box -8 -3 16 105
use FILL  FILL_3806
timestamp 1712622712
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1712622712
transform 1 0 1136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1712622712
transform 1 0 1128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1712622712
transform 1 0 1120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1712622712
transform 1 0 1112 0 -1 970
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1712622712
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1712622712
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1712622712
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1712622712
transform 1 0 1040 0 -1 970
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1712622712
transform 1 0 1032 0 -1 970
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1712622712
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use FILL  FILL_3817
timestamp 1712622712
transform 1 0 1000 0 -1 970
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1712622712
transform 1 0 992 0 -1 970
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1712622712
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1712622712
transform 1 0 944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1712622712
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1712622712
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1712622712
transform 1 0 896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1712622712
transform 1 0 888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3825
timestamp 1712622712
transform 1 0 880 0 -1 970
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1712622712
transform 1 0 840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1712622712
transform 1 0 832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1712622712
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1712622712
transform 1 0 784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1712622712
transform 1 0 776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1712622712
transform 1 0 768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1712622712
transform 1 0 760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1712622712
transform 1 0 752 0 -1 970
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1712622712
transform 1 0 744 0 -1 970
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1712622712
transform 1 0 688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1712622712
transform 1 0 680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1712622712
transform 1 0 672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1712622712
transform 1 0 664 0 -1 970
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1712622712
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1712622712
transform 1 0 584 0 -1 970
box -8 -3 16 105
use FILL  FILL_3841
timestamp 1712622712
transform 1 0 576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1712622712
transform 1 0 568 0 -1 970
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1712622712
transform 1 0 560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1712622712
transform 1 0 552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1712622712
transform 1 0 504 0 -1 970
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1712622712
transform 1 0 496 0 -1 970
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1712622712
transform 1 0 488 0 -1 970
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1712622712
transform 1 0 480 0 -1 970
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1712622712
transform 1 0 440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1712622712
transform 1 0 432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1712622712
transform 1 0 392 0 -1 970
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1712622712
transform 1 0 384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1712622712
transform 1 0 376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1712622712
transform 1 0 336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1712622712
transform 1 0 328 0 -1 970
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1712622712
transform 1 0 320 0 -1 970
box -8 -3 16 105
use FILL  FILL_3857
timestamp 1712622712
transform 1 0 288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1712622712
transform 1 0 280 0 -1 970
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1712622712
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1712622712
transform 1 0 264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1712622712
transform 1 0 240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1712622712
transform 1 0 208 0 -1 970
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1712622712
transform 1 0 200 0 -1 970
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1712622712
transform 1 0 192 0 -1 970
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1712622712
transform 1 0 184 0 -1 970
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1712622712
transform 1 0 176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1712622712
transform 1 0 168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1712622712
transform 1 0 128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1712622712
transform 1 0 120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1712622712
transform 1 0 88 0 -1 970
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1712622712
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1712622712
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1712622712
transform 1 0 3424 0 1 770
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1712622712
transform 1 0 3368 0 1 770
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1712622712
transform 1 0 3360 0 1 770
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1712622712
transform 1 0 3352 0 1 770
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1712622712
transform 1 0 3344 0 1 770
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1712622712
transform 1 0 3336 0 1 770
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1712622712
transform 1 0 3264 0 1 770
box -8 -3 16 105
use FILL  FILL_3880
timestamp 1712622712
transform 1 0 3256 0 1 770
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1712622712
transform 1 0 3248 0 1 770
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1712622712
transform 1 0 3240 0 1 770
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1712622712
transform 1 0 3232 0 1 770
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1712622712
transform 1 0 3224 0 1 770
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1712622712
transform 1 0 3176 0 1 770
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1712622712
transform 1 0 3168 0 1 770
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1712622712
transform 1 0 3160 0 1 770
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1712622712
transform 1 0 3072 0 1 770
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1712622712
transform 1 0 3064 0 1 770
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1712622712
transform 1 0 2960 0 1 770
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1712622712
transform 1 0 2952 0 1 770
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1712622712
transform 1 0 2944 0 1 770
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1712622712
transform 1 0 2856 0 1 770
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1712622712
transform 1 0 2848 0 1 770
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1712622712
transform 1 0 2840 0 1 770
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1712622712
transform 1 0 2736 0 1 770
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1712622712
transform 1 0 2728 0 1 770
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1712622712
transform 1 0 2720 0 1 770
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1712622712
transform 1 0 2712 0 1 770
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1712622712
transform 1 0 2664 0 1 770
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1712622712
transform 1 0 2656 0 1 770
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1712622712
transform 1 0 2648 0 1 770
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1712622712
transform 1 0 2640 0 1 770
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1712622712
transform 1 0 2632 0 1 770
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1712622712
transform 1 0 2600 0 1 770
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1712622712
transform 1 0 2576 0 1 770
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1712622712
transform 1 0 2568 0 1 770
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1712622712
transform 1 0 2560 0 1 770
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1712622712
transform 1 0 2552 0 1 770
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1712622712
transform 1 0 2528 0 1 770
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1712622712
transform 1 0 2520 0 1 770
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1712622712
transform 1 0 2480 0 1 770
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1712622712
transform 1 0 2472 0 1 770
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1712622712
transform 1 0 2464 0 1 770
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1712622712
transform 1 0 2456 0 1 770
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1712622712
transform 1 0 2448 0 1 770
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1712622712
transform 1 0 2440 0 1 770
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1712622712
transform 1 0 2432 0 1 770
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1712622712
transform 1 0 2376 0 1 770
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1712622712
transform 1 0 2368 0 1 770
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1712622712
transform 1 0 2360 0 1 770
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1712622712
transform 1 0 2352 0 1 770
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1712622712
transform 1 0 2320 0 1 770
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1712622712
transform 1 0 2312 0 1 770
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1712622712
transform 1 0 2304 0 1 770
box -8 -3 16 105
use FILL  FILL_3926
timestamp 1712622712
transform 1 0 2264 0 1 770
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1712622712
transform 1 0 2256 0 1 770
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1712622712
transform 1 0 2248 0 1 770
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1712622712
transform 1 0 2240 0 1 770
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1712622712
transform 1 0 2208 0 1 770
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1712622712
transform 1 0 2200 0 1 770
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1712622712
transform 1 0 2192 0 1 770
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1712622712
transform 1 0 2184 0 1 770
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1712622712
transform 1 0 2144 0 1 770
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1712622712
transform 1 0 2136 0 1 770
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1712622712
transform 1 0 2128 0 1 770
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1712622712
transform 1 0 2096 0 1 770
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1712622712
transform 1 0 2088 0 1 770
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1712622712
transform 1 0 2080 0 1 770
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1712622712
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1712622712
transform 1 0 2064 0 1 770
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1712622712
transform 1 0 2016 0 1 770
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1712622712
transform 1 0 2008 0 1 770
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1712622712
transform 1 0 2000 0 1 770
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1712622712
transform 1 0 1992 0 1 770
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1712622712
transform 1 0 1952 0 1 770
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1712622712
transform 1 0 1944 0 1 770
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1712622712
transform 1 0 1936 0 1 770
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1712622712
transform 1 0 1896 0 1 770
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1712622712
transform 1 0 1888 0 1 770
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1712622712
transform 1 0 1880 0 1 770
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1712622712
transform 1 0 1872 0 1 770
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1712622712
transform 1 0 1864 0 1 770
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1712622712
transform 1 0 1824 0 1 770
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1712622712
transform 1 0 1816 0 1 770
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1712622712
transform 1 0 1808 0 1 770
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1712622712
transform 1 0 1800 0 1 770
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1712622712
transform 1 0 1768 0 1 770
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1712622712
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1712622712
transform 1 0 1728 0 1 770
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1712622712
transform 1 0 1720 0 1 770
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1712622712
transform 1 0 1712 0 1 770
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1712622712
transform 1 0 1704 0 1 770
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1712622712
transform 1 0 1696 0 1 770
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1712622712
transform 1 0 1688 0 1 770
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1712622712
transform 1 0 1648 0 1 770
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1712622712
transform 1 0 1640 0 1 770
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1712622712
transform 1 0 1632 0 1 770
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1712622712
transform 1 0 1592 0 1 770
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1712622712
transform 1 0 1584 0 1 770
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1712622712
transform 1 0 1576 0 1 770
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1712622712
transform 1 0 1568 0 1 770
box -8 -3 16 105
use FILL  FILL_3973
timestamp 1712622712
transform 1 0 1560 0 1 770
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1712622712
transform 1 0 1552 0 1 770
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1712622712
transform 1 0 1504 0 1 770
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1712622712
transform 1 0 1496 0 1 770
box -8 -3 16 105
use FILL  FILL_3977
timestamp 1712622712
transform 1 0 1488 0 1 770
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1712622712
transform 1 0 1480 0 1 770
box -8 -3 16 105
use FILL  FILL_3979
timestamp 1712622712
transform 1 0 1440 0 1 770
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1712622712
transform 1 0 1432 0 1 770
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1712622712
transform 1 0 1424 0 1 770
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1712622712
transform 1 0 1416 0 1 770
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1712622712
transform 1 0 1368 0 1 770
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1712622712
transform 1 0 1360 0 1 770
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1712622712
transform 1 0 1352 0 1 770
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1712622712
transform 1 0 1344 0 1 770
box -8 -3 16 105
use FILL  FILL_3987
timestamp 1712622712
transform 1 0 1336 0 1 770
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1712622712
transform 1 0 1328 0 1 770
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1712622712
transform 1 0 1280 0 1 770
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1712622712
transform 1 0 1272 0 1 770
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1712622712
transform 1 0 1264 0 1 770
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1712622712
transform 1 0 1232 0 1 770
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1712622712
transform 1 0 1224 0 1 770
box -8 -3 16 105
use FILL  FILL_3994
timestamp 1712622712
transform 1 0 1216 0 1 770
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1712622712
transform 1 0 1168 0 1 770
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1712622712
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_3997
timestamp 1712622712
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1712622712
transform 1 0 1144 0 1 770
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1712622712
transform 1 0 1136 0 1 770
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1712622712
transform 1 0 1128 0 1 770
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1712622712
transform 1 0 1080 0 1 770
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1712622712
transform 1 0 1056 0 1 770
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1712622712
transform 1 0 1048 0 1 770
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1712622712
transform 1 0 1040 0 1 770
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1712622712
transform 1 0 1032 0 1 770
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1712622712
transform 1 0 992 0 1 770
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1712622712
transform 1 0 984 0 1 770
box -8 -3 16 105
use FILL  FILL_4008
timestamp 1712622712
transform 1 0 976 0 1 770
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1712622712
transform 1 0 936 0 1 770
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1712622712
transform 1 0 928 0 1 770
box -8 -3 16 105
use FILL  FILL_4011
timestamp 1712622712
transform 1 0 920 0 1 770
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1712622712
transform 1 0 912 0 1 770
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1712622712
transform 1 0 904 0 1 770
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1712622712
transform 1 0 864 0 1 770
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1712622712
transform 1 0 856 0 1 770
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1712622712
transform 1 0 848 0 1 770
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1712622712
transform 1 0 808 0 1 770
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1712622712
transform 1 0 800 0 1 770
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1712622712
transform 1 0 792 0 1 770
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1712622712
transform 1 0 784 0 1 770
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1712622712
transform 1 0 752 0 1 770
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1712622712
transform 1 0 744 0 1 770
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1712622712
transform 1 0 736 0 1 770
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1712622712
transform 1 0 696 0 1 770
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1712622712
transform 1 0 688 0 1 770
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1712622712
transform 1 0 680 0 1 770
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1712622712
transform 1 0 672 0 1 770
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1712622712
transform 1 0 632 0 1 770
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1712622712
transform 1 0 624 0 1 770
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1712622712
transform 1 0 616 0 1 770
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1712622712
transform 1 0 608 0 1 770
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1712622712
transform 1 0 600 0 1 770
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1712622712
transform 1 0 552 0 1 770
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1712622712
transform 1 0 544 0 1 770
box -8 -3 16 105
use FILL  FILL_4035
timestamp 1712622712
transform 1 0 536 0 1 770
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1712622712
transform 1 0 528 0 1 770
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1712622712
transform 1 0 480 0 1 770
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1712622712
transform 1 0 472 0 1 770
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1712622712
transform 1 0 464 0 1 770
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1712622712
transform 1 0 456 0 1 770
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1712622712
transform 1 0 448 0 1 770
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1712622712
transform 1 0 400 0 1 770
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1712622712
transform 1 0 392 0 1 770
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1712622712
transform 1 0 384 0 1 770
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1712622712
transform 1 0 376 0 1 770
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1712622712
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1712622712
transform 1 0 320 0 1 770
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1712622712
transform 1 0 312 0 1 770
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1712622712
transform 1 0 304 0 1 770
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1712622712
transform 1 0 296 0 1 770
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1712622712
transform 1 0 256 0 1 770
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1712622712
transform 1 0 248 0 1 770
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1712622712
transform 1 0 240 0 1 770
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1712622712
transform 1 0 232 0 1 770
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1712622712
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1712622712
transform 1 0 176 0 1 770
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1712622712
transform 1 0 168 0 1 770
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1712622712
transform 1 0 160 0 1 770
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1712622712
transform 1 0 152 0 1 770
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1712622712
transform 1 0 144 0 1 770
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1712622712
transform 1 0 120 0 1 770
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1712622712
transform 1 0 88 0 1 770
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1712622712
transform 1 0 80 0 1 770
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1712622712
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1712622712
transform 1 0 3424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1712622712
transform 1 0 3400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1712622712
transform 1 0 3392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1712622712
transform 1 0 3384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1712622712
transform 1 0 3376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1712622712
transform 1 0 3368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1712622712
transform 1 0 3360 0 -1 770
box -8 -3 16 105
use FILL  FILL_4072
timestamp 1712622712
transform 1 0 3352 0 -1 770
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1712622712
transform 1 0 3344 0 -1 770
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1712622712
transform 1 0 3280 0 -1 770
box -8 -3 16 105
use FILL  FILL_4075
timestamp 1712622712
transform 1 0 3272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1712622712
transform 1 0 3264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1712622712
transform 1 0 3256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4078
timestamp 1712622712
transform 1 0 3168 0 -1 770
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1712622712
transform 1 0 3160 0 -1 770
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1712622712
transform 1 0 3152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1712622712
transform 1 0 3112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1712622712
transform 1 0 3104 0 -1 770
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1712622712
transform 1 0 3096 0 -1 770
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1712622712
transform 1 0 3088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1712622712
transform 1 0 3024 0 -1 770
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1712622712
transform 1 0 3016 0 -1 770
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1712622712
transform 1 0 3008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1712622712
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1712622712
transform 1 0 2952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1712622712
transform 1 0 2944 0 -1 770
box -8 -3 16 105
use FILL  FILL_4091
timestamp 1712622712
transform 1 0 2880 0 -1 770
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1712622712
transform 1 0 2872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1712622712
transform 1 0 2768 0 -1 770
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1712622712
transform 1 0 2760 0 -1 770
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1712622712
transform 1 0 2752 0 -1 770
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1712622712
transform 1 0 2744 0 -1 770
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1712622712
transform 1 0 2736 0 -1 770
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1712622712
transform 1 0 2648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1712622712
transform 1 0 2640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1712622712
transform 1 0 2632 0 -1 770
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1712622712
transform 1 0 2624 0 -1 770
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1712622712
transform 1 0 2592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4103
timestamp 1712622712
transform 1 0 2584 0 -1 770
box -8 -3 16 105
use FILL  FILL_4104
timestamp 1712622712
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1712622712
transform 1 0 2544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1712622712
transform 1 0 2520 0 -1 770
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1712622712
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1712622712
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1712622712
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_4110
timestamp 1712622712
transform 1 0 2448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1712622712
transform 1 0 2440 0 -1 770
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1712622712
transform 1 0 2432 0 -1 770
box -8 -3 16 105
use FILL  FILL_4113
timestamp 1712622712
transform 1 0 2424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1712622712
transform 1 0 2376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1712622712
transform 1 0 2368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1712622712
transform 1 0 2360 0 -1 770
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1712622712
transform 1 0 2352 0 -1 770
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1712622712
transform 1 0 2344 0 -1 770
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1712622712
transform 1 0 2296 0 -1 770
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1712622712
transform 1 0 2288 0 -1 770
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1712622712
transform 1 0 2280 0 -1 770
box -8 -3 16 105
use FILL  FILL_4122
timestamp 1712622712
transform 1 0 2272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1712622712
transform 1 0 2224 0 -1 770
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1712622712
transform 1 0 2216 0 -1 770
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1712622712
transform 1 0 2208 0 -1 770
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1712622712
transform 1 0 2200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1712622712
transform 1 0 2152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1712622712
transform 1 0 2144 0 -1 770
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1712622712
transform 1 0 2136 0 -1 770
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1712622712
transform 1 0 2128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1712622712
transform 1 0 2088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1712622712
transform 1 0 2080 0 -1 770
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1712622712
transform 1 0 2072 0 -1 770
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1712622712
transform 1 0 2064 0 -1 770
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1712622712
transform 1 0 2008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1712622712
transform 1 0 2000 0 -1 770
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1712622712
transform 1 0 1992 0 -1 770
box -8 -3 16 105
use FILL  FILL_4138
timestamp 1712622712
transform 1 0 1984 0 -1 770
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1712622712
transform 1 0 1976 0 -1 770
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1712622712
transform 1 0 1936 0 -1 770
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1712622712
transform 1 0 1928 0 -1 770
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1712622712
transform 1 0 1920 0 -1 770
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1712622712
transform 1 0 1888 0 -1 770
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1712622712
transform 1 0 1880 0 -1 770
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1712622712
transform 1 0 1872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1712622712
transform 1 0 1848 0 -1 770
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1712622712
transform 1 0 1840 0 -1 770
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1712622712
transform 1 0 1800 0 -1 770
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1712622712
transform 1 0 1792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1712622712
transform 1 0 1784 0 -1 770
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1712622712
transform 1 0 1760 0 -1 770
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1712622712
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1712622712
transform 1 0 1744 0 -1 770
box -8 -3 16 105
use FILL  FILL_4154
timestamp 1712622712
transform 1 0 1704 0 -1 770
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1712622712
transform 1 0 1696 0 -1 770
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1712622712
transform 1 0 1688 0 -1 770
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1712622712
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1712622712
transform 1 0 1640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1712622712
transform 1 0 1632 0 -1 770
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1712622712
transform 1 0 1624 0 -1 770
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1712622712
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1712622712
transform 1 0 1560 0 -1 770
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1712622712
transform 1 0 1552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1712622712
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4165
timestamp 1712622712
transform 1 0 1536 0 -1 770
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1712622712
transform 1 0 1504 0 -1 770
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1712622712
transform 1 0 1496 0 -1 770
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1712622712
transform 1 0 1488 0 -1 770
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1712622712
transform 1 0 1448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1712622712
transform 1 0 1440 0 -1 770
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1712622712
transform 1 0 1432 0 -1 770
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1712622712
transform 1 0 1424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1712622712
transform 1 0 1384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1712622712
transform 1 0 1376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1712622712
transform 1 0 1368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1712622712
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4177
timestamp 1712622712
transform 1 0 1320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1712622712
transform 1 0 1312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1712622712
transform 1 0 1304 0 -1 770
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1712622712
transform 1 0 1264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1712622712
transform 1 0 1256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1712622712
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1712622712
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1712622712
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1712622712
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4186
timestamp 1712622712
transform 1 0 1192 0 -1 770
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1712622712
transform 1 0 1184 0 -1 770
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1712622712
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1712622712
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1712622712
transform 1 0 1104 0 -1 770
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1712622712
transform 1 0 1096 0 -1 770
box -8 -3 16 105
use FILL  FILL_4192
timestamp 1712622712
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1712622712
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1712622712
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1712622712
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1712622712
transform 1 0 1000 0 -1 770
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1712622712
transform 1 0 992 0 -1 770
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1712622712
transform 1 0 984 0 -1 770
box -8 -3 16 105
use FILL  FILL_4199
timestamp 1712622712
transform 1 0 976 0 -1 770
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1712622712
transform 1 0 968 0 -1 770
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1712622712
transform 1 0 928 0 -1 770
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1712622712
transform 1 0 896 0 -1 770
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1712622712
transform 1 0 888 0 -1 770
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1712622712
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1712622712
transform 1 0 872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1712622712
transform 1 0 848 0 -1 770
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1712622712
transform 1 0 840 0 -1 770
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1712622712
transform 1 0 832 0 -1 770
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1712622712
transform 1 0 784 0 -1 770
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1712622712
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4211
timestamp 1712622712
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1712622712
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1712622712
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1712622712
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1712622712
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1712622712
transform 1 0 704 0 -1 770
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1712622712
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1712622712
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1712622712
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1712622712
transform 1 0 592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4221
timestamp 1712622712
transform 1 0 584 0 -1 770
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1712622712
transform 1 0 576 0 -1 770
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1712622712
transform 1 0 568 0 -1 770
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1712622712
transform 1 0 536 0 -1 770
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1712622712
transform 1 0 528 0 -1 770
box -8 -3 16 105
use FILL  FILL_4226
timestamp 1712622712
transform 1 0 520 0 -1 770
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1712622712
transform 1 0 472 0 -1 770
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1712622712
transform 1 0 464 0 -1 770
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1712622712
transform 1 0 456 0 -1 770
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1712622712
transform 1 0 424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1712622712
transform 1 0 416 0 -1 770
box -8 -3 16 105
use FILL  FILL_4232
timestamp 1712622712
transform 1 0 376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1712622712
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1712622712
transform 1 0 360 0 -1 770
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1712622712
transform 1 0 352 0 -1 770
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1712622712
transform 1 0 320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1712622712
transform 1 0 312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1712622712
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1712622712
transform 1 0 264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1712622712
transform 1 0 256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1712622712
transform 1 0 248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1712622712
transform 1 0 184 0 -1 770
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1712622712
transform 1 0 176 0 -1 770
box -8 -3 16 105
use FILL  FILL_4244
timestamp 1712622712
transform 1 0 168 0 -1 770
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1712622712
transform 1 0 160 0 -1 770
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1712622712
transform 1 0 152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1712622712
transform 1 0 144 0 -1 770
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1712622712
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1712622712
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1712622712
transform 1 0 3424 0 1 570
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1712622712
transform 1 0 3416 0 1 570
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1712622712
transform 1 0 3368 0 1 570
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1712622712
transform 1 0 3360 0 1 570
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1712622712
transform 1 0 3352 0 1 570
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1712622712
transform 1 0 3344 0 1 570
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1712622712
transform 1 0 3304 0 1 570
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1712622712
transform 1 0 3264 0 1 570
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1712622712
transform 1 0 3256 0 1 570
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1712622712
transform 1 0 3248 0 1 570
box -8 -3 16 105
use FILL  FILL_4260
timestamp 1712622712
transform 1 0 3240 0 1 570
box -8 -3 16 105
use FILL  FILL_4261
timestamp 1712622712
transform 1 0 3232 0 1 570
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1712622712
transform 1 0 3224 0 1 570
box -8 -3 16 105
use FILL  FILL_4263
timestamp 1712622712
transform 1 0 3192 0 1 570
box -8 -3 16 105
use FILL  FILL_4264
timestamp 1712622712
transform 1 0 3184 0 1 570
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1712622712
transform 1 0 3144 0 1 570
box -8 -3 16 105
use FILL  FILL_4266
timestamp 1712622712
transform 1 0 3136 0 1 570
box -8 -3 16 105
use FILL  FILL_4267
timestamp 1712622712
transform 1 0 3128 0 1 570
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1712622712
transform 1 0 3120 0 1 570
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1712622712
transform 1 0 3112 0 1 570
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1712622712
transform 1 0 3064 0 1 570
box -8 -3 16 105
use FILL  FILL_4271
timestamp 1712622712
transform 1 0 3056 0 1 570
box -8 -3 16 105
use FILL  FILL_4272
timestamp 1712622712
transform 1 0 3048 0 1 570
box -8 -3 16 105
use FILL  FILL_4273
timestamp 1712622712
transform 1 0 3024 0 1 570
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1712622712
transform 1 0 3016 0 1 570
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1712622712
transform 1 0 3008 0 1 570
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1712622712
transform 1 0 2976 0 1 570
box -8 -3 16 105
use FILL  FILL_4277
timestamp 1712622712
transform 1 0 2968 0 1 570
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1712622712
transform 1 0 2960 0 1 570
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1712622712
transform 1 0 2952 0 1 570
box -8 -3 16 105
use FILL  FILL_4280
timestamp 1712622712
transform 1 0 2904 0 1 570
box -8 -3 16 105
use FILL  FILL_4281
timestamp 1712622712
transform 1 0 2896 0 1 570
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1712622712
transform 1 0 2888 0 1 570
box -8 -3 16 105
use FILL  FILL_4283
timestamp 1712622712
transform 1 0 2880 0 1 570
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1712622712
transform 1 0 2816 0 1 570
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1712622712
transform 1 0 2808 0 1 570
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1712622712
transform 1 0 2800 0 1 570
box -8 -3 16 105
use FILL  FILL_4287
timestamp 1712622712
transform 1 0 2792 0 1 570
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1712622712
transform 1 0 2768 0 1 570
box -8 -3 16 105
use FILL  FILL_4289
timestamp 1712622712
transform 1 0 2736 0 1 570
box -8 -3 16 105
use FILL  FILL_4290
timestamp 1712622712
transform 1 0 2728 0 1 570
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1712622712
transform 1 0 2720 0 1 570
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1712622712
transform 1 0 2688 0 1 570
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1712622712
transform 1 0 2680 0 1 570
box -8 -3 16 105
use FILL  FILL_4294
timestamp 1712622712
transform 1 0 2672 0 1 570
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1712622712
transform 1 0 2664 0 1 570
box -8 -3 16 105
use FILL  FILL_4296
timestamp 1712622712
transform 1 0 2656 0 1 570
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1712622712
transform 1 0 2608 0 1 570
box -8 -3 16 105
use FILL  FILL_4298
timestamp 1712622712
transform 1 0 2600 0 1 570
box -8 -3 16 105
use FILL  FILL_4299
timestamp 1712622712
transform 1 0 2592 0 1 570
box -8 -3 16 105
use FILL  FILL_4300
timestamp 1712622712
transform 1 0 2584 0 1 570
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1712622712
transform 1 0 2576 0 1 570
box -8 -3 16 105
use FILL  FILL_4302
timestamp 1712622712
transform 1 0 2528 0 1 570
box -8 -3 16 105
use FILL  FILL_4303
timestamp 1712622712
transform 1 0 2520 0 1 570
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1712622712
transform 1 0 2512 0 1 570
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1712622712
transform 1 0 2480 0 1 570
box -8 -3 16 105
use FILL  FILL_4306
timestamp 1712622712
transform 1 0 2472 0 1 570
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1712622712
transform 1 0 2464 0 1 570
box -8 -3 16 105
use FILL  FILL_4308
timestamp 1712622712
transform 1 0 2424 0 1 570
box -8 -3 16 105
use FILL  FILL_4309
timestamp 1712622712
transform 1 0 2416 0 1 570
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1712622712
transform 1 0 2408 0 1 570
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1712622712
transform 1 0 2368 0 1 570
box -8 -3 16 105
use FILL  FILL_4312
timestamp 1712622712
transform 1 0 2360 0 1 570
box -8 -3 16 105
use FILL  FILL_4313
timestamp 1712622712
transform 1 0 2352 0 1 570
box -8 -3 16 105
use FILL  FILL_4314
timestamp 1712622712
transform 1 0 2344 0 1 570
box -8 -3 16 105
use FILL  FILL_4315
timestamp 1712622712
transform 1 0 2336 0 1 570
box -8 -3 16 105
use FILL  FILL_4316
timestamp 1712622712
transform 1 0 2328 0 1 570
box -8 -3 16 105
use FILL  FILL_4317
timestamp 1712622712
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_4318
timestamp 1712622712
transform 1 0 2256 0 1 570
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1712622712
transform 1 0 2248 0 1 570
box -8 -3 16 105
use FILL  FILL_4320
timestamp 1712622712
transform 1 0 2240 0 1 570
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1712622712
transform 1 0 2232 0 1 570
box -8 -3 16 105
use FILL  FILL_4322
timestamp 1712622712
transform 1 0 2184 0 1 570
box -8 -3 16 105
use FILL  FILL_4323
timestamp 1712622712
transform 1 0 2176 0 1 570
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1712622712
transform 1 0 2168 0 1 570
box -8 -3 16 105
use FILL  FILL_4325
timestamp 1712622712
transform 1 0 2136 0 1 570
box -8 -3 16 105
use FILL  FILL_4326
timestamp 1712622712
transform 1 0 2128 0 1 570
box -8 -3 16 105
use FILL  FILL_4327
timestamp 1712622712
transform 1 0 2120 0 1 570
box -8 -3 16 105
use FILL  FILL_4328
timestamp 1712622712
transform 1 0 2088 0 1 570
box -8 -3 16 105
use FILL  FILL_4329
timestamp 1712622712
transform 1 0 2080 0 1 570
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1712622712
transform 1 0 2072 0 1 570
box -8 -3 16 105
use FILL  FILL_4331
timestamp 1712622712
transform 1 0 2032 0 1 570
box -8 -3 16 105
use FILL  FILL_4332
timestamp 1712622712
transform 1 0 2024 0 1 570
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1712622712
transform 1 0 2016 0 1 570
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1712622712
transform 1 0 2008 0 1 570
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1712622712
transform 1 0 1968 0 1 570
box -8 -3 16 105
use FILL  FILL_4336
timestamp 1712622712
transform 1 0 1960 0 1 570
box -8 -3 16 105
use FILL  FILL_4337
timestamp 1712622712
transform 1 0 1952 0 1 570
box -8 -3 16 105
use FILL  FILL_4338
timestamp 1712622712
transform 1 0 1920 0 1 570
box -8 -3 16 105
use FILL  FILL_4339
timestamp 1712622712
transform 1 0 1912 0 1 570
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1712622712
transform 1 0 1904 0 1 570
box -8 -3 16 105
use FILL  FILL_4341
timestamp 1712622712
transform 1 0 1896 0 1 570
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1712622712
transform 1 0 1864 0 1 570
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1712622712
transform 1 0 1840 0 1 570
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1712622712
transform 1 0 1832 0 1 570
box -8 -3 16 105
use FILL  FILL_4345
timestamp 1712622712
transform 1 0 1824 0 1 570
box -8 -3 16 105
use FILL  FILL_4346
timestamp 1712622712
transform 1 0 1816 0 1 570
box -8 -3 16 105
use FILL  FILL_4347
timestamp 1712622712
transform 1 0 1808 0 1 570
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1712622712
transform 1 0 1800 0 1 570
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1712622712
transform 1 0 1744 0 1 570
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1712622712
transform 1 0 1736 0 1 570
box -8 -3 16 105
use FILL  FILL_4351
timestamp 1712622712
transform 1 0 1728 0 1 570
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1712622712
transform 1 0 1688 0 1 570
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1712622712
transform 1 0 1680 0 1 570
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1712622712
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_4355
timestamp 1712622712
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_4356
timestamp 1712622712
transform 1 0 1624 0 1 570
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1712622712
transform 1 0 1592 0 1 570
box -8 -3 16 105
use FILL  FILL_4358
timestamp 1712622712
transform 1 0 1584 0 1 570
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1712622712
transform 1 0 1576 0 1 570
box -8 -3 16 105
use FILL  FILL_4360
timestamp 1712622712
transform 1 0 1568 0 1 570
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1712622712
transform 1 0 1560 0 1 570
box -8 -3 16 105
use FILL  FILL_4362
timestamp 1712622712
transform 1 0 1504 0 1 570
box -8 -3 16 105
use FILL  FILL_4363
timestamp 1712622712
transform 1 0 1496 0 1 570
box -8 -3 16 105
use FILL  FILL_4364
timestamp 1712622712
transform 1 0 1488 0 1 570
box -8 -3 16 105
use FILL  FILL_4365
timestamp 1712622712
transform 1 0 1480 0 1 570
box -8 -3 16 105
use FILL  FILL_4366
timestamp 1712622712
transform 1 0 1472 0 1 570
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1712622712
transform 1 0 1416 0 1 570
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1712622712
transform 1 0 1408 0 1 570
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1712622712
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_4370
timestamp 1712622712
transform 1 0 1392 0 1 570
box -8 -3 16 105
use FILL  FILL_4371
timestamp 1712622712
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_4372
timestamp 1712622712
transform 1 0 1312 0 1 570
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1712622712
transform 1 0 1304 0 1 570
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1712622712
transform 1 0 1296 0 1 570
box -8 -3 16 105
use FILL  FILL_4375
timestamp 1712622712
transform 1 0 1288 0 1 570
box -8 -3 16 105
use FILL  FILL_4376
timestamp 1712622712
transform 1 0 1280 0 1 570
box -8 -3 16 105
use FILL  FILL_4377
timestamp 1712622712
transform 1 0 1240 0 1 570
box -8 -3 16 105
use FILL  FILL_4378
timestamp 1712622712
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_4379
timestamp 1712622712
transform 1 0 1192 0 1 570
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1712622712
transform 1 0 1184 0 1 570
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1712622712
transform 1 0 1176 0 1 570
box -8 -3 16 105
use FILL  FILL_4382
timestamp 1712622712
transform 1 0 1144 0 1 570
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1712622712
transform 1 0 1136 0 1 570
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1712622712
transform 1 0 1112 0 1 570
box -8 -3 16 105
use FILL  FILL_4385
timestamp 1712622712
transform 1 0 1072 0 1 570
box -8 -3 16 105
use FILL  FILL_4386
timestamp 1712622712
transform 1 0 1064 0 1 570
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1712622712
transform 1 0 1024 0 1 570
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1712622712
transform 1 0 1016 0 1 570
box -8 -3 16 105
use FILL  FILL_4389
timestamp 1712622712
transform 1 0 1008 0 1 570
box -8 -3 16 105
use FILL  FILL_4390
timestamp 1712622712
transform 1 0 968 0 1 570
box -8 -3 16 105
use FILL  FILL_4391
timestamp 1712622712
transform 1 0 960 0 1 570
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1712622712
transform 1 0 952 0 1 570
box -8 -3 16 105
use FILL  FILL_4393
timestamp 1712622712
transform 1 0 912 0 1 570
box -8 -3 16 105
use FILL  FILL_4394
timestamp 1712622712
transform 1 0 904 0 1 570
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1712622712
transform 1 0 896 0 1 570
box -8 -3 16 105
use FILL  FILL_4396
timestamp 1712622712
transform 1 0 856 0 1 570
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1712622712
transform 1 0 848 0 1 570
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1712622712
transform 1 0 840 0 1 570
box -8 -3 16 105
use FILL  FILL_4399
timestamp 1712622712
transform 1 0 832 0 1 570
box -8 -3 16 105
use FILL  FILL_4400
timestamp 1712622712
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1712622712
transform 1 0 784 0 1 570
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1712622712
transform 1 0 776 0 1 570
box -8 -3 16 105
use FILL  FILL_4403
timestamp 1712622712
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_4404
timestamp 1712622712
transform 1 0 744 0 1 570
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1712622712
transform 1 0 704 0 1 570
box -8 -3 16 105
use FILL  FILL_4406
timestamp 1712622712
transform 1 0 696 0 1 570
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1712622712
transform 1 0 688 0 1 570
box -8 -3 16 105
use FILL  FILL_4408
timestamp 1712622712
transform 1 0 680 0 1 570
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1712622712
transform 1 0 640 0 1 570
box -8 -3 16 105
use FILL  FILL_4410
timestamp 1712622712
transform 1 0 632 0 1 570
box -8 -3 16 105
use FILL  FILL_4411
timestamp 1712622712
transform 1 0 624 0 1 570
box -8 -3 16 105
use FILL  FILL_4412
timestamp 1712622712
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_4413
timestamp 1712622712
transform 1 0 576 0 1 570
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1712622712
transform 1 0 568 0 1 570
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1712622712
transform 1 0 560 0 1 570
box -8 -3 16 105
use FILL  FILL_4416
timestamp 1712622712
transform 1 0 520 0 1 570
box -8 -3 16 105
use FILL  FILL_4417
timestamp 1712622712
transform 1 0 512 0 1 570
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1712622712
transform 1 0 504 0 1 570
box -8 -3 16 105
use FILL  FILL_4419
timestamp 1712622712
transform 1 0 496 0 1 570
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1712622712
transform 1 0 488 0 1 570
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1712622712
transform 1 0 480 0 1 570
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1712622712
transform 1 0 416 0 1 570
box -8 -3 16 105
use FILL  FILL_4423
timestamp 1712622712
transform 1 0 408 0 1 570
box -8 -3 16 105
use FILL  FILL_4424
timestamp 1712622712
transform 1 0 400 0 1 570
box -8 -3 16 105
use FILL  FILL_4425
timestamp 1712622712
transform 1 0 392 0 1 570
box -8 -3 16 105
use FILL  FILL_4426
timestamp 1712622712
transform 1 0 384 0 1 570
box -8 -3 16 105
use FILL  FILL_4427
timestamp 1712622712
transform 1 0 376 0 1 570
box -8 -3 16 105
use FILL  FILL_4428
timestamp 1712622712
transform 1 0 368 0 1 570
box -8 -3 16 105
use FILL  FILL_4429
timestamp 1712622712
transform 1 0 320 0 1 570
box -8 -3 16 105
use FILL  FILL_4430
timestamp 1712622712
transform 1 0 312 0 1 570
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1712622712
transform 1 0 280 0 1 570
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1712622712
transform 1 0 272 0 1 570
box -8 -3 16 105
use FILL  FILL_4433
timestamp 1712622712
transform 1 0 264 0 1 570
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1712622712
transform 1 0 256 0 1 570
box -8 -3 16 105
use FILL  FILL_4435
timestamp 1712622712
transform 1 0 248 0 1 570
box -8 -3 16 105
use FILL  FILL_4436
timestamp 1712622712
transform 1 0 240 0 1 570
box -8 -3 16 105
use FILL  FILL_4437
timestamp 1712622712
transform 1 0 192 0 1 570
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1712622712
transform 1 0 184 0 1 570
box -8 -3 16 105
use FILL  FILL_4439
timestamp 1712622712
transform 1 0 176 0 1 570
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1712622712
transform 1 0 168 0 1 570
box -8 -3 16 105
use FILL  FILL_4441
timestamp 1712622712
transform 1 0 160 0 1 570
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1712622712
transform 1 0 128 0 1 570
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1712622712
transform 1 0 120 0 1 570
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1712622712
transform 1 0 88 0 1 570
box -8 -3 16 105
use FILL  FILL_4445
timestamp 1712622712
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_4446
timestamp 1712622712
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1712622712
transform 1 0 3424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1712622712
transform 1 0 3384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4449
timestamp 1712622712
transform 1 0 3376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4450
timestamp 1712622712
transform 1 0 3368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1712622712
transform 1 0 3328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1712622712
transform 1 0 3288 0 -1 570
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1712622712
transform 1 0 3280 0 -1 570
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1712622712
transform 1 0 3272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4455
timestamp 1712622712
transform 1 0 3264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1712622712
transform 1 0 3224 0 -1 570
box -8 -3 16 105
use FILL  FILL_4457
timestamp 1712622712
transform 1 0 3216 0 -1 570
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1712622712
transform 1 0 3176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4459
timestamp 1712622712
transform 1 0 3168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1712622712
transform 1 0 3160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1712622712
transform 1 0 3152 0 -1 570
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1712622712
transform 1 0 3104 0 -1 570
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1712622712
transform 1 0 3096 0 -1 570
box -8 -3 16 105
use FILL  FILL_4464
timestamp 1712622712
transform 1 0 3056 0 -1 570
box -8 -3 16 105
use FILL  FILL_4465
timestamp 1712622712
transform 1 0 3048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1712622712
transform 1 0 3040 0 -1 570
box -8 -3 16 105
use FILL  FILL_4467
timestamp 1712622712
transform 1 0 3032 0 -1 570
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1712622712
transform 1 0 2984 0 -1 570
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1712622712
transform 1 0 2976 0 -1 570
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1712622712
transform 1 0 2936 0 -1 570
box -8 -3 16 105
use FILL  FILL_4471
timestamp 1712622712
transform 1 0 2928 0 -1 570
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1712622712
transform 1 0 2920 0 -1 570
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1712622712
transform 1 0 2896 0 -1 570
box -8 -3 16 105
use FILL  FILL_4474
timestamp 1712622712
transform 1 0 2856 0 -1 570
box -8 -3 16 105
use FILL  FILL_4475
timestamp 1712622712
transform 1 0 2848 0 -1 570
box -8 -3 16 105
use FILL  FILL_4476
timestamp 1712622712
transform 1 0 2824 0 -1 570
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1712622712
transform 1 0 2816 0 -1 570
box -8 -3 16 105
use FILL  FILL_4478
timestamp 1712622712
transform 1 0 2768 0 -1 570
box -8 -3 16 105
use FILL  FILL_4479
timestamp 1712622712
transform 1 0 2760 0 -1 570
box -8 -3 16 105
use FILL  FILL_4480
timestamp 1712622712
transform 1 0 2752 0 -1 570
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1712622712
transform 1 0 2744 0 -1 570
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1712622712
transform 1 0 2696 0 -1 570
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1712622712
transform 1 0 2688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1712622712
transform 1 0 2680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1712622712
transform 1 0 2640 0 -1 570
box -8 -3 16 105
use FILL  FILL_4486
timestamp 1712622712
transform 1 0 2632 0 -1 570
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1712622712
transform 1 0 2624 0 -1 570
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1712622712
transform 1 0 2616 0 -1 570
box -8 -3 16 105
use FILL  FILL_4489
timestamp 1712622712
transform 1 0 2568 0 -1 570
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1712622712
transform 1 0 2560 0 -1 570
box -8 -3 16 105
use FILL  FILL_4491
timestamp 1712622712
transform 1 0 2552 0 -1 570
box -8 -3 16 105
use FILL  FILL_4492
timestamp 1712622712
transform 1 0 2544 0 -1 570
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1712622712
transform 1 0 2536 0 -1 570
box -8 -3 16 105
use FILL  FILL_4494
timestamp 1712622712
transform 1 0 2480 0 -1 570
box -8 -3 16 105
use FILL  FILL_4495
timestamp 1712622712
transform 1 0 2472 0 -1 570
box -8 -3 16 105
use FILL  FILL_4496
timestamp 1712622712
transform 1 0 2464 0 -1 570
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1712622712
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4498
timestamp 1712622712
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1712622712
transform 1 0 2392 0 -1 570
box -8 -3 16 105
use FILL  FILL_4500
timestamp 1712622712
transform 1 0 2384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4501
timestamp 1712622712
transform 1 0 2376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1712622712
transform 1 0 2328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4503
timestamp 1712622712
transform 1 0 2320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1712622712
transform 1 0 2312 0 -1 570
box -8 -3 16 105
use FILL  FILL_4505
timestamp 1712622712
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1712622712
transform 1 0 2256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1712622712
transform 1 0 2248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1712622712
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1712622712
transform 1 0 2232 0 -1 570
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1712622712
transform 1 0 2184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1712622712
transform 1 0 2176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4512
timestamp 1712622712
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1712622712
transform 1 0 2128 0 -1 570
box -8 -3 16 105
use FILL  FILL_4514
timestamp 1712622712
transform 1 0 2120 0 -1 570
box -8 -3 16 105
use FILL  FILL_4515
timestamp 1712622712
transform 1 0 2112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1712622712
transform 1 0 2104 0 -1 570
box -8 -3 16 105
use FILL  FILL_4517
timestamp 1712622712
transform 1 0 2056 0 -1 570
box -8 -3 16 105
use FILL  FILL_4518
timestamp 1712622712
transform 1 0 2048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4519
timestamp 1712622712
transform 1 0 2024 0 -1 570
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1712622712
transform 1 0 2016 0 -1 570
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1712622712
transform 1 0 1968 0 -1 570
box -8 -3 16 105
use FILL  FILL_4522
timestamp 1712622712
transform 1 0 1960 0 -1 570
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1712622712
transform 1 0 1952 0 -1 570
box -8 -3 16 105
use FILL  FILL_4524
timestamp 1712622712
transform 1 0 1904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1712622712
transform 1 0 1896 0 -1 570
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1712622712
transform 1 0 1888 0 -1 570
box -8 -3 16 105
use FILL  FILL_4527
timestamp 1712622712
transform 1 0 1880 0 -1 570
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1712622712
transform 1 0 1840 0 -1 570
box -8 -3 16 105
use FILL  FILL_4529
timestamp 1712622712
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1712622712
transform 1 0 1784 0 -1 570
box -8 -3 16 105
use FILL  FILL_4531
timestamp 1712622712
transform 1 0 1776 0 -1 570
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1712622712
transform 1 0 1768 0 -1 570
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1712622712
transform 1 0 1728 0 -1 570
box -8 -3 16 105
use FILL  FILL_4534
timestamp 1712622712
transform 1 0 1688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1712622712
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4536
timestamp 1712622712
transform 1 0 1672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4537
timestamp 1712622712
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use FILL  FILL_4538
timestamp 1712622712
transform 1 0 1608 0 -1 570
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1712622712
transform 1 0 1600 0 -1 570
box -8 -3 16 105
use FILL  FILL_4540
timestamp 1712622712
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1712622712
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4542
timestamp 1712622712
transform 1 0 1520 0 -1 570
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1712622712
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1712622712
transform 1 0 1504 0 -1 570
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1712622712
transform 1 0 1496 0 -1 570
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1712622712
transform 1 0 1448 0 -1 570
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1712622712
transform 1 0 1440 0 -1 570
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1712622712
transform 1 0 1432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4549
timestamp 1712622712
transform 1 0 1384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1712622712
transform 1 0 1376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4551
timestamp 1712622712
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4552
timestamp 1712622712
transform 1 0 1336 0 -1 570
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1712622712
transform 1 0 1328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1712622712
transform 1 0 1320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4555
timestamp 1712622712
transform 1 0 1272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4556
timestamp 1712622712
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1712622712
transform 1 0 1256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1712622712
transform 1 0 1248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4559
timestamp 1712622712
transform 1 0 1192 0 -1 570
box -8 -3 16 105
use FILL  FILL_4560
timestamp 1712622712
transform 1 0 1184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4561
timestamp 1712622712
transform 1 0 1176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4562
timestamp 1712622712
transform 1 0 1168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1712622712
transform 1 0 1120 0 -1 570
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1712622712
transform 1 0 1112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1712622712
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1712622712
transform 1 0 1072 0 -1 570
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1712622712
transform 1 0 1064 0 -1 570
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1712622712
transform 1 0 1016 0 -1 570
box -8 -3 16 105
use FILL  FILL_4569
timestamp 1712622712
transform 1 0 1008 0 -1 570
box -8 -3 16 105
use FILL  FILL_4570
timestamp 1712622712
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1712622712
transform 1 0 952 0 -1 570
box -8 -3 16 105
use FILL  FILL_4572
timestamp 1712622712
transform 1 0 944 0 -1 570
box -8 -3 16 105
use FILL  FILL_4573
timestamp 1712622712
transform 1 0 936 0 -1 570
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1712622712
transform 1 0 928 0 -1 570
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1712622712
transform 1 0 904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4576
timestamp 1712622712
transform 1 0 840 0 -1 570
box -8 -3 16 105
use FILL  FILL_4577
timestamp 1712622712
transform 1 0 832 0 -1 570
box -8 -3 16 105
use FILL  FILL_4578
timestamp 1712622712
transform 1 0 824 0 -1 570
box -8 -3 16 105
use FILL  FILL_4579
timestamp 1712622712
transform 1 0 816 0 -1 570
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1712622712
transform 1 0 768 0 -1 570
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1712622712
transform 1 0 760 0 -1 570
box -8 -3 16 105
use FILL  FILL_4582
timestamp 1712622712
transform 1 0 720 0 -1 570
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1712622712
transform 1 0 712 0 -1 570
box -8 -3 16 105
use FILL  FILL_4584
timestamp 1712622712
transform 1 0 704 0 -1 570
box -8 -3 16 105
use FILL  FILL_4585
timestamp 1712622712
transform 1 0 656 0 -1 570
box -8 -3 16 105
use FILL  FILL_4586
timestamp 1712622712
transform 1 0 648 0 -1 570
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1712622712
transform 1 0 640 0 -1 570
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1712622712
transform 1 0 584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1712622712
transform 1 0 576 0 -1 570
box -8 -3 16 105
use FILL  FILL_4590
timestamp 1712622712
transform 1 0 568 0 -1 570
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1712622712
transform 1 0 560 0 -1 570
box -8 -3 16 105
use FILL  FILL_4592
timestamp 1712622712
transform 1 0 512 0 -1 570
box -8 -3 16 105
use FILL  FILL_4593
timestamp 1712622712
transform 1 0 488 0 -1 570
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1712622712
transform 1 0 480 0 -1 570
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1712622712
transform 1 0 472 0 -1 570
box -8 -3 16 105
use FILL  FILL_4596
timestamp 1712622712
transform 1 0 464 0 -1 570
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1712622712
transform 1 0 408 0 -1 570
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1712622712
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_4599
timestamp 1712622712
transform 1 0 392 0 -1 570
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1712622712
transform 1 0 384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4601
timestamp 1712622712
transform 1 0 344 0 -1 570
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1712622712
transform 1 0 304 0 -1 570
box -8 -3 16 105
use FILL  FILL_4603
timestamp 1712622712
transform 1 0 296 0 -1 570
box -8 -3 16 105
use FILL  FILL_4604
timestamp 1712622712
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_4605
timestamp 1712622712
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1712622712
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1712622712
transform 1 0 232 0 -1 570
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1712622712
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1712622712
transform 1 0 176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1712622712
transform 1 0 168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1712622712
transform 1 0 160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4612
timestamp 1712622712
transform 1 0 88 0 -1 570
box -8 -3 16 105
use FILL  FILL_4613
timestamp 1712622712
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1712622712
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1712622712
transform 1 0 3424 0 1 370
box -8 -3 16 105
use FILL  FILL_4616
timestamp 1712622712
transform 1 0 3320 0 1 370
box -8 -3 16 105
use FILL  FILL_4617
timestamp 1712622712
transform 1 0 3216 0 1 370
box -8 -3 16 105
use FILL  FILL_4618
timestamp 1712622712
transform 1 0 3208 0 1 370
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1712622712
transform 1 0 3200 0 1 370
box -8 -3 16 105
use FILL  FILL_4620
timestamp 1712622712
transform 1 0 3096 0 1 370
box -8 -3 16 105
use FILL  FILL_4621
timestamp 1712622712
transform 1 0 3056 0 1 370
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1712622712
transform 1 0 3048 0 1 370
box -8 -3 16 105
use FILL  FILL_4623
timestamp 1712622712
transform 1 0 3040 0 1 370
box -8 -3 16 105
use FILL  FILL_4624
timestamp 1712622712
transform 1 0 2936 0 1 370
box -8 -3 16 105
use FILL  FILL_4625
timestamp 1712622712
transform 1 0 2928 0 1 370
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1712622712
transform 1 0 2920 0 1 370
box -8 -3 16 105
use FILL  FILL_4627
timestamp 1712622712
transform 1 0 2848 0 1 370
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1712622712
transform 1 0 2840 0 1 370
box -8 -3 16 105
use FILL  FILL_4629
timestamp 1712622712
transform 1 0 2832 0 1 370
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1712622712
transform 1 0 2728 0 1 370
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1712622712
transform 1 0 2720 0 1 370
box -8 -3 16 105
use FILL  FILL_4632
timestamp 1712622712
transform 1 0 2712 0 1 370
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1712622712
transform 1 0 2704 0 1 370
box -8 -3 16 105
use FILL  FILL_4634
timestamp 1712622712
transform 1 0 2696 0 1 370
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1712622712
transform 1 0 2648 0 1 370
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1712622712
transform 1 0 2640 0 1 370
box -8 -3 16 105
use FILL  FILL_4637
timestamp 1712622712
transform 1 0 2632 0 1 370
box -8 -3 16 105
use FILL  FILL_4638
timestamp 1712622712
transform 1 0 2592 0 1 370
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1712622712
transform 1 0 2584 0 1 370
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1712622712
transform 1 0 2576 0 1 370
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1712622712
transform 1 0 2552 0 1 370
box -8 -3 16 105
use FILL  FILL_4642
timestamp 1712622712
transform 1 0 2544 0 1 370
box -8 -3 16 105
use FILL  FILL_4643
timestamp 1712622712
transform 1 0 2536 0 1 370
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1712622712
transform 1 0 2528 0 1 370
box -8 -3 16 105
use FILL  FILL_4645
timestamp 1712622712
transform 1 0 2488 0 1 370
box -8 -3 16 105
use FILL  FILL_4646
timestamp 1712622712
transform 1 0 2480 0 1 370
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1712622712
transform 1 0 2472 0 1 370
box -8 -3 16 105
use FILL  FILL_4648
timestamp 1712622712
transform 1 0 2464 0 1 370
box -8 -3 16 105
use FILL  FILL_4649
timestamp 1712622712
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1712622712
transform 1 0 2424 0 1 370
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1712622712
transform 1 0 2400 0 1 370
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1712622712
transform 1 0 2392 0 1 370
box -8 -3 16 105
use FILL  FILL_4653
timestamp 1712622712
transform 1 0 2360 0 1 370
box -8 -3 16 105
use FILL  FILL_4654
timestamp 1712622712
transform 1 0 2352 0 1 370
box -8 -3 16 105
use FILL  FILL_4655
timestamp 1712622712
transform 1 0 2344 0 1 370
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1712622712
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_4657
timestamp 1712622712
transform 1 0 2328 0 1 370
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1712622712
transform 1 0 2264 0 1 370
box -8 -3 16 105
use FILL  FILL_4659
timestamp 1712622712
transform 1 0 2256 0 1 370
box -8 -3 16 105
use FILL  FILL_4660
timestamp 1712622712
transform 1 0 2248 0 1 370
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1712622712
transform 1 0 2240 0 1 370
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1712622712
transform 1 0 2232 0 1 370
box -8 -3 16 105
use FILL  FILL_4663
timestamp 1712622712
transform 1 0 2184 0 1 370
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1712622712
transform 1 0 2176 0 1 370
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1712622712
transform 1 0 2168 0 1 370
box -8 -3 16 105
use FILL  FILL_4666
timestamp 1712622712
transform 1 0 2160 0 1 370
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1712622712
transform 1 0 2152 0 1 370
box -8 -3 16 105
use FILL  FILL_4668
timestamp 1712622712
transform 1 0 2104 0 1 370
box -8 -3 16 105
use FILL  FILL_4669
timestamp 1712622712
transform 1 0 2096 0 1 370
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1712622712
transform 1 0 2088 0 1 370
box -8 -3 16 105
use FILL  FILL_4671
timestamp 1712622712
transform 1 0 2080 0 1 370
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1712622712
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1712622712
transform 1 0 2024 0 1 370
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1712622712
transform 1 0 2016 0 1 370
box -8 -3 16 105
use FILL  FILL_4675
timestamp 1712622712
transform 1 0 2008 0 1 370
box -8 -3 16 105
use FILL  FILL_4676
timestamp 1712622712
transform 1 0 1976 0 1 370
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1712622712
transform 1 0 1968 0 1 370
box -8 -3 16 105
use FILL  FILL_4678
timestamp 1712622712
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1712622712
transform 1 0 1920 0 1 370
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1712622712
transform 1 0 1912 0 1 370
box -8 -3 16 105
use FILL  FILL_4681
timestamp 1712622712
transform 1 0 1904 0 1 370
box -8 -3 16 105
use FILL  FILL_4682
timestamp 1712622712
transform 1 0 1896 0 1 370
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1712622712
transform 1 0 1848 0 1 370
box -8 -3 16 105
use FILL  FILL_4684
timestamp 1712622712
transform 1 0 1840 0 1 370
box -8 -3 16 105
use FILL  FILL_4685
timestamp 1712622712
transform 1 0 1832 0 1 370
box -8 -3 16 105
use FILL  FILL_4686
timestamp 1712622712
transform 1 0 1824 0 1 370
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1712622712
transform 1 0 1784 0 1 370
box -8 -3 16 105
use FILL  FILL_4688
timestamp 1712622712
transform 1 0 1776 0 1 370
box -8 -3 16 105
use FILL  FILL_4689
timestamp 1712622712
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_4690
timestamp 1712622712
transform 1 0 1728 0 1 370
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1712622712
transform 1 0 1720 0 1 370
box -8 -3 16 105
use FILL  FILL_4692
timestamp 1712622712
transform 1 0 1712 0 1 370
box -8 -3 16 105
use FILL  FILL_4693
timestamp 1712622712
transform 1 0 1704 0 1 370
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1712622712
transform 1 0 1696 0 1 370
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1712622712
transform 1 0 1648 0 1 370
box -8 -3 16 105
use FILL  FILL_4696
timestamp 1712622712
transform 1 0 1640 0 1 370
box -8 -3 16 105
use FILL  FILL_4697
timestamp 1712622712
transform 1 0 1632 0 1 370
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1712622712
transform 1 0 1624 0 1 370
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1712622712
transform 1 0 1584 0 1 370
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1712622712
transform 1 0 1544 0 1 370
box -8 -3 16 105
use FILL  FILL_4701
timestamp 1712622712
transform 1 0 1536 0 1 370
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1712622712
transform 1 0 1528 0 1 370
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1712622712
transform 1 0 1520 0 1 370
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1712622712
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1712622712
transform 1 0 1448 0 1 370
box -8 -3 16 105
use FILL  FILL_4706
timestamp 1712622712
transform 1 0 1440 0 1 370
box -8 -3 16 105
use FILL  FILL_4707
timestamp 1712622712
transform 1 0 1432 0 1 370
box -8 -3 16 105
use FILL  FILL_4708
timestamp 1712622712
transform 1 0 1424 0 1 370
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1712622712
transform 1 0 1384 0 1 370
box -8 -3 16 105
use FILL  FILL_4710
timestamp 1712622712
transform 1 0 1336 0 1 370
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1712622712
transform 1 0 1328 0 1 370
box -8 -3 16 105
use FILL  FILL_4712
timestamp 1712622712
transform 1 0 1320 0 1 370
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1712622712
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1712622712
transform 1 0 1304 0 1 370
box -8 -3 16 105
use FILL  FILL_4715
timestamp 1712622712
transform 1 0 1240 0 1 370
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1712622712
transform 1 0 1216 0 1 370
box -8 -3 16 105
use FILL  FILL_4717
timestamp 1712622712
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1712622712
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_4719
timestamp 1712622712
transform 1 0 1192 0 1 370
box -8 -3 16 105
use FILL  FILL_4720
timestamp 1712622712
transform 1 0 1184 0 1 370
box -8 -3 16 105
use FILL  FILL_4721
timestamp 1712622712
transform 1 0 1120 0 1 370
box -8 -3 16 105
use FILL  FILL_4722
timestamp 1712622712
transform 1 0 1112 0 1 370
box -8 -3 16 105
use FILL  FILL_4723
timestamp 1712622712
transform 1 0 1104 0 1 370
box -8 -3 16 105
use FILL  FILL_4724
timestamp 1712622712
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1712622712
transform 1 0 1088 0 1 370
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1712622712
transform 1 0 1080 0 1 370
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1712622712
transform 1 0 1024 0 1 370
box -8 -3 16 105
use FILL  FILL_4728
timestamp 1712622712
transform 1 0 1016 0 1 370
box -8 -3 16 105
use FILL  FILL_4729
timestamp 1712622712
transform 1 0 1008 0 1 370
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1712622712
transform 1 0 1000 0 1 370
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1712622712
transform 1 0 952 0 1 370
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1712622712
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_4733
timestamp 1712622712
transform 1 0 936 0 1 370
box -8 -3 16 105
use FILL  FILL_4734
timestamp 1712622712
transform 1 0 904 0 1 370
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1712622712
transform 1 0 896 0 1 370
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1712622712
transform 1 0 888 0 1 370
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1712622712
transform 1 0 856 0 1 370
box -8 -3 16 105
use FILL  FILL_4738
timestamp 1712622712
transform 1 0 848 0 1 370
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1712622712
transform 1 0 808 0 1 370
box -8 -3 16 105
use FILL  FILL_4740
timestamp 1712622712
transform 1 0 800 0 1 370
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1712622712
transform 1 0 792 0 1 370
box -8 -3 16 105
use FILL  FILL_4742
timestamp 1712622712
transform 1 0 784 0 1 370
box -8 -3 16 105
use FILL  FILL_4743
timestamp 1712622712
transform 1 0 776 0 1 370
box -8 -3 16 105
use FILL  FILL_4744
timestamp 1712622712
transform 1 0 728 0 1 370
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1712622712
transform 1 0 720 0 1 370
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1712622712
transform 1 0 712 0 1 370
box -8 -3 16 105
use FILL  FILL_4747
timestamp 1712622712
transform 1 0 704 0 1 370
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1712622712
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1712622712
transform 1 0 648 0 1 370
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1712622712
transform 1 0 640 0 1 370
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1712622712
transform 1 0 632 0 1 370
box -8 -3 16 105
use FILL  FILL_4752
timestamp 1712622712
transform 1 0 624 0 1 370
box -8 -3 16 105
use FILL  FILL_4753
timestamp 1712622712
transform 1 0 600 0 1 370
box -8 -3 16 105
use FILL  FILL_4754
timestamp 1712622712
transform 1 0 576 0 1 370
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1712622712
transform 1 0 568 0 1 370
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1712622712
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_4757
timestamp 1712622712
transform 1 0 528 0 1 370
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1712622712
transform 1 0 520 0 1 370
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1712622712
transform 1 0 512 0 1 370
box -8 -3 16 105
use FILL  FILL_4760
timestamp 1712622712
transform 1 0 504 0 1 370
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1712622712
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_4762
timestamp 1712622712
transform 1 0 448 0 1 370
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1712622712
transform 1 0 440 0 1 370
box -8 -3 16 105
use FILL  FILL_4764
timestamp 1712622712
transform 1 0 432 0 1 370
box -8 -3 16 105
use FILL  FILL_4765
timestamp 1712622712
transform 1 0 392 0 1 370
box -8 -3 16 105
use FILL  FILL_4766
timestamp 1712622712
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_4767
timestamp 1712622712
transform 1 0 376 0 1 370
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1712622712
transform 1 0 368 0 1 370
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1712622712
transform 1 0 336 0 1 370
box -8 -3 16 105
use FILL  FILL_4770
timestamp 1712622712
transform 1 0 328 0 1 370
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1712622712
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1712622712
transform 1 0 288 0 1 370
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1712622712
transform 1 0 280 0 1 370
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1712622712
transform 1 0 272 0 1 370
box -8 -3 16 105
use FILL  FILL_4775
timestamp 1712622712
transform 1 0 264 0 1 370
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1712622712
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_4777
timestamp 1712622712
transform 1 0 208 0 1 370
box -8 -3 16 105
use FILL  FILL_4778
timestamp 1712622712
transform 1 0 200 0 1 370
box -8 -3 16 105
use FILL  FILL_4779
timestamp 1712622712
transform 1 0 192 0 1 370
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1712622712
transform 1 0 184 0 1 370
box -8 -3 16 105
use FILL  FILL_4781
timestamp 1712622712
transform 1 0 152 0 1 370
box -8 -3 16 105
use FILL  FILL_4782
timestamp 1712622712
transform 1 0 144 0 1 370
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1712622712
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_4784
timestamp 1712622712
transform 1 0 88 0 1 370
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1712622712
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_4786
timestamp 1712622712
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1712622712
transform 1 0 3424 0 -1 370
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1712622712
transform 1 0 3320 0 -1 370
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1712622712
transform 1 0 3312 0 -1 370
box -8 -3 16 105
use FILL  FILL_4790
timestamp 1712622712
transform 1 0 3304 0 -1 370
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1712622712
transform 1 0 3296 0 -1 370
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1712622712
transform 1 0 3288 0 -1 370
box -8 -3 16 105
use FILL  FILL_4793
timestamp 1712622712
transform 1 0 3280 0 -1 370
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1712622712
transform 1 0 3176 0 -1 370
box -8 -3 16 105
use FILL  FILL_4795
timestamp 1712622712
transform 1 0 3168 0 -1 370
box -8 -3 16 105
use FILL  FILL_4796
timestamp 1712622712
transform 1 0 3160 0 -1 370
box -8 -3 16 105
use FILL  FILL_4797
timestamp 1712622712
transform 1 0 3152 0 -1 370
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1712622712
transform 1 0 3144 0 -1 370
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1712622712
transform 1 0 3136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1712622712
transform 1 0 3032 0 -1 370
box -8 -3 16 105
use FILL  FILL_4801
timestamp 1712622712
transform 1 0 3024 0 -1 370
box -8 -3 16 105
use FILL  FILL_4802
timestamp 1712622712
transform 1 0 3016 0 -1 370
box -8 -3 16 105
use FILL  FILL_4803
timestamp 1712622712
transform 1 0 2912 0 -1 370
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1712622712
transform 1 0 2904 0 -1 370
box -8 -3 16 105
use FILL  FILL_4805
timestamp 1712622712
transform 1 0 2896 0 -1 370
box -8 -3 16 105
use FILL  FILL_4806
timestamp 1712622712
transform 1 0 2792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4807
timestamp 1712622712
transform 1 0 2784 0 -1 370
box -8 -3 16 105
use FILL  FILL_4808
timestamp 1712622712
transform 1 0 2776 0 -1 370
box -8 -3 16 105
use FILL  FILL_4809
timestamp 1712622712
transform 1 0 2768 0 -1 370
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1712622712
transform 1 0 2760 0 -1 370
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1712622712
transform 1 0 2704 0 -1 370
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1712622712
transform 1 0 2696 0 -1 370
box -8 -3 16 105
use FILL  FILL_4813
timestamp 1712622712
transform 1 0 2688 0 -1 370
box -8 -3 16 105
use FILL  FILL_4814
timestamp 1712622712
transform 1 0 2680 0 -1 370
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1712622712
transform 1 0 2672 0 -1 370
box -8 -3 16 105
use FILL  FILL_4816
timestamp 1712622712
transform 1 0 2632 0 -1 370
box -8 -3 16 105
use FILL  FILL_4817
timestamp 1712622712
transform 1 0 2624 0 -1 370
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1712622712
transform 1 0 2616 0 -1 370
box -8 -3 16 105
use FILL  FILL_4819
timestamp 1712622712
transform 1 0 2608 0 -1 370
box -8 -3 16 105
use FILL  FILL_4820
timestamp 1712622712
transform 1 0 2568 0 -1 370
box -8 -3 16 105
use FILL  FILL_4821
timestamp 1712622712
transform 1 0 2560 0 -1 370
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1712622712
transform 1 0 2536 0 -1 370
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1712622712
transform 1 0 2528 0 -1 370
box -8 -3 16 105
use FILL  FILL_4824
timestamp 1712622712
transform 1 0 2520 0 -1 370
box -8 -3 16 105
use FILL  FILL_4825
timestamp 1712622712
transform 1 0 2512 0 -1 370
box -8 -3 16 105
use FILL  FILL_4826
timestamp 1712622712
transform 1 0 2504 0 -1 370
box -8 -3 16 105
use FILL  FILL_4827
timestamp 1712622712
transform 1 0 2448 0 -1 370
box -8 -3 16 105
use FILL  FILL_4828
timestamp 1712622712
transform 1 0 2440 0 -1 370
box -8 -3 16 105
use FILL  FILL_4829
timestamp 1712622712
transform 1 0 2432 0 -1 370
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1712622712
transform 1 0 2424 0 -1 370
box -8 -3 16 105
use FILL  FILL_4831
timestamp 1712622712
transform 1 0 2416 0 -1 370
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1712622712
transform 1 0 2368 0 -1 370
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1712622712
transform 1 0 2360 0 -1 370
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1712622712
transform 1 0 2352 0 -1 370
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1712622712
transform 1 0 2344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4836
timestamp 1712622712
transform 1 0 2312 0 -1 370
box -8 -3 16 105
use FILL  FILL_4837
timestamp 1712622712
transform 1 0 2304 0 -1 370
box -8 -3 16 105
use FILL  FILL_4838
timestamp 1712622712
transform 1 0 2296 0 -1 370
box -8 -3 16 105
use FILL  FILL_4839
timestamp 1712622712
transform 1 0 2288 0 -1 370
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1712622712
transform 1 0 2256 0 -1 370
box -8 -3 16 105
use FILL  FILL_4841
timestamp 1712622712
transform 1 0 2216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1712622712
transform 1 0 2208 0 -1 370
box -8 -3 16 105
use FILL  FILL_4843
timestamp 1712622712
transform 1 0 2200 0 -1 370
box -8 -3 16 105
use FILL  FILL_4844
timestamp 1712622712
transform 1 0 2192 0 -1 370
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1712622712
transform 1 0 2184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4846
timestamp 1712622712
transform 1 0 2176 0 -1 370
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1712622712
transform 1 0 2128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1712622712
transform 1 0 2120 0 -1 370
box -8 -3 16 105
use FILL  FILL_4849
timestamp 1712622712
transform 1 0 2112 0 -1 370
box -8 -3 16 105
use FILL  FILL_4850
timestamp 1712622712
transform 1 0 2104 0 -1 370
box -8 -3 16 105
use FILL  FILL_4851
timestamp 1712622712
transform 1 0 2064 0 -1 370
box -8 -3 16 105
use FILL  FILL_4852
timestamp 1712622712
transform 1 0 2056 0 -1 370
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1712622712
transform 1 0 2048 0 -1 370
box -8 -3 16 105
use FILL  FILL_4854
timestamp 1712622712
transform 1 0 2016 0 -1 370
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1712622712
transform 1 0 2008 0 -1 370
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1712622712
transform 1 0 2000 0 -1 370
box -8 -3 16 105
use FILL  FILL_4857
timestamp 1712622712
transform 1 0 1992 0 -1 370
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1712622712
transform 1 0 1984 0 -1 370
box -8 -3 16 105
use FILL  FILL_4859
timestamp 1712622712
transform 1 0 1936 0 -1 370
box -8 -3 16 105
use FILL  FILL_4860
timestamp 1712622712
transform 1 0 1928 0 -1 370
box -8 -3 16 105
use FILL  FILL_4861
timestamp 1712622712
transform 1 0 1920 0 -1 370
box -8 -3 16 105
use FILL  FILL_4862
timestamp 1712622712
transform 1 0 1912 0 -1 370
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1712622712
transform 1 0 1904 0 -1 370
box -8 -3 16 105
use FILL  FILL_4864
timestamp 1712622712
transform 1 0 1864 0 -1 370
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1712622712
transform 1 0 1856 0 -1 370
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1712622712
transform 1 0 1848 0 -1 370
box -8 -3 16 105
use FILL  FILL_4867
timestamp 1712622712
transform 1 0 1816 0 -1 370
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1712622712
transform 1 0 1808 0 -1 370
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1712622712
transform 1 0 1800 0 -1 370
box -8 -3 16 105
use FILL  FILL_4870
timestamp 1712622712
transform 1 0 1792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4871
timestamp 1712622712
transform 1 0 1760 0 -1 370
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1712622712
transform 1 0 1752 0 -1 370
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1712622712
transform 1 0 1704 0 -1 370
box -8 -3 16 105
use FILL  FILL_4874
timestamp 1712622712
transform 1 0 1696 0 -1 370
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1712622712
transform 1 0 1688 0 -1 370
box -8 -3 16 105
use FILL  FILL_4876
timestamp 1712622712
transform 1 0 1680 0 -1 370
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1712622712
transform 1 0 1672 0 -1 370
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1712622712
transform 1 0 1640 0 -1 370
box -8 -3 16 105
use FILL  FILL_4879
timestamp 1712622712
transform 1 0 1632 0 -1 370
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1712622712
transform 1 0 1584 0 -1 370
box -8 -3 16 105
use FILL  FILL_4881
timestamp 1712622712
transform 1 0 1576 0 -1 370
box -8 -3 16 105
use FILL  FILL_4882
timestamp 1712622712
transform 1 0 1568 0 -1 370
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1712622712
transform 1 0 1560 0 -1 370
box -8 -3 16 105
use FILL  FILL_4884
timestamp 1712622712
transform 1 0 1552 0 -1 370
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1712622712
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_4886
timestamp 1712622712
transform 1 0 1480 0 -1 370
box -8 -3 16 105
use FILL  FILL_4887
timestamp 1712622712
transform 1 0 1472 0 -1 370
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1712622712
transform 1 0 1464 0 -1 370
box -8 -3 16 105
use FILL  FILL_4889
timestamp 1712622712
transform 1 0 1456 0 -1 370
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1712622712
transform 1 0 1448 0 -1 370
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1712622712
transform 1 0 1440 0 -1 370
box -8 -3 16 105
use FILL  FILL_4892
timestamp 1712622712
transform 1 0 1384 0 -1 370
box -8 -3 16 105
use FILL  FILL_4893
timestamp 1712622712
transform 1 0 1376 0 -1 370
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1712622712
transform 1 0 1368 0 -1 370
box -8 -3 16 105
use FILL  FILL_4895
timestamp 1712622712
transform 1 0 1360 0 -1 370
box -8 -3 16 105
use FILL  FILL_4896
timestamp 1712622712
transform 1 0 1352 0 -1 370
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1712622712
transform 1 0 1344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1712622712
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1712622712
transform 1 0 1328 0 -1 370
box -8 -3 16 105
use FILL  FILL_4900
timestamp 1712622712
transform 1 0 1264 0 -1 370
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1712622712
transform 1 0 1256 0 -1 370
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1712622712
transform 1 0 1248 0 -1 370
box -8 -3 16 105
use FILL  FILL_4903
timestamp 1712622712
transform 1 0 1240 0 -1 370
box -8 -3 16 105
use FILL  FILL_4904
timestamp 1712622712
transform 1 0 1232 0 -1 370
box -8 -3 16 105
use FILL  FILL_4905
timestamp 1712622712
transform 1 0 1208 0 -1 370
box -8 -3 16 105
use FILL  FILL_4906
timestamp 1712622712
transform 1 0 1200 0 -1 370
box -8 -3 16 105
use FILL  FILL_4907
timestamp 1712622712
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1712622712
transform 1 0 1144 0 -1 370
box -8 -3 16 105
use FILL  FILL_4909
timestamp 1712622712
transform 1 0 1136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4910
timestamp 1712622712
transform 1 0 1128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1712622712
transform 1 0 1120 0 -1 370
box -8 -3 16 105
use FILL  FILL_4912
timestamp 1712622712
transform 1 0 1080 0 -1 370
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1712622712
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_4914
timestamp 1712622712
transform 1 0 1064 0 -1 370
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1712622712
transform 1 0 1032 0 -1 370
box -8 -3 16 105
use FILL  FILL_4916
timestamp 1712622712
transform 1 0 1024 0 -1 370
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1712622712
transform 1 0 1016 0 -1 370
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1712622712
transform 1 0 1008 0 -1 370
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1712622712
transform 1 0 976 0 -1 370
box -8 -3 16 105
use FILL  FILL_4920
timestamp 1712622712
transform 1 0 968 0 -1 370
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1712622712
transform 1 0 960 0 -1 370
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1712622712
transform 1 0 912 0 -1 370
box -8 -3 16 105
use FILL  FILL_4923
timestamp 1712622712
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1712622712
transform 1 0 896 0 -1 370
box -8 -3 16 105
use FILL  FILL_4925
timestamp 1712622712
transform 1 0 888 0 -1 370
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1712622712
transform 1 0 880 0 -1 370
box -8 -3 16 105
use FILL  FILL_4927
timestamp 1712622712
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_4928
timestamp 1712622712
transform 1 0 840 0 -1 370
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1712622712
transform 1 0 832 0 -1 370
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1712622712
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1712622712
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1712622712
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_4933
timestamp 1712622712
transform 1 0 744 0 -1 370
box -8 -3 16 105
use FILL  FILL_4934
timestamp 1712622712
transform 1 0 736 0 -1 370
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1712622712
transform 1 0 728 0 -1 370
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1712622712
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1712622712
transform 1 0 712 0 -1 370
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1712622712
transform 1 0 704 0 -1 370
box -8 -3 16 105
use FILL  FILL_4939
timestamp 1712622712
transform 1 0 696 0 -1 370
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1712622712
transform 1 0 632 0 -1 370
box -8 -3 16 105
use FILL  FILL_4941
timestamp 1712622712
transform 1 0 624 0 -1 370
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1712622712
transform 1 0 616 0 -1 370
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1712622712
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_4944
timestamp 1712622712
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1712622712
transform 1 0 568 0 -1 370
box -8 -3 16 105
use FILL  FILL_4946
timestamp 1712622712
transform 1 0 560 0 -1 370
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1712622712
transform 1 0 552 0 -1 370
box -8 -3 16 105
use FILL  FILL_4948
timestamp 1712622712
transform 1 0 504 0 -1 370
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1712622712
transform 1 0 496 0 -1 370
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1712622712
transform 1 0 488 0 -1 370
box -8 -3 16 105
use FILL  FILL_4951
timestamp 1712622712
transform 1 0 480 0 -1 370
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1712622712
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1712622712
transform 1 0 424 0 -1 370
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1712622712
transform 1 0 416 0 -1 370
box -8 -3 16 105
use FILL  FILL_4955
timestamp 1712622712
transform 1 0 408 0 -1 370
box -8 -3 16 105
use FILL  FILL_4956
timestamp 1712622712
transform 1 0 400 0 -1 370
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1712622712
transform 1 0 352 0 -1 370
box -8 -3 16 105
use FILL  FILL_4958
timestamp 1712622712
transform 1 0 344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4959
timestamp 1712622712
transform 1 0 336 0 -1 370
box -8 -3 16 105
use FILL  FILL_4960
timestamp 1712622712
transform 1 0 296 0 -1 370
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1712622712
transform 1 0 288 0 -1 370
box -8 -3 16 105
use FILL  FILL_4962
timestamp 1712622712
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_4963
timestamp 1712622712
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1712622712
transform 1 0 264 0 -1 370
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1712622712
transform 1 0 232 0 -1 370
box -8 -3 16 105
use FILL  FILL_4966
timestamp 1712622712
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_4967
timestamp 1712622712
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1712622712
transform 1 0 176 0 -1 370
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1712622712
transform 1 0 168 0 -1 370
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1712622712
transform 1 0 160 0 -1 370
box -8 -3 16 105
use FILL  FILL_4971
timestamp 1712622712
transform 1 0 152 0 -1 370
box -8 -3 16 105
use FILL  FILL_4972
timestamp 1712622712
transform 1 0 88 0 -1 370
box -8 -3 16 105
use FILL  FILL_4973
timestamp 1712622712
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1712622712
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_4975
timestamp 1712622712
transform 1 0 3368 0 1 170
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1712622712
transform 1 0 3360 0 1 170
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1712622712
transform 1 0 3352 0 1 170
box -8 -3 16 105
use FILL  FILL_4978
timestamp 1712622712
transform 1 0 3344 0 1 170
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1712622712
transform 1 0 3256 0 1 170
box -8 -3 16 105
use FILL  FILL_4980
timestamp 1712622712
transform 1 0 3248 0 1 170
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1712622712
transform 1 0 3240 0 1 170
box -8 -3 16 105
use FILL  FILL_4982
timestamp 1712622712
transform 1 0 3232 0 1 170
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1712622712
transform 1 0 3224 0 1 170
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1712622712
transform 1 0 3168 0 1 170
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1712622712
transform 1 0 3160 0 1 170
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1712622712
transform 1 0 3152 0 1 170
box -8 -3 16 105
use FILL  FILL_4987
timestamp 1712622712
transform 1 0 3088 0 1 170
box -8 -3 16 105
use FILL  FILL_4988
timestamp 1712622712
transform 1 0 3080 0 1 170
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1712622712
transform 1 0 3072 0 1 170
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1712622712
transform 1 0 3040 0 1 170
box -8 -3 16 105
use FILL  FILL_4991
timestamp 1712622712
transform 1 0 3032 0 1 170
box -8 -3 16 105
use FILL  FILL_4992
timestamp 1712622712
transform 1 0 2968 0 1 170
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1712622712
transform 1 0 2960 0 1 170
box -8 -3 16 105
use FILL  FILL_4994
timestamp 1712622712
transform 1 0 2952 0 1 170
box -8 -3 16 105
use FILL  FILL_4995
timestamp 1712622712
transform 1 0 2928 0 1 170
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1712622712
transform 1 0 2888 0 1 170
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1712622712
transform 1 0 2880 0 1 170
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1712622712
transform 1 0 2872 0 1 170
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1712622712
transform 1 0 2864 0 1 170
box -8 -3 16 105
use FILL  FILL_5000
timestamp 1712622712
transform 1 0 2800 0 1 170
box -8 -3 16 105
use FILL  FILL_5001
timestamp 1712622712
transform 1 0 2776 0 1 170
box -8 -3 16 105
use FILL  FILL_5002
timestamp 1712622712
transform 1 0 2768 0 1 170
box -8 -3 16 105
use FILL  FILL_5003
timestamp 1712622712
transform 1 0 2728 0 1 170
box -8 -3 16 105
use FILL  FILL_5004
timestamp 1712622712
transform 1 0 2720 0 1 170
box -8 -3 16 105
use FILL  FILL_5005
timestamp 1712622712
transform 1 0 2712 0 1 170
box -8 -3 16 105
use FILL  FILL_5006
timestamp 1712622712
transform 1 0 2704 0 1 170
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1712622712
transform 1 0 2696 0 1 170
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1712622712
transform 1 0 2688 0 1 170
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1712622712
transform 1 0 2680 0 1 170
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1712622712
transform 1 0 2624 0 1 170
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1712622712
transform 1 0 2616 0 1 170
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1712622712
transform 1 0 2608 0 1 170
box -8 -3 16 105
use FILL  FILL_5013
timestamp 1712622712
transform 1 0 2600 0 1 170
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1712622712
transform 1 0 2592 0 1 170
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1712622712
transform 1 0 2584 0 1 170
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1712622712
transform 1 0 2576 0 1 170
box -8 -3 16 105
use FILL  FILL_5017
timestamp 1712622712
transform 1 0 2520 0 1 170
box -8 -3 16 105
use FILL  FILL_5018
timestamp 1712622712
transform 1 0 2512 0 1 170
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1712622712
transform 1 0 2504 0 1 170
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1712622712
transform 1 0 2496 0 1 170
box -8 -3 16 105
use FILL  FILL_5021
timestamp 1712622712
transform 1 0 2488 0 1 170
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1712622712
transform 1 0 2480 0 1 170
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1712622712
transform 1 0 2440 0 1 170
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1712622712
transform 1 0 2432 0 1 170
box -8 -3 16 105
use FILL  FILL_5025
timestamp 1712622712
transform 1 0 2424 0 1 170
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1712622712
transform 1 0 2384 0 1 170
box -8 -3 16 105
use FILL  FILL_5027
timestamp 1712622712
transform 1 0 2376 0 1 170
box -8 -3 16 105
use FILL  FILL_5028
timestamp 1712622712
transform 1 0 2368 0 1 170
box -8 -3 16 105
use FILL  FILL_5029
timestamp 1712622712
transform 1 0 2360 0 1 170
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1712622712
transform 1 0 2352 0 1 170
box -8 -3 16 105
use FILL  FILL_5031
timestamp 1712622712
transform 1 0 2304 0 1 170
box -8 -3 16 105
use FILL  FILL_5032
timestamp 1712622712
transform 1 0 2296 0 1 170
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1712622712
transform 1 0 2288 0 1 170
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1712622712
transform 1 0 2280 0 1 170
box -8 -3 16 105
use FILL  FILL_5035
timestamp 1712622712
transform 1 0 2272 0 1 170
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1712622712
transform 1 0 2264 0 1 170
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1712622712
transform 1 0 2216 0 1 170
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1712622712
transform 1 0 2208 0 1 170
box -8 -3 16 105
use FILL  FILL_5039
timestamp 1712622712
transform 1 0 2200 0 1 170
box -8 -3 16 105
use FILL  FILL_5040
timestamp 1712622712
transform 1 0 2192 0 1 170
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1712622712
transform 1 0 2160 0 1 170
box -8 -3 16 105
use FILL  FILL_5042
timestamp 1712622712
transform 1 0 2152 0 1 170
box -8 -3 16 105
use FILL  FILL_5043
timestamp 1712622712
transform 1 0 2144 0 1 170
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1712622712
transform 1 0 2136 0 1 170
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1712622712
transform 1 0 2128 0 1 170
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1712622712
transform 1 0 2080 0 1 170
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1712622712
transform 1 0 2072 0 1 170
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1712622712
transform 1 0 2064 0 1 170
box -8 -3 16 105
use FILL  FILL_5049
timestamp 1712622712
transform 1 0 2056 0 1 170
box -8 -3 16 105
use FILL  FILL_5050
timestamp 1712622712
transform 1 0 2048 0 1 170
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1712622712
transform 1 0 2016 0 1 170
box -8 -3 16 105
use FILL  FILL_5052
timestamp 1712622712
transform 1 0 1992 0 1 170
box -8 -3 16 105
use FILL  FILL_5053
timestamp 1712622712
transform 1 0 1984 0 1 170
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1712622712
transform 1 0 1976 0 1 170
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1712622712
transform 1 0 1968 0 1 170
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1712622712
transform 1 0 1960 0 1 170
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1712622712
transform 1 0 1912 0 1 170
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1712622712
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1712622712
transform 1 0 1896 0 1 170
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1712622712
transform 1 0 1888 0 1 170
box -8 -3 16 105
use FILL  FILL_5061
timestamp 1712622712
transform 1 0 1840 0 1 170
box -8 -3 16 105
use FILL  FILL_5062
timestamp 1712622712
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_5063
timestamp 1712622712
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_5064
timestamp 1712622712
transform 1 0 1816 0 1 170
box -8 -3 16 105
use FILL  FILL_5065
timestamp 1712622712
transform 1 0 1808 0 1 170
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1712622712
transform 1 0 1784 0 1 170
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1712622712
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_5068
timestamp 1712622712
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1712622712
transform 1 0 1736 0 1 170
box -8 -3 16 105
use FILL  FILL_5070
timestamp 1712622712
transform 1 0 1704 0 1 170
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1712622712
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1712622712
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_5073
timestamp 1712622712
transform 1 0 1680 0 1 170
box -8 -3 16 105
use FILL  FILL_5074
timestamp 1712622712
transform 1 0 1632 0 1 170
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1712622712
transform 1 0 1624 0 1 170
box -8 -3 16 105
use FILL  FILL_5076
timestamp 1712622712
transform 1 0 1616 0 1 170
box -8 -3 16 105
use FILL  FILL_5077
timestamp 1712622712
transform 1 0 1608 0 1 170
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1712622712
transform 1 0 1600 0 1 170
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1712622712
transform 1 0 1592 0 1 170
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1712622712
transform 1 0 1528 0 1 170
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1712622712
transform 1 0 1520 0 1 170
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1712622712
transform 1 0 1512 0 1 170
box -8 -3 16 105
use FILL  FILL_5083
timestamp 1712622712
transform 1 0 1504 0 1 170
box -8 -3 16 105
use FILL  FILL_5084
timestamp 1712622712
transform 1 0 1496 0 1 170
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1712622712
transform 1 0 1448 0 1 170
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1712622712
transform 1 0 1440 0 1 170
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1712622712
transform 1 0 1432 0 1 170
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1712622712
transform 1 0 1392 0 1 170
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1712622712
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1712622712
transform 1 0 1376 0 1 170
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1712622712
transform 1 0 1336 0 1 170
box -8 -3 16 105
use FILL  FILL_5092
timestamp 1712622712
transform 1 0 1328 0 1 170
box -8 -3 16 105
use FILL  FILL_5093
timestamp 1712622712
transform 1 0 1320 0 1 170
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1712622712
transform 1 0 1312 0 1 170
box -8 -3 16 105
use FILL  FILL_5095
timestamp 1712622712
transform 1 0 1264 0 1 170
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1712622712
transform 1 0 1256 0 1 170
box -8 -3 16 105
use FILL  FILL_5097
timestamp 1712622712
transform 1 0 1248 0 1 170
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1712622712
transform 1 0 1240 0 1 170
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1712622712
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_5100
timestamp 1712622712
transform 1 0 1184 0 1 170
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1712622712
transform 1 0 1176 0 1 170
box -8 -3 16 105
use FILL  FILL_5102
timestamp 1712622712
transform 1 0 1168 0 1 170
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1712622712
transform 1 0 1128 0 1 170
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1712622712
transform 1 0 1120 0 1 170
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1712622712
transform 1 0 1088 0 1 170
box -8 -3 16 105
use FILL  FILL_5106
timestamp 1712622712
transform 1 0 1080 0 1 170
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1712622712
transform 1 0 1072 0 1 170
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1712622712
transform 1 0 1064 0 1 170
box -8 -3 16 105
use FILL  FILL_5109
timestamp 1712622712
transform 1 0 1016 0 1 170
box -8 -3 16 105
use FILL  FILL_5110
timestamp 1712622712
transform 1 0 1008 0 1 170
box -8 -3 16 105
use FILL  FILL_5111
timestamp 1712622712
transform 1 0 1000 0 1 170
box -8 -3 16 105
use FILL  FILL_5112
timestamp 1712622712
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1712622712
transform 1 0 952 0 1 170
box -8 -3 16 105
use FILL  FILL_5114
timestamp 1712622712
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1712622712
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1712622712
transform 1 0 928 0 1 170
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1712622712
transform 1 0 888 0 1 170
box -8 -3 16 105
use FILL  FILL_5118
timestamp 1712622712
transform 1 0 856 0 1 170
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1712622712
transform 1 0 848 0 1 170
box -8 -3 16 105
use FILL  FILL_5120
timestamp 1712622712
transform 1 0 840 0 1 170
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1712622712
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_5122
timestamp 1712622712
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_5123
timestamp 1712622712
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_5124
timestamp 1712622712
transform 1 0 768 0 1 170
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1712622712
transform 1 0 736 0 1 170
box -8 -3 16 105
use FILL  FILL_5126
timestamp 1712622712
transform 1 0 728 0 1 170
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1712622712
transform 1 0 720 0 1 170
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1712622712
transform 1 0 712 0 1 170
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1712622712
transform 1 0 664 0 1 170
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1712622712
transform 1 0 656 0 1 170
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1712622712
transform 1 0 648 0 1 170
box -8 -3 16 105
use FILL  FILL_5132
timestamp 1712622712
transform 1 0 640 0 1 170
box -8 -3 16 105
use FILL  FILL_5133
timestamp 1712622712
transform 1 0 600 0 1 170
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1712622712
transform 1 0 592 0 1 170
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1712622712
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1712622712
transform 1 0 552 0 1 170
box -8 -3 16 105
use FILL  FILL_5137
timestamp 1712622712
transform 1 0 544 0 1 170
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1712622712
transform 1 0 536 0 1 170
box -8 -3 16 105
use FILL  FILL_5139
timestamp 1712622712
transform 1 0 488 0 1 170
box -8 -3 16 105
use FILL  FILL_5140
timestamp 1712622712
transform 1 0 480 0 1 170
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1712622712
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_5142
timestamp 1712622712
transform 1 0 464 0 1 170
box -8 -3 16 105
use FILL  FILL_5143
timestamp 1712622712
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_5144
timestamp 1712622712
transform 1 0 424 0 1 170
box -8 -3 16 105
use FILL  FILL_5145
timestamp 1712622712
transform 1 0 416 0 1 170
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1712622712
transform 1 0 376 0 1 170
box -8 -3 16 105
use FILL  FILL_5147
timestamp 1712622712
transform 1 0 368 0 1 170
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1712622712
transform 1 0 360 0 1 170
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1712622712
transform 1 0 320 0 1 170
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1712622712
transform 1 0 312 0 1 170
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1712622712
transform 1 0 304 0 1 170
box -8 -3 16 105
use FILL  FILL_5152
timestamp 1712622712
transform 1 0 296 0 1 170
box -8 -3 16 105
use FILL  FILL_5153
timestamp 1712622712
transform 1 0 288 0 1 170
box -8 -3 16 105
use FILL  FILL_5154
timestamp 1712622712
transform 1 0 240 0 1 170
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1712622712
transform 1 0 232 0 1 170
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1712622712
transform 1 0 224 0 1 170
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1712622712
transform 1 0 216 0 1 170
box -8 -3 16 105
use FILL  FILL_5158
timestamp 1712622712
transform 1 0 176 0 1 170
box -8 -3 16 105
use FILL  FILL_5159
timestamp 1712622712
transform 1 0 168 0 1 170
box -8 -3 16 105
use FILL  FILL_5160
timestamp 1712622712
transform 1 0 160 0 1 170
box -8 -3 16 105
use FILL  FILL_5161
timestamp 1712622712
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_5162
timestamp 1712622712
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_5163
timestamp 1712622712
transform 1 0 96 0 1 170
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1712622712
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1712622712
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_5166
timestamp 1712622712
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1712622712
transform 1 0 3424 0 -1 170
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1712622712
transform 1 0 3400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1712622712
transform 1 0 3392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5170
timestamp 1712622712
transform 1 0 3384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1712622712
transform 1 0 3376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5172
timestamp 1712622712
transform 1 0 3312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1712622712
transform 1 0 3304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5174
timestamp 1712622712
transform 1 0 3296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5175
timestamp 1712622712
transform 1 0 3288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1712622712
transform 1 0 3280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5177
timestamp 1712622712
transform 1 0 3272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1712622712
transform 1 0 3224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1712622712
transform 1 0 3216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1712622712
transform 1 0 3208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1712622712
transform 1 0 3168 0 -1 170
box -8 -3 16 105
use FILL  FILL_5182
timestamp 1712622712
transform 1 0 3160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1712622712
transform 1 0 3152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5184
timestamp 1712622712
transform 1 0 3144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1712622712
transform 1 0 3136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1712622712
transform 1 0 3128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1712622712
transform 1 0 3064 0 -1 170
box -8 -3 16 105
use FILL  FILL_5188
timestamp 1712622712
transform 1 0 3056 0 -1 170
box -8 -3 16 105
use FILL  FILL_5189
timestamp 1712622712
transform 1 0 3048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1712622712
transform 1 0 3040 0 -1 170
box -8 -3 16 105
use FILL  FILL_5191
timestamp 1712622712
transform 1 0 3032 0 -1 170
box -8 -3 16 105
use FILL  FILL_5192
timestamp 1712622712
transform 1 0 3024 0 -1 170
box -8 -3 16 105
use FILL  FILL_5193
timestamp 1712622712
transform 1 0 2944 0 -1 170
box -8 -3 16 105
use FILL  FILL_5194
timestamp 1712622712
transform 1 0 2936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1712622712
transform 1 0 2928 0 -1 170
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1712622712
transform 1 0 2896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1712622712
transform 1 0 2856 0 -1 170
box -8 -3 16 105
use FILL  FILL_5198
timestamp 1712622712
transform 1 0 2848 0 -1 170
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1712622712
transform 1 0 2840 0 -1 170
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1712622712
transform 1 0 2776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5201
timestamp 1712622712
transform 1 0 2768 0 -1 170
box -8 -3 16 105
use FILL  FILL_5202
timestamp 1712622712
transform 1 0 2736 0 -1 170
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1712622712
transform 1 0 2728 0 -1 170
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1712622712
transform 1 0 2720 0 -1 170
box -8 -3 16 105
use FILL  FILL_5205
timestamp 1712622712
transform 1 0 2696 0 -1 170
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1712622712
transform 1 0 2688 0 -1 170
box -8 -3 16 105
use FILL  FILL_5207
timestamp 1712622712
transform 1 0 2664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1712622712
transform 1 0 2656 0 -1 170
box -8 -3 16 105
use FILL  FILL_5209
timestamp 1712622712
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5210
timestamp 1712622712
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1712622712
transform 1 0 2600 0 -1 170
box -8 -3 16 105
use FILL  FILL_5212
timestamp 1712622712
transform 1 0 2592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5213
timestamp 1712622712
transform 1 0 2584 0 -1 170
box -8 -3 16 105
use FILL  FILL_5214
timestamp 1712622712
transform 1 0 2544 0 -1 170
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1712622712
transform 1 0 2536 0 -1 170
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1712622712
transform 1 0 2528 0 -1 170
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1712622712
transform 1 0 2504 0 -1 170
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1712622712
transform 1 0 2496 0 -1 170
box -8 -3 16 105
use FILL  FILL_5219
timestamp 1712622712
transform 1 0 2488 0 -1 170
box -8 -3 16 105
use FILL  FILL_5220
timestamp 1712622712
transform 1 0 2480 0 -1 170
box -8 -3 16 105
use FILL  FILL_5221
timestamp 1712622712
transform 1 0 2432 0 -1 170
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1712622712
transform 1 0 2424 0 -1 170
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1712622712
transform 1 0 2416 0 -1 170
box -8 -3 16 105
use FILL  FILL_5224
timestamp 1712622712
transform 1 0 2408 0 -1 170
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1712622712
transform 1 0 2400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5226
timestamp 1712622712
transform 1 0 2352 0 -1 170
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1712622712
transform 1 0 2344 0 -1 170
box -8 -3 16 105
use FILL  FILL_5228
timestamp 1712622712
transform 1 0 2336 0 -1 170
box -8 -3 16 105
use FILL  FILL_5229
timestamp 1712622712
transform 1 0 2328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5230
timestamp 1712622712
transform 1 0 2320 0 -1 170
box -8 -3 16 105
use FILL  FILL_5231
timestamp 1712622712
transform 1 0 2272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1712622712
transform 1 0 2264 0 -1 170
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1712622712
transform 1 0 2256 0 -1 170
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1712622712
transform 1 0 2216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1712622712
transform 1 0 2208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5236
timestamp 1712622712
transform 1 0 2200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1712622712
transform 1 0 2192 0 -1 170
box -8 -3 16 105
use FILL  FILL_5238
timestamp 1712622712
transform 1 0 2184 0 -1 170
box -8 -3 16 105
use FILL  FILL_5239
timestamp 1712622712
transform 1 0 2144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1712622712
transform 1 0 2112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1712622712
transform 1 0 2104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5242
timestamp 1712622712
transform 1 0 2096 0 -1 170
box -8 -3 16 105
use FILL  FILL_5243
timestamp 1712622712
transform 1 0 2088 0 -1 170
box -8 -3 16 105
use FILL  FILL_5244
timestamp 1712622712
transform 1 0 2080 0 -1 170
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1712622712
transform 1 0 2032 0 -1 170
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1712622712
transform 1 0 2024 0 -1 170
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1712622712
transform 1 0 2016 0 -1 170
box -8 -3 16 105
use FILL  FILL_5248
timestamp 1712622712
transform 1 0 2008 0 -1 170
box -8 -3 16 105
use FILL  FILL_5249
timestamp 1712622712
transform 1 0 2000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1712622712
transform 1 0 1960 0 -1 170
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1712622712
transform 1 0 1952 0 -1 170
box -8 -3 16 105
use FILL  FILL_5252
timestamp 1712622712
transform 1 0 1944 0 -1 170
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1712622712
transform 1 0 1904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1712622712
transform 1 0 1896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5255
timestamp 1712622712
transform 1 0 1888 0 -1 170
box -8 -3 16 105
use FILL  FILL_5256
timestamp 1712622712
transform 1 0 1864 0 -1 170
box -8 -3 16 105
use FILL  FILL_5257
timestamp 1712622712
transform 1 0 1856 0 -1 170
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1712622712
transform 1 0 1832 0 -1 170
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1712622712
transform 1 0 1800 0 -1 170
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1712622712
transform 1 0 1792 0 -1 170
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1712622712
transform 1 0 1784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5262
timestamp 1712622712
transform 1 0 1776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5263
timestamp 1712622712
transform 1 0 1728 0 -1 170
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1712622712
transform 1 0 1720 0 -1 170
box -8 -3 16 105
use FILL  FILL_5265
timestamp 1712622712
transform 1 0 1712 0 -1 170
box -8 -3 16 105
use FILL  FILL_5266
timestamp 1712622712
transform 1 0 1704 0 -1 170
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1712622712
transform 1 0 1696 0 -1 170
box -8 -3 16 105
use FILL  FILL_5268
timestamp 1712622712
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_5269
timestamp 1712622712
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1712622712
transform 1 0 1608 0 -1 170
box -8 -3 16 105
use FILL  FILL_5271
timestamp 1712622712
transform 1 0 1600 0 -1 170
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1712622712
transform 1 0 1592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1712622712
transform 1 0 1584 0 -1 170
box -8 -3 16 105
use FILL  FILL_5274
timestamp 1712622712
transform 1 0 1560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5275
timestamp 1712622712
transform 1 0 1552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5276
timestamp 1712622712
transform 1 0 1520 0 -1 170
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1712622712
transform 1 0 1512 0 -1 170
box -8 -3 16 105
use FILL  FILL_5278
timestamp 1712622712
transform 1 0 1480 0 -1 170
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1712622712
transform 1 0 1472 0 -1 170
box -8 -3 16 105
use FILL  FILL_5280
timestamp 1712622712
transform 1 0 1464 0 -1 170
box -8 -3 16 105
use FILL  FILL_5281
timestamp 1712622712
transform 1 0 1456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1712622712
transform 1 0 1448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5283
timestamp 1712622712
transform 1 0 1400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5284
timestamp 1712622712
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5285
timestamp 1712622712
transform 1 0 1384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5286
timestamp 1712622712
transform 1 0 1376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1712622712
transform 1 0 1344 0 -1 170
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1712622712
transform 1 0 1336 0 -1 170
box -8 -3 16 105
use FILL  FILL_5289
timestamp 1712622712
transform 1 0 1328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5290
timestamp 1712622712
transform 1 0 1320 0 -1 170
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1712622712
transform 1 0 1280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5292
timestamp 1712622712
transform 1 0 1272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5293
timestamp 1712622712
transform 1 0 1264 0 -1 170
box -8 -3 16 105
use FILL  FILL_5294
timestamp 1712622712
transform 1 0 1256 0 -1 170
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1712622712
transform 1 0 1216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1712622712
transform 1 0 1208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1712622712
transform 1 0 1200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1712622712
transform 1 0 1192 0 -1 170
box -8 -3 16 105
use FILL  FILL_5299
timestamp 1712622712
transform 1 0 1152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5300
timestamp 1712622712
transform 1 0 1144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1712622712
transform 1 0 1136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5302
timestamp 1712622712
transform 1 0 1128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5303
timestamp 1712622712
transform 1 0 1120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5304
timestamp 1712622712
transform 1 0 1072 0 -1 170
box -8 -3 16 105
use FILL  FILL_5305
timestamp 1712622712
transform 1 0 1064 0 -1 170
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1712622712
transform 1 0 1056 0 -1 170
box -8 -3 16 105
use FILL  FILL_5307
timestamp 1712622712
transform 1 0 1048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1712622712
transform 1 0 1008 0 -1 170
box -8 -3 16 105
use FILL  FILL_5309
timestamp 1712622712
transform 1 0 1000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1712622712
transform 1 0 992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1712622712
transform 1 0 984 0 -1 170
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1712622712
transform 1 0 936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1712622712
transform 1 0 928 0 -1 170
box -8 -3 16 105
use FILL  FILL_5314
timestamp 1712622712
transform 1 0 920 0 -1 170
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1712622712
transform 1 0 912 0 -1 170
box -8 -3 16 105
use FILL  FILL_5316
timestamp 1712622712
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5317
timestamp 1712622712
transform 1 0 856 0 -1 170
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1712622712
transform 1 0 848 0 -1 170
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1712622712
transform 1 0 840 0 -1 170
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1712622712
transform 1 0 808 0 -1 170
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1712622712
transform 1 0 800 0 -1 170
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1712622712
transform 1 0 792 0 -1 170
box -8 -3 16 105
use FILL  FILL_5323
timestamp 1712622712
transform 1 0 784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5324
timestamp 1712622712
transform 1 0 776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1712622712
transform 1 0 728 0 -1 170
box -8 -3 16 105
use FILL  FILL_5326
timestamp 1712622712
transform 1 0 720 0 -1 170
box -8 -3 16 105
use FILL  FILL_5327
timestamp 1712622712
transform 1 0 712 0 -1 170
box -8 -3 16 105
use FILL  FILL_5328
timestamp 1712622712
transform 1 0 704 0 -1 170
box -8 -3 16 105
use FILL  FILL_5329
timestamp 1712622712
transform 1 0 696 0 -1 170
box -8 -3 16 105
use FILL  FILL_5330
timestamp 1712622712
transform 1 0 688 0 -1 170
box -8 -3 16 105
use FILL  FILL_5331
timestamp 1712622712
transform 1 0 648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5332
timestamp 1712622712
transform 1 0 624 0 -1 170
box -8 -3 16 105
use FILL  FILL_5333
timestamp 1712622712
transform 1 0 616 0 -1 170
box -8 -3 16 105
use FILL  FILL_5334
timestamp 1712622712
transform 1 0 608 0 -1 170
box -8 -3 16 105
use FILL  FILL_5335
timestamp 1712622712
transform 1 0 600 0 -1 170
box -8 -3 16 105
use FILL  FILL_5336
timestamp 1712622712
transform 1 0 592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5337
timestamp 1712622712
transform 1 0 560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5338
timestamp 1712622712
transform 1 0 552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5339
timestamp 1712622712
transform 1 0 544 0 -1 170
box -8 -3 16 105
use FILL  FILL_5340
timestamp 1712622712
transform 1 0 496 0 -1 170
box -8 -3 16 105
use FILL  FILL_5341
timestamp 1712622712
transform 1 0 488 0 -1 170
box -8 -3 16 105
use FILL  FILL_5342
timestamp 1712622712
transform 1 0 480 0 -1 170
box -8 -3 16 105
use FILL  FILL_5343
timestamp 1712622712
transform 1 0 472 0 -1 170
box -8 -3 16 105
use FILL  FILL_5344
timestamp 1712622712
transform 1 0 464 0 -1 170
box -8 -3 16 105
use FILL  FILL_5345
timestamp 1712622712
transform 1 0 456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5346
timestamp 1712622712
transform 1 0 448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5347
timestamp 1712622712
transform 1 0 400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5348
timestamp 1712622712
transform 1 0 392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5349
timestamp 1712622712
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5350
timestamp 1712622712
transform 1 0 376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5351
timestamp 1712622712
transform 1 0 368 0 -1 170
box -8 -3 16 105
use FILL  FILL_5352
timestamp 1712622712
transform 1 0 360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5353
timestamp 1712622712
transform 1 0 312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5354
timestamp 1712622712
transform 1 0 304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5355
timestamp 1712622712
transform 1 0 296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5356
timestamp 1712622712
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5357
timestamp 1712622712
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5358
timestamp 1712622712
transform 1 0 272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5359
timestamp 1712622712
transform 1 0 224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5360
timestamp 1712622712
transform 1 0 216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5361
timestamp 1712622712
transform 1 0 208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5362
timestamp 1712622712
transform 1 0 200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5363
timestamp 1712622712
transform 1 0 168 0 -1 170
box -8 -3 16 105
use FILL  FILL_5364
timestamp 1712622712
transform 1 0 160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5365
timestamp 1712622712
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5366
timestamp 1712622712
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5367
timestamp 1712622712
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5368
timestamp 1712622712
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5369
timestamp 1712622712
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5370
timestamp 1712622712
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5371
timestamp 1712622712
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5372
timestamp 1712622712
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_5373
timestamp 1712622712
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_5374
timestamp 1712622712
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_5375
timestamp 1712622712
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1712622712
transform 1 0 2864 0 1 770
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1712622712
transform 1 0 3080 0 1 770
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1712622712
transform 1 0 3176 0 -1 770
box -5 -3 84 105
use INVX2  INVX2_0
timestamp 1712622712
transform 1 0 3352 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1712622712
transform 1 0 3256 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1712622712
transform 1 0 3328 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1712622712
transform 1 0 3136 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1712622712
transform 1 0 1480 0 1 970
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1712622712
transform 1 0 2784 0 1 170
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1712622712
transform 1 0 2936 0 1 170
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1712622712
transform 1 0 3008 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1712622712
transform 1 0 3256 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1712622712
transform 1 0 3408 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1712622712
transform 1 0 1440 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1712622712
transform 1 0 2960 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1712622712
transform 1 0 2960 0 1 970
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1712622712
transform 1 0 928 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1712622712
transform 1 0 1064 0 1 770
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1712622712
transform 1 0 1960 0 1 970
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1712622712
transform 1 0 2744 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1712622712
transform 1 0 1464 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1712622712
transform 1 0 768 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1712622712
transform 1 0 1768 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1712622712
transform 1 0 2848 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1712622712
transform 1 0 1504 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1712622712
transform 1 0 576 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1712622712
transform 1 0 1848 0 1 570
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1712622712
transform 1 0 2488 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1712622712
transform 1 0 2640 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1712622712
transform 1 0 1256 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1712622712
transform 1 0 1072 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1712622712
transform 1 0 1392 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1712622712
transform 1 0 1552 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1712622712
transform 1 0 2768 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1712622712
transform 1 0 1344 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1712622712
transform 1 0 2984 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1712622712
transform 1 0 728 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1712622712
transform 1 0 1544 0 1 570
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1712622712
transform 1 0 2384 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1712622712
transform 1 0 1280 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1712622712
transform 1 0 1560 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1712622712
transform 1 0 896 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1712622712
transform 1 0 1568 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1712622712
transform 1 0 2728 0 1 970
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1712622712
transform 1 0 3048 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1712622712
transform 1 0 1360 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1712622712
transform 1 0 1072 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1712622712
transform 1 0 1016 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1712622712
transform 1 0 1912 0 1 970
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1712622712
transform 1 0 2736 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1712622712
transform 1 0 912 0 1 970
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1712622712
transform 1 0 1728 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1712622712
transform 1 0 2720 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1712622712
transform 1 0 2632 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1712622712
transform 1 0 1536 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1712622712
transform 1 0 1672 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1712622712
transform 1 0 2776 0 1 570
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1712622712
transform 1 0 2728 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1712622712
transform 1 0 2704 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1712622712
transform 1 0 2400 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1712622712
transform 1 0 2744 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1712622712
transform 1 0 2544 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1712622712
transform 1 0 1008 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1712622712
transform 1 0 424 0 1 570
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1712622712
transform 1 0 1792 0 1 170
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1712622712
transform 1 0 2056 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1712622712
transform 1 0 2496 0 1 370
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1712622712
transform 1 0 536 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1712622712
transform 1 0 1408 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1712622712
transform 1 0 2944 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1712622712
transform 1 0 2656 0 1 370
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1712622712
transform 1 0 592 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1712622712
transform 1 0 2648 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1712622712
transform 1 0 2664 0 1 170
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1712622712
transform 1 0 1192 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1712622712
transform 1 0 312 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1712622712
transform 1 0 608 0 1 370
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1712622712
transform 1 0 2672 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1712622712
transform 1 0 2512 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1712622712
transform 1 0 976 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1712622712
transform 1 0 1544 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1712622712
transform 1 0 816 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1712622712
transform 1 0 544 0 1 570
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1712622712
transform 1 0 520 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1712622712
transform 1 0 2064 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1712622712
transform 1 0 1536 0 1 170
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1712622712
transform 1 0 2000 0 1 170
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1712622712
transform 1 0 2896 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1712622712
transform 1 0 2560 0 1 170
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1712622712
transform 1 0 840 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1712622712
transform 1 0 240 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1712622712
transform 1 0 744 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1712622712
transform 1 0 488 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1712622712
transform 1 0 680 0 1 370
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1712622712
transform 1 0 768 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1712622712
transform 1 0 2672 0 1 770
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1712622712
transform 1 0 3032 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1712622712
transform 1 0 2512 0 1 370
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1712622712
transform 1 0 808 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1712622712
transform 1 0 248 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1712622712
transform 1 0 480 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1712622712
transform 1 0 528 0 1 570
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1712622712
transform 1 0 1224 0 1 370
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1712622712
transform 1 0 1304 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1712622712
transform 1 0 2928 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1712622712
transform 1 0 2648 0 1 970
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1712622712
transform 1 0 1872 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1712622712
transform 1 0 2560 0 1 370
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1712622712
transform 1 0 1408 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1712622712
transform 1 0 1056 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1712622712
transform 1 0 584 0 1 370
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1712622712
transform 1 0 912 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1712622712
transform 1 0 496 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1712622712
transform 1 0 2576 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1712622712
transform 1 0 2408 0 1 370
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1712622712
transform 1 0 2528 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1712622712
transform 1 0 1696 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1712622712
transform 1 0 1088 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1712622712
transform 1 0 880 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1712622712
transform 1 0 544 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1712622712
transform 1 0 584 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1712622712
transform 1 0 416 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1712622712
transform 1 0 368 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1712622712
transform 1 0 384 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1712622712
transform 1 0 328 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1712622712
transform 1 0 200 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1712622712
transform 1 0 80 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1712622712
transform 1 0 192 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1712622712
transform 1 0 1016 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1712622712
transform 1 0 1128 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1712622712
transform 1 0 1224 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1712622712
transform 1 0 1344 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1712622712
transform 1 0 1328 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1712622712
transform 1 0 1496 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1712622712
transform 1 0 1608 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1712622712
transform 1 0 1848 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1712622712
transform 1 0 1720 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1712622712
transform 1 0 2072 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1712622712
transform 1 0 2128 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1712622712
transform 1 0 2336 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1712622712
transform 1 0 2016 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1712622712
transform 1 0 2400 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1712622712
transform 1 0 2712 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1712622712
transform 1 0 2720 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1712622712
transform 1 0 2560 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1712622712
transform 1 0 2824 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1712622712
transform 1 0 3176 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1712622712
transform 1 0 2688 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1712622712
transform 1 0 3088 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1712622712
transform 1 0 3048 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1712622712
transform 1 0 2976 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1712622712
transform 1 0 3248 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1712622712
transform 1 0 3280 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1712622712
transform 1 0 3072 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1712622712
transform 1 0 3312 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1712622712
transform 1 0 3192 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1712622712
transform 1 0 3400 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1712622712
transform 1 0 2832 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1712622712
transform 1 0 2904 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1712622712
transform 1 0 3032 0 1 570
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1712622712
transform 1 0 3168 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1712622712
transform 1 0 3344 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1712622712
transform 1 0 3208 0 1 770
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1712622712
transform 1 0 3288 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1712622712
transform 1 0 3184 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1712622712
transform 1 0 3288 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1712622712
transform 1 0 2040 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1712622712
transform 1 0 2224 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1712622712
transform 1 0 1960 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1712622712
transform 1 0 1960 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1712622712
transform 1 0 2048 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1712622712
transform 1 0 1984 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1712622712
transform 1 0 2144 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1712622712
transform 1 0 1912 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1712622712
transform 1 0 2304 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1712622712
transform 1 0 2208 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1712622712
transform 1 0 2280 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1712622712
transform 1 0 2240 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1712622712
transform 1 0 2400 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1712622712
transform 1 0 2392 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1712622712
transform 1 0 2488 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1712622712
transform 1 0 2496 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1712622712
transform 1 0 2488 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1712622712
transform 1 0 2560 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1712622712
transform 1 0 2424 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1712622712
transform 1 0 2032 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1712622712
transform 1 0 1680 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1712622712
transform 1 0 2640 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1712622712
transform 1 0 2440 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1712622712
transform 1 0 2416 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1712622712
transform 1 0 1344 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1712622712
transform 1 0 1632 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1712622712
transform 1 0 992 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1712622712
transform 1 0 992 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1712622712
transform 1 0 1456 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1712622712
transform 1 0 1024 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1712622712
transform 1 0 1664 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1712622712
transform 1 0 872 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1712622712
transform 1 0 2840 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1712622712
transform 1 0 1064 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1712622712
transform 1 0 1472 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1712622712
transform 1 0 1696 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1712622712
transform 1 0 712 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1712622712
transform 1 0 1376 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1712622712
transform 1 0 1208 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1712622712
transform 1 0 648 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1712622712
transform 1 0 800 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1712622712
transform 1 0 640 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1712622712
transform 1 0 1096 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1712622712
transform 1 0 568 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1712622712
transform 1 0 720 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1712622712
transform 1 0 512 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1712622712
transform 1 0 568 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1712622712
transform 1 0 552 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1712622712
transform 1 0 80 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1712622712
transform 1 0 496 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1712622712
transform 1 0 288 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1712622712
transform 1 0 528 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1712622712
transform 1 0 792 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1712622712
transform 1 0 168 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1712622712
transform 1 0 304 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1712622712
transform 1 0 728 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1712622712
transform 1 0 664 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1712622712
transform 1 0 496 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1712622712
transform 1 0 448 0 1 970
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1712622712
transform 1 0 96 0 1 970
box -9 -3 26 105
use INVX2  INVX2_223
timestamp 1712622712
transform 1 0 192 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1712622712
transform 1 0 368 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_225
timestamp 1712622712
transform 1 0 88 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_226
timestamp 1712622712
transform 1 0 672 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_227
timestamp 1712622712
transform 1 0 560 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_228
timestamp 1712622712
transform 1 0 88 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_229
timestamp 1712622712
transform 1 0 128 0 1 770
box -9 -3 26 105
use INVX2  INVX2_230
timestamp 1712622712
transform 1 0 728 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1712622712
transform 1 0 760 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_232
timestamp 1712622712
transform 1 0 1688 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1712622712
transform 1 0 880 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_234
timestamp 1712622712
transform 1 0 752 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_235
timestamp 1712622712
transform 1 0 688 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_236
timestamp 1712622712
transform 1 0 520 0 1 970
box -9 -3 26 105
use INVX2  INVX2_237
timestamp 1712622712
transform 1 0 448 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1712622712
transform 1 0 872 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_239
timestamp 1712622712
transform 1 0 2536 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1712622712
transform 1 0 520 0 1 170
box -9 -3 26 105
use INVX2  INVX2_241
timestamp 1712622712
transform 1 0 856 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_242
timestamp 1712622712
transform 1 0 1040 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_243
timestamp 1712622712
transform 1 0 432 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_244
timestamp 1712622712
transform 1 0 632 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_245
timestamp 1712622712
transform 1 0 760 0 1 570
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1712622712
transform 1 0 1080 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_247
timestamp 1712622712
transform 1 0 1160 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_248
timestamp 1712622712
transform 1 0 1176 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_249
timestamp 1712622712
transform 1 0 1120 0 1 570
box -9 -3 26 105
use INVX2  INVX2_250
timestamp 1712622712
transform 1 0 1240 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_251
timestamp 1712622712
transform 1 0 1352 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_252
timestamp 1712622712
transform 1 0 1328 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_253
timestamp 1712622712
transform 1 0 1056 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_254
timestamp 1712622712
transform 1 0 1216 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_255
timestamp 1712622712
transform 1 0 1312 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_256
timestamp 1712622712
transform 1 0 1272 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_257
timestamp 1712622712
transform 1 0 1528 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_258
timestamp 1712622712
transform 1 0 1368 0 1 370
box -9 -3 26 105
use INVX2  INVX2_259
timestamp 1712622712
transform 1 0 1456 0 1 570
box -9 -3 26 105
use INVX2  INVX2_260
timestamp 1712622712
transform 1 0 1616 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_261
timestamp 1712622712
transform 1 0 1544 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_262
timestamp 1712622712
transform 1 0 1664 0 1 170
box -9 -3 26 105
use INVX2  INVX2_263
timestamp 1712622712
transform 1 0 1680 0 1 370
box -9 -3 26 105
use INVX2  INVX2_264
timestamp 1712622712
transform 1 0 1872 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_265
timestamp 1712622712
transform 1 0 1840 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_266
timestamp 1712622712
transform 1 0 1752 0 1 570
box -9 -3 26 105
use INVX2  INVX2_267
timestamp 1712622712
transform 1 0 1672 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_268
timestamp 1712622712
transform 1 0 2040 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_269
timestamp 1712622712
transform 1 0 2112 0 1 370
box -9 -3 26 105
use INVX2  INVX2_270
timestamp 1712622712
transform 1 0 2032 0 1 370
box -9 -3 26 105
use INVX2  INVX2_271
timestamp 1712622712
transform 1 0 1856 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_272
timestamp 1712622712
transform 1 0 1760 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_273
timestamp 1712622712
transform 1 0 2032 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_274
timestamp 1712622712
transform 1 0 1840 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_275
timestamp 1712622712
transform 1 0 1560 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_276
timestamp 1712622712
transform 1 0 1672 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_277
timestamp 1712622712
transform 1 0 2720 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_278
timestamp 1712622712
transform 1 0 2096 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_279
timestamp 1712622712
transform 1 0 1832 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_280
timestamp 1712622712
transform 1 0 2208 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_281
timestamp 1712622712
transform 1 0 1840 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_282
timestamp 1712622712
transform 1 0 992 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_283
timestamp 1712622712
transform 1 0 2424 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_284
timestamp 1712622712
transform 1 0 2200 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_285
timestamp 1712622712
transform 1 0 2416 0 1 770
box -9 -3 26 105
use INVX2  INVX2_286
timestamp 1712622712
transform 1 0 2104 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_287
timestamp 1712622712
transform 1 0 2176 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_288
timestamp 1712622712
transform 1 0 2448 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_289
timestamp 1712622712
transform 1 0 2256 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_290
timestamp 1712622712
transform 1 0 2272 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_291
timestamp 1712622712
transform 1 0 2488 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_292
timestamp 1712622712
transform 1 0 2800 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_293
timestamp 1712622712
transform 1 0 2464 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_294
timestamp 1712622712
transform 1 0 3408 0 1 770
box -9 -3 26 105
use INVX2  INVX2_295
timestamp 1712622712
transform 1 0 3272 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_296
timestamp 1712622712
transform 1 0 3296 0 1 770
box -9 -3 26 105
use INVX2  INVX2_297
timestamp 1712622712
transform 1 0 3288 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_298
timestamp 1712622712
transform 1 0 3384 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_299
timestamp 1712622712
transform 1 0 3344 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_300
timestamp 1712622712
transform 1 0 3400 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_301
timestamp 1712622712
transform 1 0 3400 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_302
timestamp 1712622712
transform 1 0 3304 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_303
timestamp 1712622712
transform 1 0 2952 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_304
timestamp 1712622712
transform 1 0 3256 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_305
timestamp 1712622712
transform 1 0 2792 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_306
timestamp 1712622712
transform 1 0 2368 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_307
timestamp 1712622712
transform 1 0 3136 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_308
timestamp 1712622712
transform 1 0 1288 0 1 970
box -9 -3 26 105
use INVX2  INVX2_309
timestamp 1712622712
transform 1 0 3208 0 1 170
box -9 -3 26 105
use INVX2  INVX2_310
timestamp 1712622712
transform 1 0 2432 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_311
timestamp 1712622712
transform 1 0 1264 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_312
timestamp 1712622712
transform 1 0 2944 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_313
timestamp 1712622712
transform 1 0 2344 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_314
timestamp 1712622712
transform 1 0 2616 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_315
timestamp 1712622712
transform 1 0 2584 0 1 770
box -9 -3 26 105
use INVX2  INVX2_316
timestamp 1712622712
transform 1 0 2672 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_317
timestamp 1712622712
transform 1 0 2824 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_318
timestamp 1712622712
transform 1 0 1704 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_319
timestamp 1712622712
transform 1 0 2632 0 1 970
box -9 -3 26 105
use INVX2  INVX2_320
timestamp 1712622712
transform 1 0 2584 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_321
timestamp 1712622712
transform 1 0 3248 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_322
timestamp 1712622712
transform 1 0 328 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_323
timestamp 1712622712
transform 1 0 312 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_324
timestamp 1712622712
transform 1 0 472 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_325
timestamp 1712622712
transform 1 0 2264 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_326
timestamp 1712622712
transform 1 0 1568 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_327
timestamp 1712622712
transform 1 0 2728 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_328
timestamp 1712622712
transform 1 0 752 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_329
timestamp 1712622712
transform 1 0 2960 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_330
timestamp 1712622712
transform 1 0 3024 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_331
timestamp 1712622712
transform 1 0 2832 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_332
timestamp 1712622712
transform 1 0 2584 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_333
timestamp 1712622712
transform 1 0 2824 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_334
timestamp 1712622712
transform 1 0 2480 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_335
timestamp 1712622712
transform 1 0 2552 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_336
timestamp 1712622712
transform 1 0 2536 0 1 770
box -9 -3 26 105
use INVX2  INVX2_337
timestamp 1712622712
transform 1 0 2584 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_338
timestamp 1712622712
transform 1 0 3256 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_339
timestamp 1712622712
transform 1 0 3200 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_340
timestamp 1712622712
transform 1 0 3240 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_341
timestamp 1712622712
transform 1 0 3008 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_342
timestamp 1712622712
transform 1 0 1272 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_343
timestamp 1712622712
transform 1 0 2512 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_344
timestamp 1712622712
transform 1 0 2808 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_345
timestamp 1712622712
transform 1 0 2360 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_346
timestamp 1712622712
transform 1 0 2472 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_347
timestamp 1712622712
transform 1 0 2936 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_348
timestamp 1712622712
transform 1 0 1712 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_349
timestamp 1712622712
transform 1 0 2568 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_350
timestamp 1712622712
transform 1 0 3408 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_351
timestamp 1712622712
transform 1 0 3208 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_352
timestamp 1712622712
transform 1 0 3352 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_353
timestamp 1712622712
transform 1 0 3400 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_354
timestamp 1712622712
transform 1 0 3304 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_355
timestamp 1712622712
transform 1 0 3392 0 -1 2370
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1712622712
transform 1 0 3204 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1712622712
transform 1 0 3092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1712622712
transform 1 0 3108 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1712622712
transform 1 0 2876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1712622712
transform 1 0 2900 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1712622712
transform 1 0 2892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1712622712
transform 1 0 3140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1712622712
transform 1 0 2988 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1712622712
transform 1 0 2988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1712622712
transform 1 0 2924 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1712622712
transform 1 0 2884 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1712622712
transform 1 0 2852 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1712622712
transform 1 0 3140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1712622712
transform 1 0 2980 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1712622712
transform 1 0 2964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1712622712
transform 1 0 2940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1712622712
transform 1 0 2924 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1712622712
transform 1 0 2828 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1712622712
transform 1 0 2812 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1712622712
transform 1 0 3060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1712622712
transform 1 0 2988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1712622712
transform 1 0 2964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1712622712
transform 1 0 2852 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1712622712
transform 1 0 2812 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1712622712
transform 1 0 2804 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1712622712
transform 1 0 2836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1712622712
transform 1 0 2772 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1712622712
transform 1 0 1412 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1712622712
transform 1 0 1380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1712622712
transform 1 0 2868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1712622712
transform 1 0 2804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1712622712
transform 1 0 1524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1712622712
transform 1 0 1420 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1712622712
transform 1 0 1364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1712622712
transform 1 0 3268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1712622712
transform 1 0 2980 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1712622712
transform 1 0 2684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1712622712
transform 1 0 2676 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1712622712
transform 1 0 2668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1712622712
transform 1 0 2588 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1712622712
transform 1 0 2564 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1712622712
transform 1 0 2404 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1712622712
transform 1 0 1972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1712622712
transform 1 0 1964 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1712622712
transform 1 0 1380 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1712622712
transform 1 0 1300 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1712622712
transform 1 0 1292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1712622712
transform 1 0 1084 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1712622712
transform 1 0 1028 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1712622712
transform 1 0 740 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1712622712
transform 1 0 708 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1712622712
transform 1 0 700 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1712622712
transform 1 0 684 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1712622712
transform 1 0 668 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1712622712
transform 1 0 652 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1712622712
transform 1 0 596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1712622712
transform 1 0 596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1712622712
transform 1 0 3188 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1712622712
transform 1 0 2964 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1712622712
transform 1 0 2684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1712622712
transform 1 0 2684 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1712622712
transform 1 0 2628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1712622712
transform 1 0 3276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1712622712
transform 1 0 3252 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1712622712
transform 1 0 3236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1712622712
transform 1 0 3132 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1712622712
transform 1 0 3100 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1712622712
transform 1 0 2988 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1712622712
transform 1 0 2956 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1712622712
transform 1 0 2932 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1712622712
transform 1 0 2868 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1712622712
transform 1 0 3036 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1712622712
transform 1 0 3004 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1712622712
transform 1 0 2932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1712622712
transform 1 0 2876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1712622712
transform 1 0 2892 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1712622712
transform 1 0 2788 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1712622712
transform 1 0 2788 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1712622712
transform 1 0 3404 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1712622712
transform 1 0 3300 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1712622712
transform 1 0 3292 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1712622712
transform 1 0 3284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1712622712
transform 1 0 3260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1712622712
transform 1 0 3420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1712622712
transform 1 0 3348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1712622712
transform 1 0 3284 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1712622712
transform 1 0 2692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1712622712
transform 1 0 2692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1712622712
transform 1 0 2980 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1712622712
transform 1 0 2916 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1712622712
transform 1 0 3188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1712622712
transform 1 0 3180 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1712622712
transform 1 0 2900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1712622712
transform 1 0 2828 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1712622712
transform 1 0 2692 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1712622712
transform 1 0 2564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1712622712
transform 1 0 2772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1712622712
transform 1 0 2724 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1712622712
transform 1 0 2820 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1712622712
transform 1 0 2716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1712622712
transform 1 0 2508 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1712622712
transform 1 0 2404 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1712622712
transform 1 0 2148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1712622712
transform 1 0 2020 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1712622712
transform 1 0 2236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1712622712
transform 1 0 2132 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1712622712
transform 1 0 1772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1712622712
transform 1 0 1724 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1712622712
transform 1 0 1924 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1712622712
transform 1 0 1852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1712622712
transform 1 0 1612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1712622712
transform 1 0 1612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1712622712
transform 1 0 1564 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1712622712
transform 1 0 1500 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1712622712
transform 1 0 1444 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1712622712
transform 1 0 1332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1712622712
transform 1 0 1468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1712622712
transform 1 0 1348 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1712622712
transform 1 0 1292 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1712622712
transform 1 0 1228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1712622712
transform 1 0 1148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1712622712
transform 1 0 1020 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1712622712
transform 1 0 228 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1712622712
transform 1 0 84 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1712622712
transform 1 0 3388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1712622712
transform 1 0 3348 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1712622712
transform 1 0 3292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1712622712
transform 1 0 3276 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1712622712
transform 1 0 3428 0 1 2455
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1712622712
transform 1 0 3292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1712622712
transform 1 0 3436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1712622712
transform 1 0 3388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1712622712
transform 1 0 3196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1712622712
transform 1 0 3156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1712622712
transform 1 0 3428 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1712622712
transform 1 0 3404 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1712622712
transform 1 0 3396 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1712622712
transform 1 0 3332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1712622712
transform 1 0 3052 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1712622712
transform 1 0 2828 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1712622712
transform 1 0 3364 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1712622712
transform 1 0 3348 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1712622712
transform 1 0 3332 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1712622712
transform 1 0 3324 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1712622712
transform 1 0 3044 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1712622712
transform 1 0 2980 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1712622712
transform 1 0 2756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1712622712
transform 1 0 2668 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1712622712
transform 1 0 2948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1712622712
transform 1 0 2884 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1712622712
transform 1 0 3052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1712622712
transform 1 0 2828 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1712622712
transform 1 0 2852 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1712622712
transform 1 0 2740 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1712622712
transform 1 0 2652 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1712622712
transform 1 0 2596 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1712622712
transform 1 0 2556 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1712622712
transform 1 0 2508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1712622712
transform 1 0 2460 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1712622712
transform 1 0 2388 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1712622712
transform 1 0 2164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1712622712
transform 1 0 2140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1712622712
transform 1 0 1964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1712622712
transform 1 0 1964 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1712622712
transform 1 0 2260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1712622712
transform 1 0 2220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1712622712
transform 1 0 2356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1712622712
transform 1 0 2316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1712622712
transform 1 0 2060 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1712622712
transform 1 0 2036 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1712622712
transform 1 0 1860 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1712622712
transform 1 0 1836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1712622712
transform 1 0 1748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1712622712
transform 1 0 1732 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1712622712
transform 1 0 1628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1712622712
transform 1 0 1620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1712622712
transform 1 0 1484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1712622712
transform 1 0 1460 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1712622712
transform 1 0 1444 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1712622712
transform 1 0 1356 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1712622712
transform 1 0 1188 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1712622712
transform 1 0 1140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1712622712
transform 1 0 1060 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1712622712
transform 1 0 956 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1712622712
transform 1 0 764 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1712622712
transform 1 0 628 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1712622712
transform 1 0 180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1712622712
transform 1 0 156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1712622712
transform 1 0 180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1712622712
transform 1 0 84 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1712622712
transform 1 0 236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1712622712
transform 1 0 236 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1712622712
transform 1 0 292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1712622712
transform 1 0 292 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1712622712
transform 1 0 412 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1712622712
transform 1 0 412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1712622712
transform 1 0 508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1712622712
transform 1 0 500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1712622712
transform 1 0 724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1712622712
transform 1 0 612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1712622712
transform 1 0 836 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1712622712
transform 1 0 716 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1712622712
transform 1 0 948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1712622712
transform 1 0 868 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1712622712
transform 1 0 1244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1712622712
transform 1 0 1148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1712622712
transform 1 0 2740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1712622712
transform 1 0 2740 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1712622712
transform 1 0 2972 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1712622712
transform 1 0 2924 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1712622712
transform 1 0 3036 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1712622712
transform 1 0 2876 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1712622712
transform 1 0 2844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1712622712
transform 1 0 2828 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1712622712
transform 1 0 2660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1712622712
transform 1 0 2636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1712622712
transform 1 0 2612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1712622712
transform 1 0 2596 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1712622712
transform 1 0 2548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1712622712
transform 1 0 2444 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1712622712
transform 1 0 2436 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1712622712
transform 1 0 2204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1712622712
transform 1 0 2004 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1712622712
transform 1 0 2004 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1712622712
transform 1 0 2308 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1712622712
transform 1 0 2260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1712622712
transform 1 0 2348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1712622712
transform 1 0 2268 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1712622712
transform 1 0 2116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1712622712
transform 1 0 2108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1712622712
transform 1 0 1884 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1712622712
transform 1 0 1884 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1712622712
transform 1 0 1996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1712622712
transform 1 0 1828 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1712622712
transform 1 0 1772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1712622712
transform 1 0 1716 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1712622712
transform 1 0 1660 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1712622712
transform 1 0 1660 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1712622712
transform 1 0 1532 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1712622712
transform 1 0 1532 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1712622712
transform 1 0 1476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1712622712
transform 1 0 1436 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1712622712
transform 1 0 1308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1712622712
transform 1 0 1244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1712622712
transform 1 0 1084 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1712622712
transform 1 0 1020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1712622712
transform 1 0 988 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1712622712
transform 1 0 860 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1712622712
transform 1 0 204 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1712622712
transform 1 0 204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1712622712
transform 1 0 172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1712622712
transform 1 0 148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1712622712
transform 1 0 284 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1712622712
transform 1 0 284 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1712622712
transform 1 0 332 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1712622712
transform 1 0 332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1712622712
transform 1 0 396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1712622712
transform 1 0 364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1712622712
transform 1 0 444 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1712622712
transform 1 0 444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1712622712
transform 1 0 532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1712622712
transform 1 0 492 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1712622712
transform 1 0 660 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1712622712
transform 1 0 652 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1712622712
transform 1 0 764 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1712622712
transform 1 0 756 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1712622712
transform 1 0 908 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1712622712
transform 1 0 884 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1712622712
transform 1 0 1196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1712622712
transform 1 0 1196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1712622712
transform 1 0 3348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1712622712
transform 1 0 3204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1712622712
transform 1 0 3196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1712622712
transform 1 0 3180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1712622712
transform 1 0 3172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1712622712
transform 1 0 3124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1712622712
transform 1 0 3100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1712622712
transform 1 0 3244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1712622712
transform 1 0 3204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1712622712
transform 1 0 3196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1712622712
transform 1 0 3188 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1712622712
transform 1 0 3164 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1712622712
transform 1 0 3164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1712622712
transform 1 0 3148 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1712622712
transform 1 0 3116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1712622712
transform 1 0 3108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1712622712
transform 1 0 3100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1712622712
transform 1 0 3068 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1712622712
transform 1 0 3028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1712622712
transform 1 0 3028 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1712622712
transform 1 0 3012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1712622712
transform 1 0 2964 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1712622712
transform 1 0 2916 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1712622712
transform 1 0 2908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1712622712
transform 1 0 2844 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1712622712
transform 1 0 2804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1712622712
transform 1 0 2948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1712622712
transform 1 0 2884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1712622712
transform 1 0 2828 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1712622712
transform 1 0 2828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1712622712
transform 1 0 2828 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1712622712
transform 1 0 3404 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1712622712
transform 1 0 3396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1712622712
transform 1 0 3188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1712622712
transform 1 0 3188 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1712622712
transform 1 0 3308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1712622712
transform 1 0 3252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1712622712
transform 1 0 3148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1712622712
transform 1 0 3404 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1712622712
transform 1 0 3404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1712622712
transform 1 0 3380 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1712622712
transform 1 0 3380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1712622712
transform 1 0 3340 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1712622712
transform 1 0 3348 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1712622712
transform 1 0 3348 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1712622712
transform 1 0 3300 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1712622712
transform 1 0 3300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1712622712
transform 1 0 3428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1712622712
transform 1 0 3364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1712622712
transform 1 0 3252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1712622712
transform 1 0 3236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1712622712
transform 1 0 3420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1712622712
transform 1 0 3348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1712622712
transform 1 0 3316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1712622712
transform 1 0 3316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1712622712
transform 1 0 3228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1712622712
transform 1 0 3212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1712622712
transform 1 0 3196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1712622712
transform 1 0 3148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1712622712
transform 1 0 3068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1712622712
transform 1 0 3036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1712622712
transform 1 0 2980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1712622712
transform 1 0 2892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1712622712
transform 1 0 2844 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1712622712
transform 1 0 2812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1712622712
transform 1 0 3332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1712622712
transform 1 0 3316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1712622712
transform 1 0 3300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1712622712
transform 1 0 3284 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1712622712
transform 1 0 3220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1712622712
transform 1 0 3220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1712622712
transform 1 0 3204 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1712622712
transform 1 0 3180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1712622712
transform 1 0 3172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1712622712
transform 1 0 3148 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1712622712
transform 1 0 3148 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1712622712
transform 1 0 3420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1712622712
transform 1 0 3300 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1712622712
transform 1 0 3284 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1712622712
transform 1 0 3164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1712622712
transform 1 0 3164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1712622712
transform 1 0 3268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1712622712
transform 1 0 3252 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1712622712
transform 1 0 3220 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1712622712
transform 1 0 3212 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1712622712
transform 1 0 3212 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1712622712
transform 1 0 3164 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1712622712
transform 1 0 3140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1712622712
transform 1 0 3140 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1712622712
transform 1 0 2948 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1712622712
transform 1 0 2916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1712622712
transform 1 0 3188 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1712622712
transform 1 0 3100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1712622712
transform 1 0 3036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1712622712
transform 1 0 3196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1712622712
transform 1 0 3156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1712622712
transform 1 0 3156 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1712622712
transform 1 0 3156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1712622712
transform 1 0 3252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1712622712
transform 1 0 3172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1712622712
transform 1 0 2676 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1712622712
transform 1 0 2604 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1712622712
transform 1 0 2404 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1712622712
transform 1 0 1668 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1712622712
transform 1 0 1452 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1712622712
transform 1 0 1268 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1712622712
transform 1 0 3396 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1712622712
transform 1 0 3276 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1712622712
transform 1 0 3260 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1712622712
transform 1 0 3260 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1712622712
transform 1 0 3268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1712622712
transform 1 0 3172 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1712622712
transform 1 0 3068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1712622712
transform 1 0 3068 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1712622712
transform 1 0 2964 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1712622712
transform 1 0 2956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1712622712
transform 1 0 3332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1712622712
transform 1 0 3332 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1712622712
transform 1 0 3324 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1712622712
transform 1 0 3308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1712622712
transform 1 0 3300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1712622712
transform 1 0 3284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1712622712
transform 1 0 3228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1712622712
transform 1 0 3124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1712622712
transform 1 0 3124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1712622712
transform 1 0 3068 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1712622712
transform 1 0 3012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1712622712
transform 1 0 2788 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1712622712
transform 1 0 2684 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1712622712
transform 1 0 2644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1712622712
transform 1 0 2612 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1712622712
transform 1 0 2420 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1712622712
transform 1 0 2252 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1712622712
transform 1 0 1908 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1712622712
transform 1 0 1820 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1712622712
transform 1 0 1748 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1712622712
transform 1 0 1748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1712622712
transform 1 0 1684 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1712622712
transform 1 0 1396 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1712622712
transform 1 0 1324 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1712622712
transform 1 0 1044 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1712622712
transform 1 0 1028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1712622712
transform 1 0 852 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1712622712
transform 1 0 796 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1712622712
transform 1 0 796 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1712622712
transform 1 0 2660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1712622712
transform 1 0 2580 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1712622712
transform 1 0 2540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1712622712
transform 1 0 2404 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1712622712
transform 1 0 2348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1712622712
transform 1 0 2124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1712622712
transform 1 0 1556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1712622712
transform 1 0 1484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1712622712
transform 1 0 1476 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1712622712
transform 1 0 1468 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1712622712
transform 1 0 1452 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1712622712
transform 1 0 1396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1712622712
transform 1 0 1396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1712622712
transform 1 0 1340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1712622712
transform 1 0 1300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1712622712
transform 1 0 1020 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1712622712
transform 1 0 972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1712622712
transform 1 0 932 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1712622712
transform 1 0 932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1712622712
transform 1 0 1492 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1712622712
transform 1 0 1492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1712622712
transform 1 0 1452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1712622712
transform 1 0 1156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1712622712
transform 1 0 2860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1712622712
transform 1 0 2772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1712622712
transform 1 0 2748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1712622712
transform 1 0 3028 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1712622712
transform 1 0 2932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1712622712
transform 1 0 2908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1712622712
transform 1 0 3108 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1712622712
transform 1 0 3076 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1712622712
transform 1 0 3316 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1712622712
transform 1 0 3316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1712622712
transform 1 0 3252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1712622712
transform 1 0 3188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1712622712
transform 1 0 3428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1712622712
transform 1 0 3428 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1712622712
transform 1 0 3380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1712622712
transform 1 0 3332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1712622712
transform 1 0 2948 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1712622712
transform 1 0 2948 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1712622712
transform 1 0 2932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1712622712
transform 1 0 2868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1712622712
transform 1 0 2844 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1712622712
transform 1 0 2844 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1712622712
transform 1 0 2812 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1712622712
transform 1 0 2812 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1712622712
transform 1 0 2804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1712622712
transform 1 0 2804 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1712622712
transform 1 0 2772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1712622712
transform 1 0 2748 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1712622712
transform 1 0 2740 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1712622712
transform 1 0 1500 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1712622712
transform 1 0 1436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1712622712
transform 1 0 1428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1712622712
transform 1 0 2540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1712622712
transform 1 0 2452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1712622712
transform 1 0 2452 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1712622712
transform 1 0 2420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1712622712
transform 1 0 2372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1712622712
transform 1 0 2220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1712622712
transform 1 0 2060 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1712622712
transform 1 0 1980 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1712622712
transform 1 0 1980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1712622712
transform 1 0 1924 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1712622712
transform 1 0 1892 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1712622712
transform 1 0 1812 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1712622712
transform 1 0 1700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1712622712
transform 1 0 1628 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1712622712
transform 1 0 1628 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1712622712
transform 1 0 1604 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1712622712
transform 1 0 1596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1712622712
transform 1 0 2940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1712622712
transform 1 0 2884 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1712622712
transform 1 0 2884 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1712622712
transform 1 0 2860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1712622712
transform 1 0 2852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1712622712
transform 1 0 2948 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1712622712
transform 1 0 2876 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1712622712
transform 1 0 2876 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1712622712
transform 1 0 2844 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1712622712
transform 1 0 2836 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1712622712
transform 1 0 2796 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1712622712
transform 1 0 1020 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1712622712
transform 1 0 924 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1712622712
transform 1 0 868 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1712622712
transform 1 0 1268 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1712622712
transform 1 0 1060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1712622712
transform 1 0 1036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1712622712
transform 1 0 1036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1712622712
transform 1 0 1036 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1712622712
transform 1 0 828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1712622712
transform 1 0 2004 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1712622712
transform 1 0 1932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1712622712
transform 1 0 1868 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1712622712
transform 1 0 1740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1712622712
transform 1 0 1740 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1712622712
transform 1 0 2700 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1712622712
transform 1 0 2652 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1712622712
transform 1 0 1476 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1712622712
transform 1 0 1420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1712622712
transform 1 0 772 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1712622712
transform 1 0 692 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1712622712
transform 1 0 628 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1712622712
transform 1 0 1780 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1712622712
transform 1 0 1780 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1712622712
transform 1 0 1748 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1712622712
transform 1 0 1644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1712622712
transform 1 0 1644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1712622712
transform 1 0 3036 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1712622712
transform 1 0 2932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1712622712
transform 1 0 2844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1712622712
transform 1 0 2796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1712622712
transform 1 0 2620 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1712622712
transform 1 0 2436 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1712622712
transform 1 0 2436 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1712622712
transform 1 0 2420 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1712622712
transform 1 0 2404 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1712622712
transform 1 0 2396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1712622712
transform 1 0 1652 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1712622712
transform 1 0 1556 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1712622712
transform 1 0 1556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1712622712
transform 1 0 1524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1712622712
transform 1 0 1460 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1712622712
transform 1 0 1460 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1712622712
transform 1 0 596 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1712622712
transform 1 0 596 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1712622712
transform 1 0 1900 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1712622712
transform 1 0 1804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1712622712
transform 1 0 1780 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1712622712
transform 1 0 2652 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1712622712
transform 1 0 2564 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1712622712
transform 1 0 2468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1712622712
transform 1 0 2460 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1712622712
transform 1 0 2764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1712622712
transform 1 0 2668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1712622712
transform 1 0 1268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1712622712
transform 1 0 1268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1712622712
transform 1 0 1092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1712622712
transform 1 0 1092 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1712622712
transform 1 0 876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1712622712
transform 1 0 1396 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1712622712
transform 1 0 1164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1712622712
transform 1 0 2660 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1712622712
transform 1 0 1564 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1712622712
transform 1 0 1540 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1712622712
transform 1 0 2980 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1712622712
transform 1 0 2724 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1712622712
transform 1 0 1916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1712622712
transform 1 0 1524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1712622712
transform 1 0 1380 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1712622712
transform 1 0 1324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1712622712
transform 1 0 1276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1712622712
transform 1 0 1212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1712622712
transform 1 0 1188 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1712622712
transform 1 0 2980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1712622712
transform 1 0 2900 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1712622712
transform 1 0 2844 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1712622712
transform 1 0 2804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1712622712
transform 1 0 2796 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1712622712
transform 1 0 740 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1712622712
transform 1 0 708 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1712622712
transform 1 0 1620 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1712622712
transform 1 0 1556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1712622712
transform 1 0 1524 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1712622712
transform 1 0 2372 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1712622712
transform 1 0 2372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1712622712
transform 1 0 2348 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1712622712
transform 1 0 1284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1712622712
transform 1 0 1260 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1712622712
transform 1 0 908 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1712622712
transform 1 0 900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1712622712
transform 1 0 732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1712622712
transform 1 0 692 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1712622712
transform 1 0 1588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1712622712
transform 1 0 1580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1712622712
transform 1 0 1516 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1712622712
transform 1 0 1364 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1712622712
transform 1 0 1284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1712622712
transform 1 0 2780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1712622712
transform 1 0 2740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1712622712
transform 1 0 1708 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1712622712
transform 1 0 3076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1712622712
transform 1 0 3076 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1712622712
transform 1 0 3076 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1712622712
transform 1 0 2996 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1712622712
transform 1 0 2332 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1712622712
transform 1 0 2156 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1712622712
transform 1 0 2156 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1712622712
transform 1 0 1420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1712622712
transform 1 0 1364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1712622712
transform 1 0 1364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1712622712
transform 1 0 1324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1712622712
transform 1 0 1244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1712622712
transform 1 0 1084 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1712622712
transform 1 0 1084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1712622712
transform 1 0 1052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1712622712
transform 1 0 1044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1712622712
transform 1 0 1092 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1712622712
transform 1 0 1004 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1712622712
transform 1 0 812 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1712622712
transform 1 0 668 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1712622712
transform 1 0 644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1712622712
transform 1 0 1956 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1712622712
transform 1 0 1900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1712622712
transform 1 0 1852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1712622712
transform 1 0 1812 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1712622712
transform 1 0 1812 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1712622712
transform 1 0 2868 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1712622712
transform 1 0 2852 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1712622712
transform 1 0 2764 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1712622712
transform 1 0 2748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1712622712
transform 1 0 2580 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1712622712
transform 1 0 2540 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1712622712
transform 1 0 2540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1712622712
transform 1 0 1100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1712622712
transform 1 0 900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1712622712
transform 1 0 708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1712622712
transform 1 0 1820 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1712622712
transform 1 0 1740 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1712622712
transform 1 0 1460 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1712622712
transform 1 0 2700 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1712622712
transform 1 0 2676 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1712622712
transform 1 0 2596 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1712622712
transform 1 0 2740 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1712622712
transform 1 0 2628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1712622712
transform 1 0 1596 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1712622712
transform 1 0 1596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1712622712
transform 1 0 1580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1712622712
transform 1 0 1580 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1712622712
transform 1 0 1524 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1712622712
transform 1 0 1524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1712622712
transform 1 0 1660 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1712622712
transform 1 0 1660 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1712622712
transform 1 0 3372 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1712622712
transform 1 0 3324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1712622712
transform 1 0 3260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1712622712
transform 1 0 3252 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1712622712
transform 1 0 3148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1712622712
transform 1 0 3092 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1712622712
transform 1 0 3092 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1712622712
transform 1 0 2924 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1712622712
transform 1 0 2868 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1712622712
transform 1 0 2764 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1712622712
transform 1 0 2740 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1712622712
transform 1 0 2812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1712622712
transform 1 0 2812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1712622712
transform 1 0 2764 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1712622712
transform 1 0 2708 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1712622712
transform 1 0 3028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1712622712
transform 1 0 2740 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1712622712
transform 1 0 2740 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1712622712
transform 1 0 2676 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1712622712
transform 1 0 2692 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1712622712
transform 1 0 2692 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1712622712
transform 1 0 2588 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1712622712
transform 1 0 2564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1712622712
transform 1 0 2540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1712622712
transform 1 0 2428 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1712622712
transform 1 0 2396 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1712622712
transform 1 0 3156 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1712622712
transform 1 0 2756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1712622712
transform 1 0 2676 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1712622712
transform 1 0 2652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1712622712
transform 1 0 2612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1712622712
transform 1 0 2580 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1712622712
transform 1 0 2580 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1712622712
transform 1 0 2500 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1712622712
transform 1 0 1380 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1712622712
transform 1 0 1340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1712622712
transform 1 0 1188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1712622712
transform 1 0 1156 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1712622712
transform 1 0 1044 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1712622712
transform 1 0 1020 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1712622712
transform 1 0 900 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1712622712
transform 1 0 884 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1712622712
transform 1 0 644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1712622712
transform 1 0 508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1712622712
transform 1 0 1244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1712622712
transform 1 0 884 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1712622712
transform 1 0 516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1712622712
transform 1 0 436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1712622712
transform 1 0 236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1712622712
transform 1 0 228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1712622712
transform 1 0 148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1712622712
transform 1 0 132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1712622712
transform 1 0 1788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1712622712
transform 1 0 1764 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1712622712
transform 1 0 1740 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1712622712
transform 1 0 1628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1712622712
transform 1 0 1628 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1712622712
transform 1 0 1580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1712622712
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1712622712
transform 1 0 2108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1712622712
transform 1 0 2100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1712622712
transform 1 0 2092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1712622712
transform 1 0 2068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1712622712
transform 1 0 2060 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1712622712
transform 1 0 2044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1712622712
transform 1 0 2036 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1712622712
transform 1 0 2036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1712622712
transform 1 0 2012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1712622712
transform 1 0 2516 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1712622712
transform 1 0 2492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1712622712
transform 1 0 2372 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1712622712
transform 1 0 1108 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1712622712
transform 1 0 1060 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1712622712
transform 1 0 1372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1712622712
transform 1 0 1284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1712622712
transform 1 0 676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1712622712
transform 1 0 620 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1712622712
transform 1 0 580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1712622712
transform 1 0 1380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1712622712
transform 1 0 1356 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1712622712
transform 1 0 1332 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1712622712
transform 1 0 1012 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1712622712
transform 1 0 884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1712622712
transform 1 0 772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1712622712
transform 1 0 676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1712622712
transform 1 0 3132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1712622712
transform 1 0 3068 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1712622712
transform 1 0 2900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1712622712
transform 1 0 2724 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1712622712
transform 1 0 2276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1712622712
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1712622712
transform 1 0 1900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1712622712
transform 1 0 2652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1712622712
transform 1 0 2628 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1712622712
transform 1 0 2284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1712622712
transform 1 0 1300 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1712622712
transform 1 0 1244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1712622712
transform 1 0 1292 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1712622712
transform 1 0 1244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1712622712
transform 1 0 1140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1712622712
transform 1 0 964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1712622712
transform 1 0 900 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1712622712
transform 1 0 604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1712622712
transform 1 0 588 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1712622712
transform 1 0 500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1712622712
transform 1 0 3004 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1712622712
transform 1 0 2660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1712622712
transform 1 0 2444 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1712622712
transform 1 0 2380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1712622712
transform 1 0 2252 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1712622712
transform 1 0 2252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1712622712
transform 1 0 2700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1712622712
transform 1 0 2700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1712622712
transform 1 0 2676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1712622712
transform 1 0 2484 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1712622712
transform 1 0 1244 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1712622712
transform 1 0 1228 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1712622712
transform 1 0 1324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1712622712
transform 1 0 1268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1712622712
transform 1 0 1196 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1712622712
transform 1 0 1196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1712622712
transform 1 0 1164 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1712622712
transform 1 0 1612 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1712622712
transform 1 0 932 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1712622712
transform 1 0 876 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1712622712
transform 1 0 732 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1712622712
transform 1 0 668 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1712622712
transform 1 0 324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1712622712
transform 1 0 324 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1712622712
transform 1 0 324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1712622712
transform 1 0 276 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1712622712
transform 1 0 604 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1712622712
transform 1 0 564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1712622712
transform 1 0 188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1712622712
transform 1 0 100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1712622712
transform 1 0 2644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1712622712
transform 1 0 2620 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1712622712
transform 1 0 2612 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1712622712
transform 1 0 2588 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1712622712
transform 1 0 2588 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1712622712
transform 1 0 2564 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1712622712
transform 1 0 2524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1712622712
transform 1 0 2516 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1712622712
transform 1 0 2508 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1712622712
transform 1 0 1124 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1712622712
transform 1 0 1092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1712622712
transform 1 0 1076 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1712622712
transform 1 0 972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1712622712
transform 1 0 972 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1712622712
transform 1 0 940 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1712622712
transform 1 0 1596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1712622712
transform 1 0 1556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1712622712
transform 1 0 1228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1712622712
transform 1 0 836 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1712622712
transform 1 0 116 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1712622712
transform 1 0 100 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1712622712
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1712622712
transform 1 0 532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1712622712
transform 1 0 412 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1712622712
transform 1 0 412 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1712622712
transform 1 0 356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1712622712
transform 1 0 540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1712622712
transform 1 0 516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1712622712
transform 1 0 436 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1712622712
transform 1 0 420 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1712622712
transform 1 0 388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1712622712
transform 1 0 2052 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1712622712
transform 1 0 2020 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1712622712
transform 1 0 2012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1712622712
transform 1 0 2004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1712622712
transform 1 0 1780 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1712622712
transform 1 0 1556 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1712622712
transform 1 0 1556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1712622712
transform 1 0 1500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1712622712
transform 1 0 1284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1712622712
transform 1 0 1244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1712622712
transform 1 0 1212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1712622712
transform 1 0 1956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1712622712
transform 1 0 1924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1712622712
transform 1 0 2932 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1712622712
transform 1 0 2892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1712622712
transform 1 0 2404 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1712622712
transform 1 0 2236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1712622712
transform 1 0 2076 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1712622712
transform 1 0 2020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1712622712
transform 1 0 2668 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1712622712
transform 1 0 2572 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1712622712
transform 1 0 1404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1712622712
transform 1 0 1220 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1712622712
transform 1 0 1172 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1712622712
transform 1 0 1164 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1712622712
transform 1 0 1132 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1712622712
transform 1 0 1556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1712622712
transform 1 0 1532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1712622712
transform 1 0 1220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1712622712
transform 1 0 820 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1712622712
transform 1 0 660 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1712622712
transform 1 0 748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1712622712
transform 1 0 684 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1712622712
transform 1 0 668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1712622712
transform 1 0 508 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1712622712
transform 1 0 476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1712622712
transform 1 0 292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1712622712
transform 1 0 284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1712622712
transform 1 0 228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1712622712
transform 1 0 1052 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1712622712
transform 1 0 892 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1712622712
transform 1 0 844 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1712622712
transform 1 0 780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1712622712
transform 1 0 780 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1712622712
transform 1 0 516 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1712622712
transform 1 0 476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1712622712
transform 1 0 476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1712622712
transform 1 0 452 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1712622712
transform 1 0 444 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1712622712
transform 1 0 436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1712622712
transform 1 0 692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1712622712
transform 1 0 500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1712622712
transform 1 0 388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1712622712
transform 1 0 292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1712622712
transform 1 0 796 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1712622712
transform 1 0 772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1712622712
transform 1 0 444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1712622712
transform 1 0 340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1712622712
transform 1 0 260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1712622712
transform 1 0 2644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1712622712
transform 1 0 2628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1712622712
transform 1 0 2620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1712622712
transform 1 0 2388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1712622712
transform 1 0 2388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1712622712
transform 1 0 3020 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1712622712
transform 1 0 2660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1712622712
transform 1 0 2620 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1712622712
transform 1 0 2396 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1712622712
transform 1 0 2372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1712622712
transform 1 0 2532 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1712622712
transform 1 0 2516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1712622712
transform 1 0 1564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1712622712
transform 1 0 1116 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1712622712
transform 1 0 1116 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1712622712
transform 1 0 1404 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1712622712
transform 1 0 1404 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1712622712
transform 1 0 820 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1712622712
transform 1 0 644 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1712622712
transform 1 0 596 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1712622712
transform 1 0 492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1712622712
transform 1 0 492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1712622712
transform 1 0 380 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1712622712
transform 1 0 260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1712622712
transform 1 0 196 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1712622712
transform 1 0 188 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1712622712
transform 1 0 172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1712622712
transform 1 0 92 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1712622712
transform 1 0 532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1712622712
transform 1 0 476 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1712622712
transform 1 0 476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1712622712
transform 1 0 468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1712622712
transform 1 0 460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1712622712
transform 1 0 412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1712622712
transform 1 0 1300 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1712622712
transform 1 0 572 0 1 1495
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1712622712
transform 1 0 548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1712622712
transform 1 0 460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1712622712
transform 1 0 404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1712622712
transform 1 0 1196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1712622712
transform 1 0 1004 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1712622712
transform 1 0 996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1712622712
transform 1 0 1308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1712622712
transform 1 0 1300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1712622712
transform 1 0 1228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1712622712
transform 1 0 1060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1712622712
transform 1 0 964 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1712622712
transform 1 0 3004 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1712622712
transform 1 0 2964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1712622712
transform 1 0 2756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1712622712
transform 1 0 2236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1712622712
transform 1 0 2076 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1712622712
transform 1 0 2020 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1712622712
transform 1 0 1988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1712622712
transform 1 0 1940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1712622712
transform 1 0 2660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1712622712
transform 1 0 2596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1712622712
transform 1 0 2540 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1712622712
transform 1 0 2420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1712622712
transform 1 0 2372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1712622712
transform 1 0 1884 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1712622712
transform 1 0 1884 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1712622712
transform 1 0 1860 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1712622712
transform 1 0 1812 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1712622712
transform 1 0 1620 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1712622712
transform 1 0 1564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1712622712
transform 1 0 2644 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1712622712
transform 1 0 2636 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1712622712
transform 1 0 2612 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1712622712
transform 1 0 2540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1712622712
transform 1 0 2444 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1712622712
transform 1 0 1372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1712622712
transform 1 0 1764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1712622712
transform 1 0 1372 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1712622712
transform 1 0 1260 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1712622712
transform 1 0 1524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1712622712
transform 1 0 1076 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1712622712
transform 1 0 1068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1712622712
transform 1 0 852 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1712622712
transform 1 0 628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1712622712
transform 1 0 612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1712622712
transform 1 0 580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1712622712
transform 1 0 508 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1712622712
transform 1 0 260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1712622712
transform 1 0 164 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1712622712
transform 1 0 164 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1712622712
transform 1 0 2084 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1712622712
transform 1 0 924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1712622712
transform 1 0 468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1712622712
transform 1 0 444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1712622712
transform 1 0 404 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1712622712
transform 1 0 396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1712622712
transform 1 0 356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1712622712
transform 1 0 524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1712622712
transform 1 0 468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1712622712
transform 1 0 468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1712622712
transform 1 0 340 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1712622712
transform 1 0 332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1712622712
transform 1 0 2620 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1712622712
transform 1 0 2612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1712622712
transform 1 0 2572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1712622712
transform 1 0 2564 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1712622712
transform 1 0 2564 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1712622712
transform 1 0 2332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1712622712
transform 1 0 2300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1712622712
transform 1 0 2268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1712622712
transform 1 0 2260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1712622712
transform 1 0 2468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1712622712
transform 1 0 2428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1712622712
transform 1 0 2388 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1712622712
transform 1 0 1892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1712622712
transform 1 0 1868 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1712622712
transform 1 0 2652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1712622712
transform 1 0 2500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1712622712
transform 1 0 2436 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1712622712
transform 1 0 2412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1712622712
transform 1 0 2404 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1712622712
transform 1 0 2372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1712622712
transform 1 0 2884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1712622712
transform 1 0 2204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1712622712
transform 1 0 1708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1712622712
transform 1 0 1588 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1712622712
transform 1 0 1556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1712622712
transform 1 0 1476 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1712622712
transform 1 0 1108 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1712622712
transform 1 0 964 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1712622712
transform 1 0 900 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1712622712
transform 1 0 868 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1712622712
transform 1 0 676 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1712622712
transform 1 0 556 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1712622712
transform 1 0 604 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1712622712
transform 1 0 548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1712622712
transform 1 0 476 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1712622712
transform 1 0 444 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1712622712
transform 1 0 404 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1712622712
transform 1 0 396 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1712622712
transform 1 0 452 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1712622712
transform 1 0 412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1712622712
transform 1 0 372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1712622712
transform 1 0 348 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1712622712
transform 1 0 260 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1712622712
transform 1 0 212 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1712622712
transform 1 0 148 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1712622712
transform 1 0 228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1712622712
transform 1 0 76 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1712622712
transform 1 0 76 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1712622712
transform 1 0 204 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1712622712
transform 1 0 124 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1712622712
transform 1 0 1156 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1712622712
transform 1 0 1012 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1712622712
transform 1 0 932 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1712622712
transform 1 0 1140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1712622712
transform 1 0 1140 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1712622712
transform 1 0 1204 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1712622712
transform 1 0 1204 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1712622712
transform 1 0 1340 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1712622712
transform 1 0 1324 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1712622712
transform 1 0 1324 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1712622712
transform 1 0 1388 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1712622712
transform 1 0 1348 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1712622712
transform 1 0 1348 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1712622712
transform 1 0 1572 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1712622712
transform 1 0 1564 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1712622712
transform 1 0 1516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1712622712
transform 1 0 1644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1712622712
transform 1 0 1644 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1712622712
transform 1 0 1940 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1712622712
transform 1 0 1860 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1712622712
transform 1 0 1820 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1712622712
transform 1 0 1780 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1712622712
transform 1 0 1780 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1712622712
transform 1 0 1764 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1712622712
transform 1 0 2084 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1712622712
transform 1 0 2068 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1712622712
transform 1 0 2164 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1712622712
transform 1 0 2156 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1712622712
transform 1 0 2140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1712622712
transform 1 0 2348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1712622712
transform 1 0 2324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1712622712
transform 1 0 2316 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1712622712
transform 1 0 2028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1712622712
transform 1 0 2020 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1712622712
transform 1 0 1996 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1712622712
transform 1 0 2412 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1712622712
transform 1 0 2388 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1712622712
transform 1 0 2380 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1712622712
transform 1 0 2708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1712622712
transform 1 0 2708 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1712622712
transform 1 0 2532 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1712622712
transform 1 0 2724 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1712622712
transform 1 0 2700 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1712622712
transform 1 0 2572 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1712622712
transform 1 0 2548 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1712622712
transform 1 0 2540 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1712622712
transform 1 0 2828 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1712622712
transform 1 0 2804 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1712622712
transform 1 0 2772 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1712622712
transform 1 0 2756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1712622712
transform 1 0 3188 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1712622712
transform 1 0 3108 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1712622712
transform 1 0 3068 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1712622712
transform 1 0 2716 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1712622712
transform 1 0 2708 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1712622712
transform 1 0 3100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1712622712
transform 1 0 3100 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1712622712
transform 1 0 3036 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1712622712
transform 1 0 3028 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1712622712
transform 1 0 2988 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1712622712
transform 1 0 2972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1712622712
transform 1 0 2964 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1712622712
transform 1 0 2916 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1712622712
transform 1 0 2900 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1712622712
transform 1 0 2884 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1712622712
transform 1 0 3236 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1712622712
transform 1 0 3236 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1712622712
transform 1 0 3236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1712622712
transform 1 0 3180 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1712622712
transform 1 0 3164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1712622712
transform 1 0 3156 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1712622712
transform 1 0 3404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1712622712
transform 1 0 3324 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1712622712
transform 1 0 3292 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1712622712
transform 1 0 3228 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1712622712
transform 1 0 3140 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1712622712
transform 1 0 3124 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1712622712
transform 1 0 3124 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1712622712
transform 1 0 3036 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1712622712
transform 1 0 3268 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1712622712
transform 1 0 3244 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1712622712
transform 1 0 3092 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1712622712
transform 1 0 3324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1712622712
transform 1 0 3324 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1712622712
transform 1 0 3292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1712622712
transform 1 0 3252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1712622712
transform 1 0 3164 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1712622712
transform 1 0 3204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1712622712
transform 1 0 3172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1712622712
transform 1 0 3420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1712622712
transform 1 0 3380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1712622712
transform 1 0 3292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1712622712
transform 1 0 3260 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1712622712
transform 1 0 3236 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1712622712
transform 1 0 2820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1712622712
transform 1 0 2788 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1712622712
transform 1 0 2972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1712622712
transform 1 0 2948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1712622712
transform 1 0 3220 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1712622712
transform 1 0 3164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1712622712
transform 1 0 3164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1712622712
transform 1 0 3116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1712622712
transform 1 0 3060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1712622712
transform 1 0 3060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1712622712
transform 1 0 3412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1712622712
transform 1 0 3404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1712622712
transform 1 0 3364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1712622712
transform 1 0 3348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1712622712
transform 1 0 3196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1712622712
transform 1 0 3180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1712622712
transform 1 0 3396 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1712622712
transform 1 0 3364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1712622712
transform 1 0 3316 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1712622712
transform 1 0 3212 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1712622712
transform 1 0 3268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1712622712
transform 1 0 3244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1712622712
transform 1 0 3244 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1712622712
transform 1 0 3204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1712622712
transform 1 0 3172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1712622712
transform 1 0 3124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1712622712
transform 1 0 3076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1712622712
transform 1 0 3188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1712622712
transform 1 0 3172 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1712622712
transform 1 0 3084 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1712622712
transform 1 0 2644 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1712622712
transform 1 0 1716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1712622712
transform 1 0 3356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1712622712
transform 1 0 3300 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1712622712
transform 1 0 3292 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1712622712
transform 1 0 3172 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1712622712
transform 1 0 3164 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1712622712
transform 1 0 3132 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1712622712
transform 1 0 3132 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1712622712
transform 1 0 2148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1712622712
transform 1 0 2092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1712622712
transform 1 0 2124 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1712622712
transform 1 0 1972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1712622712
transform 1 0 2060 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1712622712
transform 1 0 2060 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1712622712
transform 1 0 1964 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1712622712
transform 1 0 1964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1712622712
transform 1 0 1948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1712622712
transform 1 0 2140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1712622712
transform 1 0 1972 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1712622712
transform 1 0 1956 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1712622712
transform 1 0 1900 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1712622712
transform 1 0 1860 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1712622712
transform 1 0 1860 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1712622712
transform 1 0 1924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1712622712
transform 1 0 1924 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1712622712
transform 1 0 2276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1712622712
transform 1 0 2132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1712622712
transform 1 0 2132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1712622712
transform 1 0 2220 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1712622712
transform 1 0 2220 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1712622712
transform 1 0 2220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1712622712
transform 1 0 2188 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1712622712
transform 1 0 2156 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1712622712
transform 1 0 2420 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1712622712
transform 1 0 2412 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1712622712
transform 1 0 2524 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1712622712
transform 1 0 2508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1712622712
transform 1 0 2532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1712622712
transform 1 0 2412 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1712622712
transform 1 0 2380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1712622712
transform 1 0 2500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1712622712
transform 1 0 2460 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1712622712
transform 1 0 2380 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1712622712
transform 1 0 2380 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1712622712
transform 1 0 2348 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1712622712
transform 1 0 2340 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1712622712
transform 1 0 2580 0 1 1695
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1712622712
transform 1 0 2564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1712622712
transform 1 0 2044 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1712622712
transform 1 0 2044 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1712622712
transform 1 0 2020 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1712622712
transform 1 0 1996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1712622712
transform 1 0 1660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1712622712
transform 1 0 1636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1712622712
transform 1 0 2668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1712622712
transform 1 0 2628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1712622712
transform 1 0 2580 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1712622712
transform 1 0 1420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1712622712
transform 1 0 1348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1712622712
transform 1 0 1348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1712622712
transform 1 0 1316 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1712622712
transform 1 0 1284 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1712622712
transform 1 0 1244 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1712622712
transform 1 0 900 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1712622712
transform 1 0 1636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1712622712
transform 1 0 1588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1712622712
transform 1 0 1172 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1712622712
transform 1 0 1116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1712622712
transform 1 0 1052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1712622712
transform 1 0 1004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1712622712
transform 1 0 996 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1712622712
transform 1 0 1452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1712622712
transform 1 0 1420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1712622712
transform 1 0 1020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1712622712
transform 1 0 1020 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1712622712
transform 1 0 1700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1712622712
transform 1 0 1684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1712622712
transform 1 0 1124 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1712622712
transform 1 0 1116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1712622712
transform 1 0 1092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1712622712
transform 1 0 1084 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1712622712
transform 1 0 1476 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1712622712
transform 1 0 1444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1712622712
transform 1 0 1748 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1712622712
transform 1 0 1716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1712622712
transform 1 0 1212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1712622712
transform 1 0 1172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1712622712
transform 1 0 684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1712622712
transform 1 0 604 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1712622712
transform 1 0 516 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1712622712
transform 1 0 1196 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1712622712
transform 1 0 1108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1712622712
transform 1 0 804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1712622712
transform 1 0 748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1712622712
transform 1 0 804 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1712622712
transform 1 0 604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1712622712
transform 1 0 892 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1712622712
transform 1 0 556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1712622712
transform 1 0 284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1712622712
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1712622712
transform 1 0 812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1712622712
transform 1 0 812 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1712622712
transform 1 0 236 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1712622712
transform 1 0 204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1712622712
transform 1 0 316 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1712622712
transform 1 0 316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1712622712
transform 1 0 204 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1712622712
transform 1 0 204 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1712622712
transform 1 0 172 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1712622712
transform 1 0 172 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1712622712
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1712622712
transform 1 0 708 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1712622712
transform 1 0 516 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1712622712
transform 1 0 508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1712622712
transform 1 0 444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1712622712
transform 1 0 404 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1712622712
transform 1 0 252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1712622712
transform 1 0 116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1712622712
transform 1 0 116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1712622712
transform 1 0 300 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1712622712
transform 1 0 276 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1712622712
transform 1 0 172 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1712622712
transform 1 0 140 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1712622712
transform 1 0 420 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1712622712
transform 1 0 388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1712622712
transform 1 0 124 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1712622712
transform 1 0 68 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1712622712
transform 1 0 660 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1712622712
transform 1 0 644 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1712622712
transform 1 0 116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1712622712
transform 1 0 68 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1712622712
transform 1 0 252 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1712622712
transform 1 0 228 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1712622712
transform 1 0 212 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1712622712
transform 1 0 180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1712622712
transform 1 0 732 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1712622712
transform 1 0 716 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1712622712
transform 1 0 1868 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1712622712
transform 1 0 1692 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1712622712
transform 1 0 1652 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1712622712
transform 1 0 900 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1712622712
transform 1 0 892 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1712622712
transform 1 0 860 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1712622712
transform 1 0 820 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1712622712
transform 1 0 772 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1712622712
transform 1 0 708 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1712622712
transform 1 0 708 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1712622712
transform 1 0 684 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1712622712
transform 1 0 772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1712622712
transform 1 0 732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1712622712
transform 1 0 564 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1712622712
transform 1 0 564 0 1 1045
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1712622712
transform 1 0 460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1712622712
transform 1 0 444 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1712622712
transform 1 0 596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1712622712
transform 1 0 564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1712622712
transform 1 0 924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1712622712
transform 1 0 900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1712622712
transform 1 0 836 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1712622712
transform 1 0 788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1712622712
transform 1 0 988 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1712622712
transform 1 0 500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1712622712
transform 1 0 828 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1712622712
transform 1 0 804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1712622712
transform 1 0 804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1712622712
transform 1 0 1196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1712622712
transform 1 0 1180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1712622712
transform 1 0 1252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1712622712
transform 1 0 1188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1712622712
transform 1 0 1404 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1712622712
transform 1 0 1132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1712622712
transform 1 0 1132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1712622712
transform 1 0 1508 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1712622712
transform 1 0 1380 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1712622712
transform 1 0 1708 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1712622712
transform 1 0 1580 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1712622712
transform 1 0 1340 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1712622712
transform 1 0 1028 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1712622712
transform 1 0 1556 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1712622712
transform 1 0 1268 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1712622712
transform 1 0 1156 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1712622712
transform 1 0 1068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1712622712
transform 1 0 1068 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1712622712
transform 1 0 1004 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1712622712
transform 1 0 1588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1712622712
transform 1 0 1260 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1712622712
transform 1 0 1316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1712622712
transform 1 0 1284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1712622712
transform 1 0 1540 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1712622712
transform 1 0 1500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1712622712
transform 1 0 1412 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1712622712
transform 1 0 1380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1712622712
transform 1 0 1380 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1712622712
transform 1 0 1364 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1712622712
transform 1 0 1796 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1712622712
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1712622712
transform 1 0 1660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1712622712
transform 1 0 1644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1712622712
transform 1 0 1684 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1712622712
transform 1 0 1684 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1712622712
transform 1 0 1676 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1712622712
transform 1 0 1652 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1712622712
transform 1 0 1636 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1712622712
transform 1 0 1948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1712622712
transform 1 0 1884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1712622712
transform 1 0 1892 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1712622712
transform 1 0 1876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1712622712
transform 1 0 1772 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1712622712
transform 1 0 1764 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1712622712
transform 1 0 2076 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1712622712
transform 1 0 2060 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1712622712
transform 1 0 2164 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1712622712
transform 1 0 2124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1712622712
transform 1 0 2188 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1712622712
transform 1 0 2172 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1712622712
transform 1 0 2044 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1712622712
transform 1 0 1852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1712622712
transform 1 0 1820 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1712622712
transform 1 0 2044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1712622712
transform 1 0 2044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1712622712
transform 1 0 1612 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1712622712
transform 1 0 1588 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1712622712
transform 1 0 1548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1712622712
transform 1 0 1516 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1712622712
transform 1 0 1756 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1712622712
transform 1 0 1732 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1712622712
transform 1 0 1692 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1712622712
transform 1 0 1684 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1712622712
transform 1 0 2724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1712622712
transform 1 0 2708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1712622712
transform 1 0 1892 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1712622712
transform 1 0 1844 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1712622712
transform 1 0 1836 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1712622712
transform 1 0 1772 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1712622712
transform 1 0 1684 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1712622712
transform 1 0 2028 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1712622712
transform 1 0 1828 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1712622712
transform 1 0 1748 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1712622712
transform 1 0 1740 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1712622712
transform 1 0 980 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1712622712
transform 1 0 948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1712622712
transform 1 0 2604 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1712622712
transform 1 0 2412 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1712622712
transform 1 0 2396 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1712622712
transform 1 0 2212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1712622712
transform 1 0 2180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1712622712
transform 1 0 2428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1712622712
transform 1 0 2412 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1712622712
transform 1 0 2140 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1712622712
transform 1 0 2084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1712622712
transform 1 0 2060 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1712622712
transform 1 0 2852 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1712622712
transform 1 0 2516 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1712622712
transform 1 0 2460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1712622712
transform 1 0 2268 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1712622712
transform 1 0 2180 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1712622712
transform 1 0 2020 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1712622712
transform 1 0 2844 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1712622712
transform 1 0 2636 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1712622712
transform 1 0 2292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1712622712
transform 1 0 2564 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1712622712
transform 1 0 2476 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1712622712
transform 1 0 2468 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1712622712
transform 1 0 2812 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1712622712
transform 1 0 2812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1712622712
transform 1 0 3412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1712622712
transform 1 0 3340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1712622712
transform 1 0 3300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1712622712
transform 1 0 3412 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1712622712
transform 1 0 3356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1712622712
transform 1 0 3316 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1712622712
transform 1 0 3252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1712622712
transform 1 0 3252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1712622712
transform 1 0 3340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1712622712
transform 1 0 3316 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1712622712
transform 1 0 3292 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1712622712
transform 1 0 3252 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1712622712
transform 1 0 3388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1712622712
transform 1 0 3388 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1712622712
transform 1 0 3412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1712622712
transform 1 0 3356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1712622712
transform 1 0 3324 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1712622712
transform 1 0 3300 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1712622712
transform 1 0 3260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1712622712
transform 1 0 2964 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1712622712
transform 1 0 2964 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1712622712
transform 1 0 2948 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1712622712
transform 1 0 2900 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1712622712
transform 1 0 2692 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1712622712
transform 1 0 2692 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1712622712
transform 1 0 3356 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1712622712
transform 1 0 3284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1712622712
transform 1 0 3268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1712622712
transform 1 0 3252 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1712622712
transform 1 0 3188 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1712622712
transform 1 0 3148 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1712622712
transform 1 0 3132 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1712622712
transform 1 0 2852 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1712622712
transform 1 0 2780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1712622712
transform 1 0 2780 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1712622712
transform 1 0 2340 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1712622712
transform 1 0 1452 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1712622712
transform 1 0 1284 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1712622712
transform 1 0 836 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1712622712
transform 1 0 3236 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1712622712
transform 1 0 3196 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1712622712
transform 1 0 3180 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1712622712
transform 1 0 3228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1712622712
transform 1 0 3228 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1712622712
transform 1 0 3204 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1712622712
transform 1 0 3204 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1712622712
transform 1 0 3348 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1712622712
transform 1 0 3308 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1712622712
transform 1 0 3284 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1712622712
transform 1 0 2428 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1712622712
transform 1 0 2252 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1712622712
transform 1 0 2156 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1712622712
transform 1 0 2068 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1712622712
transform 1 0 1988 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1712622712
transform 1 0 1844 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1712622712
transform 1 0 1692 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1712622712
transform 1 0 1532 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1712622712
transform 1 0 1484 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1712622712
transform 1 0 1388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1712622712
transform 1 0 1364 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1712622712
transform 1 0 1212 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1712622712
transform 1 0 1028 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1712622712
transform 1 0 3212 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1712622712
transform 1 0 3212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1712622712
transform 1 0 3068 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1712622712
transform 1 0 3060 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1712622712
transform 1 0 1068 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1712622712
transform 1 0 964 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1712622712
transform 1 0 780 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1712622712
transform 1 0 476 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1712622712
transform 1 0 436 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1712622712
transform 1 0 316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1712622712
transform 1 0 276 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1712622712
transform 1 0 260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1712622712
transform 1 0 212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1712622712
transform 1 0 148 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1712622712
transform 1 0 92 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1712622712
transform 1 0 92 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1712622712
transform 1 0 3348 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1712622712
transform 1 0 3340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1712622712
transform 1 0 3340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1712622712
transform 1 0 3324 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1712622712
transform 1 0 3220 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1712622712
transform 1 0 3196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1712622712
transform 1 0 3164 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1712622712
transform 1 0 3156 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1712622712
transform 1 0 3108 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1712622712
transform 1 0 3108 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1712622712
transform 1 0 3060 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1712622712
transform 1 0 3052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1712622712
transform 1 0 2980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1712622712
transform 1 0 2932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1712622712
transform 1 0 2812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1712622712
transform 1 0 2788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1712622712
transform 1 0 2756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1712622712
transform 1 0 2740 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1712622712
transform 1 0 3348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1712622712
transform 1 0 3340 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1712622712
transform 1 0 3244 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1712622712
transform 1 0 3244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1712622712
transform 1 0 3172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1712622712
transform 1 0 2956 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1712622712
transform 1 0 2892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1712622712
transform 1 0 2764 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1712622712
transform 1 0 2652 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1712622712
transform 1 0 2580 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1712622712
transform 1 0 2532 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1712622712
transform 1 0 2468 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1712622712
transform 1 0 2356 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1712622712
transform 1 0 2356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1712622712
transform 1 0 2220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1712622712
transform 1 0 2156 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1712622712
transform 1 0 2156 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1712622712
transform 1 0 2036 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1712622712
transform 1 0 1916 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1712622712
transform 1 0 1908 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1712622712
transform 1 0 1804 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1712622712
transform 1 0 1692 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1712622712
transform 1 0 1580 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1712622712
transform 1 0 1428 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1712622712
transform 1 0 1332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1712622712
transform 1 0 1220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1712622712
transform 1 0 1004 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1712622712
transform 1 0 900 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1712622712
transform 1 0 3004 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1712622712
transform 1 0 2908 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1712622712
transform 1 0 2316 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1712622712
transform 1 0 1116 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1712622712
transform 1 0 796 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1712622712
transform 1 0 684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1712622712
transform 1 0 580 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1712622712
transform 1 0 380 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1712622712
transform 1 0 364 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1712622712
transform 1 0 316 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1712622712
transform 1 0 244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1712622712
transform 1 0 204 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1712622712
transform 1 0 124 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1712622712
transform 1 0 92 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1712622712
transform 1 0 2972 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1712622712
transform 1 0 2868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1712622712
transform 1 0 2772 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1712622712
transform 1 0 2676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1712622712
transform 1 0 2572 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1712622712
transform 1 0 2476 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1712622712
transform 1 0 2380 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1712622712
transform 1 0 2276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1712622712
transform 1 0 2180 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1712622712
transform 1 0 2084 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1712622712
transform 1 0 1980 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1712622712
transform 1 0 1908 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1712622712
transform 1 0 1884 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1712622712
transform 1 0 1780 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1712622712
transform 1 0 1756 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1712622712
transform 1 0 1644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1712622712
transform 1 0 1532 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1712622712
transform 1 0 1476 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1712622712
transform 1 0 1372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1712622712
transform 1 0 1268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1712622712
transform 1 0 1036 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1712622712
transform 1 0 980 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1712622712
transform 1 0 540 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1712622712
transform 1 0 212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1712622712
transform 1 0 204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1712622712
transform 1 0 140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1712622712
transform 1 0 100 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1712622712
transform 1 0 92 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1712622712
transform 1 0 3348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1712622712
transform 1 0 3340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1712622712
transform 1 0 3236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1712622712
transform 1 0 3124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1712622712
transform 1 0 3116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1712622712
transform 1 0 2956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1712622712
transform 1 0 2748 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1712622712
transform 1 0 1756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1712622712
transform 1 0 1164 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1712622712
transform 1 0 868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1712622712
transform 1 0 756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1712622712
transform 1 0 644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1712622712
transform 1 0 428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1712622712
transform 1 0 316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1712622712
transform 1 0 2324 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1712622712
transform 1 0 2300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1712622712
transform 1 0 2140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1712622712
transform 1 0 1932 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1712622712
transform 1 0 1892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1712622712
transform 1 0 1740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1712622712
transform 1 0 1724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1712622712
transform 1 0 2452 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1712622712
transform 1 0 2444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1712622712
transform 1 0 2412 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1712622712
transform 1 0 2388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1712622712
transform 1 0 2276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1712622712
transform 1 0 2116 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1712622712
transform 1 0 2628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1712622712
transform 1 0 2468 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1712622712
transform 1 0 2292 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1712622712
transform 1 0 2268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1712622712
transform 1 0 2132 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1712622712
transform 1 0 1996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1712622712
transform 1 0 1844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1712622712
transform 1 0 1764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1712622712
transform 1 0 1668 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1712622712
transform 1 0 1564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1712622712
transform 1 0 1476 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1712622712
transform 1 0 1452 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1712622712
transform 1 0 2852 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1712622712
transform 1 0 2292 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1712622712
transform 1 0 1212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1712622712
transform 1 0 916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1712622712
transform 1 0 748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1712622712
transform 1 0 188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1712622712
transform 1 0 132 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1712622712
transform 1 0 100 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1712622712
transform 1 0 2836 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1712622712
transform 1 0 2428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1712622712
transform 1 0 724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1712622712
transform 1 0 628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1712622712
transform 1 0 508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1712622712
transform 1 0 372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1712622712
transform 1 0 308 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1712622712
transform 1 0 308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1712622712
transform 1 0 2756 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1712622712
transform 1 0 2404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1712622712
transform 1 0 1124 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1712622712
transform 1 0 884 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1712622712
transform 1 0 2604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1712622712
transform 1 0 2476 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1712622712
transform 1 0 2468 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1712622712
transform 1 0 2396 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1712622712
transform 1 0 2284 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1712622712
transform 1 0 2172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1712622712
transform 1 0 2148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1712622712
transform 1 0 1972 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1712622712
transform 1 0 2852 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1712622712
transform 1 0 2772 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1712622712
transform 1 0 2484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1712622712
transform 1 0 1172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1712622712
transform 1 0 900 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1712622712
transform 1 0 740 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1712622712
transform 1 0 644 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1712622712
transform 1 0 524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1712622712
transform 1 0 436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1712622712
transform 1 0 356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1712622712
transform 1 0 356 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1712622712
transform 1 0 324 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1712622712
transform 1 0 260 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1712622712
transform 1 0 180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1712622712
transform 1 0 116 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1712622712
transform 1 0 2980 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1712622712
transform 1 0 2964 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1712622712
transform 1 0 3044 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1712622712
transform 1 0 2996 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1712622712
transform 1 0 2924 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1712622712
transform 1 0 3084 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1712622712
transform 1 0 2972 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1712622712
transform 1 0 2724 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1712622712
transform 1 0 2572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1712622712
transform 1 0 2556 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1712622712
transform 1 0 2036 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1712622712
transform 1 0 1844 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1712622712
transform 1 0 1668 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1712622712
transform 1 0 1580 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1712622712
transform 1 0 1364 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1712622712
transform 1 0 1340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1712622712
transform 1 0 1324 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1712622712
transform 1 0 1156 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1712622712
transform 1 0 948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1712622712
transform 1 0 364 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1712622712
transform 1 0 164 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1712622712
transform 1 0 140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1712622712
transform 1 0 124 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1712622712
transform 1 0 3020 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1712622712
transform 1 0 2932 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1712622712
transform 1 0 2828 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1712622712
transform 1 0 2492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1712622712
transform 1 0 2484 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1712622712
transform 1 0 2556 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1712622712
transform 1 0 2524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1712622712
transform 1 0 2308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1712622712
transform 1 0 2236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1712622712
transform 1 0 2148 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1712622712
transform 1 0 2028 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1712622712
transform 1 0 1956 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1712622712
transform 1 0 1828 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1712622712
transform 1 0 1732 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1712622712
transform 1 0 1652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1712622712
transform 1 0 1484 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1712622712
transform 1 0 1372 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1712622712
transform 1 0 1276 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1712622712
transform 1 0 1212 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1712622712
transform 1 0 1156 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1712622712
transform 1 0 988 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1712622712
transform 1 0 988 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1712622712
transform 1 0 868 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1712622712
transform 1 0 684 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1712622712
transform 1 0 676 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1712622712
transform 1 0 620 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1712622712
transform 1 0 572 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1712622712
transform 1 0 548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1712622712
transform 1 0 516 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1712622712
transform 1 0 516 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1712622712
transform 1 0 484 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1712622712
transform 1 0 2860 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1712622712
transform 1 0 2860 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1712622712
transform 1 0 2828 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1712622712
transform 1 0 2812 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1712622712
transform 1 0 3036 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1712622712
transform 1 0 2884 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1712622712
transform 1 0 2788 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1712622712
transform 1 0 2748 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1712622712
transform 1 0 2708 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1712622712
transform 1 0 2532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1712622712
transform 1 0 2396 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1712622712
transform 1 0 2316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1712622712
transform 1 0 2180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1712622712
transform 1 0 2092 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1712622712
transform 1 0 1988 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1712622712
transform 1 0 1932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1712622712
transform 1 0 1788 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1712622712
transform 1 0 1620 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1712622712
transform 1 0 1572 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1712622712
transform 1 0 1396 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1712622712
transform 1 0 1300 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1712622712
transform 1 0 1188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1712622712
transform 1 0 1156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1712622712
transform 1 0 1148 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1712622712
transform 1 0 2364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1712622712
transform 1 0 2276 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1712622712
transform 1 0 2196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1712622712
transform 1 0 2196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1712622712
transform 1 0 2140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1712622712
transform 1 0 2132 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1712622712
transform 1 0 2100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1712622712
transform 1 0 2044 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1712622712
transform 1 0 1860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1712622712
transform 1 0 1780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1712622712
transform 1 0 1756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1712622712
transform 1 0 1716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1712622712
transform 1 0 1684 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1712622712
transform 1 0 1492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1712622712
transform 1 0 1012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1712622712
transform 1 0 796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1712622712
transform 1 0 684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1712622712
transform 1 0 644 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1712622712
transform 1 0 604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1712622712
transform 1 0 508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1712622712
transform 1 0 236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1712622712
transform 1 0 108 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1712622712
transform 1 0 100 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1712622712
transform 1 0 100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1712622712
transform 1 0 92 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1712622712
transform 1 0 92 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1712622712
transform 1 0 68 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1712622712
transform 1 0 68 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1712622712
transform 1 0 68 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1712622712
transform 1 0 2220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1712622712
transform 1 0 1716 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1712622712
transform 1 0 1716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1712622712
transform 1 0 1436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1712622712
transform 1 0 572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1712622712
transform 1 0 412 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1712622712
transform 1 0 356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1712622712
transform 1 0 316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1712622712
transform 1 0 300 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1712622712
transform 1 0 299 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1712622712
transform 1 0 292 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1712622712
transform 1 0 276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1712622712
transform 1 0 276 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1712622712
transform 1 0 260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1712622712
transform 1 0 252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1712622712
transform 1 0 252 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1712622712
transform 1 0 252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1712622712
transform 1 0 2396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1712622712
transform 1 0 2364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1712622712
transform 1 0 2356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1712622712
transform 1 0 2356 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1712622712
transform 1 0 2268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1712622712
transform 1 0 2204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1712622712
transform 1 0 1948 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1712622712
transform 1 0 1836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1712622712
transform 1 0 1772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1712622712
transform 1 0 1604 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1712622712
transform 1 0 1492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1712622712
transform 1 0 1116 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1712622712
transform 1 0 900 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1712622712
transform 1 0 2148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1712622712
transform 1 0 2068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1712622712
transform 1 0 1964 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1712622712
transform 1 0 1948 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1712622712
transform 1 0 1316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1712622712
transform 1 0 604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1712622712
transform 1 0 540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1712622712
transform 1 0 300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1712622712
transform 1 0 172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1712622712
transform 1 0 164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1712622712
transform 1 0 148 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1712622712
transform 1 0 132 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1712622712
transform 1 0 132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1712622712
transform 1 0 132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1712622712
transform 1 0 124 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1712622712
transform 1 0 2308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1712622712
transform 1 0 2228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1712622712
transform 1 0 2228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1712622712
transform 1 0 2220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1712622712
transform 1 0 2172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1712622712
transform 1 0 2164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1712622712
transform 1 0 1924 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1712622712
transform 1 0 1908 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1712622712
transform 1 0 1836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1712622712
transform 1 0 1748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1712622712
transform 1 0 1692 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1712622712
transform 1 0 1532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1712622712
transform 1 0 1060 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1712622712
transform 1 0 868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1712622712
transform 1 0 2740 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1712622712
transform 1 0 2708 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1712622712
transform 1 0 3012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1712622712
transform 1 0 2972 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1712622712
transform 1 0 2956 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1712622712
transform 1 0 2852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1712622712
transform 1 0 2636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1712622712
transform 1 0 2556 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1712622712
transform 1 0 1764 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1712622712
transform 1 0 1412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1712622712
transform 1 0 1164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1712622712
transform 1 0 1148 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1712622712
transform 1 0 2564 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1712622712
transform 1 0 2492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1712622712
transform 1 0 2484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1712622712
transform 1 0 2476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1712622712
transform 1 0 2476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1712622712
transform 1 0 2348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1712622712
transform 1 0 2340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1712622712
transform 1 0 2044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1712622712
transform 1 0 1948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1712622712
transform 1 0 1844 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1712622712
transform 1 0 1732 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1712622712
transform 1 0 1556 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1712622712
transform 1 0 1492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1712622712
transform 1 0 1164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1712622712
transform 1 0 1036 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1712622712
transform 1 0 996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1712622712
transform 1 0 948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1712622712
transform 1 0 836 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1712622712
transform 1 0 836 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1712622712
transform 1 0 804 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1712622712
transform 1 0 724 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1712622712
transform 1 0 692 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1712622712
transform 1 0 604 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1712622712
transform 1 0 604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1712622712
transform 1 0 596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1712622712
transform 1 0 588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1712622712
transform 1 0 580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1712622712
transform 1 0 564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1712622712
transform 1 0 548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1712622712
transform 1 0 3164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1712622712
transform 1 0 2844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1712622712
transform 1 0 2828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1712622712
transform 1 0 3140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1712622712
transform 1 0 3132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1712622712
transform 1 0 3092 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1712622712
transform 1 0 3060 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1712622712
transform 1 0 2892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1712622712
transform 1 0 2588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1712622712
transform 1 0 3228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1712622712
transform 1 0 3140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1712622712
transform 1 0 2836 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1712622712
transform 1 0 2804 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1712622712
transform 1 0 2540 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1712622712
transform 1 0 2452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1712622712
transform 1 0 2444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1712622712
transform 1 0 2444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1712622712
transform 1 0 2436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1712622712
transform 1 0 2308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1712622712
transform 1 0 2300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1712622712
transform 1 0 1916 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1712622712
transform 1 0 1772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1712622712
transform 1 0 1700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1712622712
transform 1 0 1452 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1712622712
transform 1 0 1108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1712622712
transform 1 0 940 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1712622712
transform 1 0 764 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1712622712
transform 1 0 668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1712622712
transform 1 0 660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1712622712
transform 1 0 2828 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1712622712
transform 1 0 2740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1712622712
transform 1 0 2596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1712622712
transform 1 0 2012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1712622712
transform 1 0 1460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1712622712
transform 1 0 1428 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1712622712
transform 1 0 1236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1712622712
transform 1 0 1220 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1712622712
transform 1 0 1212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1712622712
transform 1 0 956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1712622712
transform 1 0 916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1712622712
transform 1 0 564 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1712622712
transform 1 0 548 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1712622712
transform 1 0 532 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1712622712
transform 1 0 532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1712622712
transform 1 0 524 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1712622712
transform 1 0 524 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1712622712
transform 1 0 516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1712622712
transform 1 0 508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1712622712
transform 1 0 508 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1712622712
transform 1 0 2740 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1712622712
transform 1 0 2484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1712622712
transform 1 0 3148 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1712622712
transform 1 0 3076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1712622712
transform 1 0 3004 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1712622712
transform 1 0 2988 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1712622712
transform 1 0 2476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1712622712
transform 1 0 2332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1712622712
transform 1 0 2316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1712622712
transform 1 0 2308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1712622712
transform 1 0 2284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1712622712
transform 1 0 2284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1712622712
transform 1 0 2228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1712622712
transform 1 0 2196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1712622712
transform 1 0 2172 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1712622712
transform 1 0 2172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1712622712
transform 1 0 2156 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1712622712
transform 1 0 1876 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1712622712
transform 1 0 1788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1712622712
transform 1 0 1708 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1712622712
transform 1 0 1452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1712622712
transform 1 0 1084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1712622712
transform 1 0 836 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1712622712
transform 1 0 356 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1712622712
transform 1 0 324 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1712622712
transform 1 0 228 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1712622712
transform 1 0 2668 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1712622712
transform 1 0 2556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1712622712
transform 1 0 2172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1712622712
transform 1 0 1500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1712622712
transform 1 0 1428 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1712622712
transform 1 0 1396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1712622712
transform 1 0 1172 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1712622712
transform 1 0 1172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1712622712
transform 1 0 852 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1712622712
transform 1 0 844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1712622712
transform 1 0 628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1712622712
transform 1 0 268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1712622712
transform 1 0 244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1712622712
transform 1 0 244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1712622712
transform 1 0 212 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1712622712
transform 1 0 204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1712622712
transform 1 0 188 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1712622712
transform 1 0 188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1712622712
transform 1 0 2868 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1712622712
transform 1 0 2812 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1712622712
transform 1 0 2588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1712622712
transform 1 0 1636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1712622712
transform 1 0 1524 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1712622712
transform 1 0 1356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1712622712
transform 1 0 1340 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1712622712
transform 1 0 2596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1712622712
transform 1 0 2596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1712622712
transform 1 0 2580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1712622712
transform 1 0 2556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1712622712
transform 1 0 2412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1712622712
transform 1 0 2372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1712622712
transform 1 0 2180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1712622712
transform 1 0 2124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1712622712
transform 1 0 2012 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1712622712
transform 1 0 1948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1712622712
transform 1 0 1884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1712622712
transform 1 0 1780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1712622712
transform 1 0 1436 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1712622712
transform 1 0 1332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1712622712
transform 1 0 1220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1712622712
transform 1 0 956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1712622712
transform 1 0 812 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1712622712
transform 1 0 756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1712622712
transform 1 0 756 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1712622712
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1712622712
transform 1 0 516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1712622712
transform 1 0 500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1712622712
transform 1 0 492 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1712622712
transform 1 0 484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1712622712
transform 1 0 476 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1712622712
transform 1 0 460 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1712622712
transform 1 0 460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1712622712
transform 1 0 412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1712622712
transform 1 0 412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1712622712
transform 1 0 380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1712622712
transform 1 0 3188 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1712622712
transform 1 0 3140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1712622712
transform 1 0 3020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1712622712
transform 1 0 3012 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1712622712
transform 1 0 3308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1712622712
transform 1 0 3268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1712622712
transform 1 0 3236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1712622712
transform 1 0 2804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1712622712
transform 1 0 3076 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1712622712
transform 1 0 3004 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1712622712
transform 1 0 2932 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1712622712
transform 1 0 2884 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1712622712
transform 1 0 2788 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1712622712
transform 1 0 2572 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1712622712
transform 1 0 2452 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1712622712
transform 1 0 2356 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1712622712
transform 1 0 2348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1712622712
transform 1 0 2300 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1712622712
transform 1 0 2252 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1712622712
transform 1 0 2204 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1712622712
transform 1 0 2132 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1712622712
transform 1 0 2116 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1712622712
transform 1 0 2004 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1712622712
transform 1 0 1900 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1712622712
transform 1 0 1772 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1712622712
transform 1 0 1756 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1712622712
transform 1 0 1556 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1712622712
transform 1 0 1524 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1712622712
transform 1 0 1284 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1712622712
transform 1 0 1156 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1712622712
transform 1 0 1116 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1712622712
transform 1 0 868 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1712622712
transform 1 0 844 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1712622712
transform 1 0 692 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1712622712
transform 1 0 612 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1712622712
transform 1 0 420 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1712622712
transform 1 0 324 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1712622712
transform 1 0 292 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1712622712
transform 1 0 244 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1712622712
transform 1 0 236 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1712622712
transform 1 0 228 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1712622712
transform 1 0 188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1712622712
transform 1 0 164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1712622712
transform 1 0 164 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1712622712
transform 1 0 148 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1712622712
transform 1 0 2732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1712622712
transform 1 0 2716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1712622712
transform 1 0 2700 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1712622712
transform 1 0 2684 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1712622712
transform 1 0 2668 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1712622712
transform 1 0 2644 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1712622712
transform 1 0 2596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1712622712
transform 1 0 2572 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1712622712
transform 1 0 2540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1712622712
transform 1 0 2052 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1712622712
transform 1 0 1892 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1712622712
transform 1 0 1588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1712622712
transform 1 0 1260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1712622712
transform 1 0 1204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1712622712
transform 1 0 1204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1712622712
transform 1 0 1180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1712622712
transform 1 0 1164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1712622712
transform 1 0 1164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1712622712
transform 1 0 1116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1712622712
transform 1 0 2700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1712622712
transform 1 0 2580 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1712622712
transform 1 0 2540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1712622712
transform 1 0 2316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1712622712
transform 1 0 2148 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1712622712
transform 1 0 2028 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1712622712
transform 1 0 2028 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1712622712
transform 1 0 2004 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1712622712
transform 1 0 2004 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1712622712
transform 1 0 1836 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1712622712
transform 1 0 1652 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1712622712
transform 1 0 1644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1712622712
transform 1 0 1564 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1712622712
transform 1 0 1236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1712622712
transform 1 0 1180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1712622712
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1712622712
transform 1 0 1132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1712622712
transform 1 0 1124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1712622712
transform 1 0 1092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1712622712
transform 1 0 3324 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1712622712
transform 1 0 3268 0 1 655
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1712622712
transform 1 0 3268 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1712622712
transform 1 0 3228 0 1 655
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1712622712
transform 1 0 3204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1712622712
transform 1 0 1732 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1712622712
transform 1 0 1068 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1712622712
transform 1 0 932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1712622712
transform 1 0 884 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1712622712
transform 1 0 692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1712622712
transform 1 0 628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1712622712
transform 1 0 508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1712622712
transform 1 0 428 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1712622712
transform 1 0 356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1712622712
transform 1 0 308 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1712622712
transform 1 0 260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1712622712
transform 1 0 188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1712622712
transform 1 0 140 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1712622712
transform 1 0 84 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1712622712
transform 1 0 2868 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1712622712
transform 1 0 2676 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1712622712
transform 1 0 2332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1712622712
transform 1 0 2268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1712622712
transform 1 0 2236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1712622712
transform 1 0 2084 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1712622712
transform 1 0 2044 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1712622712
transform 1 0 1884 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1712622712
transform 1 0 1828 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1712622712
transform 1 0 1772 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1712622712
transform 1 0 1660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1712622712
transform 1 0 1444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1712622712
transform 1 0 1372 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1712622712
transform 1 0 1292 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1712622712
transform 1 0 3340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1712622712
transform 1 0 3284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1712622712
transform 1 0 3220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1712622712
transform 1 0 3172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1712622712
transform 1 0 3108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1712622712
transform 1 0 3108 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1712622712
transform 1 0 2996 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1712622712
transform 1 0 2956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1712622712
transform 1 0 2804 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1712622712
transform 1 0 2780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1712622712
transform 1 0 2684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1712622712
transform 1 0 2604 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1712622712
transform 1 0 2452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1712622712
transform 1 0 1340 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1712622712
transform 1 0 1780 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1712622712
transform 1 0 1468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1712622712
transform 1 0 1244 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1712622712
transform 1 0 1180 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1712622712
transform 1 0 1100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1712622712
transform 1 0 924 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1712622712
transform 1 0 636 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1712622712
transform 1 0 612 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1712622712
transform 1 0 588 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1712622712
transform 1 0 524 0 1 3095
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1712622712
transform 1 0 492 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1712622712
transform 1 0 484 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1712622712
transform 1 0 436 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1712622712
transform 1 0 428 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1712622712
transform 1 0 2524 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1712622712
transform 1 0 2516 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1712622712
transform 1 0 2484 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1712622712
transform 1 0 2444 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1712622712
transform 1 0 2252 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1712622712
transform 1 0 2196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1712622712
transform 1 0 2116 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1712622712
transform 1 0 1988 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1712622712
transform 1 0 1924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1712622712
transform 1 0 1668 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1712622712
transform 1 0 1620 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1712622712
transform 1 0 1444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1712622712
transform 1 0 1324 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1712622712
transform 1 0 1324 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1712622712
transform 1 0 956 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1712622712
transform 1 0 3340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1712622712
transform 1 0 3332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1712622712
transform 1 0 3308 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1712622712
transform 1 0 3292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1712622712
transform 1 0 3252 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1712622712
transform 1 0 3220 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1712622712
transform 1 0 3196 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1712622712
transform 1 0 3188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1712622712
transform 1 0 3164 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1712622712
transform 1 0 3060 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1712622712
transform 1 0 3052 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1712622712
transform 1 0 2908 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1712622712
transform 1 0 2620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1712622712
transform 1 0 1628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1712622712
transform 1 0 1468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1712622712
transform 1 0 1444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1712622712
transform 1 0 1404 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1712622712
transform 1 0 2964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1712622712
transform 1 0 2868 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1712622712
transform 1 0 2820 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1712622712
transform 1 0 2628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1712622712
transform 1 0 2556 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1712622712
transform 1 0 2420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1712622712
transform 1 0 2140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1712622712
transform 1 0 1588 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1712622712
transform 1 0 1540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1712622712
transform 1 0 1500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1712622712
transform 1 0 1452 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1712622712
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1712622712
transform 1 0 1316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1712622712
transform 1 0 1244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1712622712
transform 1 0 1060 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1712622712
transform 1 0 1044 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1712622712
transform 1 0 956 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1712622712
transform 1 0 956 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1712622712
transform 1 0 2652 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1712622712
transform 1 0 2572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1712622712
transform 1 0 2412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1712622712
transform 1 0 2364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1712622712
transform 1 0 2188 0 1 1295
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1712622712
transform 1 0 1836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1712622712
transform 1 0 1796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1712622712
transform 1 0 1756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1712622712
transform 1 0 1628 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1712622712
transform 1 0 1420 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1712622712
transform 1 0 1276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1712622712
transform 1 0 1148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1712622712
transform 1 0 1060 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1712622712
transform 1 0 988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1712622712
transform 1 0 892 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1712622712
transform 1 0 812 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1712622712
transform 1 0 812 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1712622712
transform 1 0 3116 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1712622712
transform 1 0 3084 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1712622712
transform 1 0 3084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1712622712
transform 1 0 3028 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1712622712
transform 1 0 2444 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1712622712
transform 1 0 2172 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1712622712
transform 1 0 2172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1712622712
transform 1 0 2156 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1712622712
transform 1 0 2124 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1712622712
transform 1 0 2012 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1712622712
transform 1 0 1980 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1712622712
transform 1 0 1940 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1712622712
transform 1 0 3052 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1712622712
transform 1 0 2988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1712622712
transform 1 0 2948 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1712622712
transform 1 0 2740 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1712622712
transform 1 0 2108 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1712622712
transform 1 0 1908 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1712622712
transform 1 0 1836 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1712622712
transform 1 0 1756 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1712622712
transform 1 0 1732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1712622712
transform 1 0 1716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1712622712
transform 1 0 2436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1712622712
transform 1 0 2396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1712622712
transform 1 0 2396 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1712622712
transform 1 0 2348 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1712622712
transform 1 0 2276 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1712622712
transform 1 0 2276 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1712622712
transform 1 0 2276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1712622712
transform 1 0 2252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1712622712
transform 1 0 2244 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1712622712
transform 1 0 2244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1712622712
transform 1 0 2156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1712622712
transform 1 0 2132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1712622712
transform 1 0 2188 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1712622712
transform 1 0 2180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1712622712
transform 1 0 2156 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1712622712
transform 1 0 2076 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1712622712
transform 1 0 1892 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1712622712
transform 1 0 1860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1712622712
transform 1 0 1812 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1712622712
transform 1 0 1780 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1712622712
transform 1 0 1612 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1712622712
transform 1 0 1604 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1712622712
transform 1 0 2388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1712622712
transform 1 0 2308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1712622712
transform 1 0 2284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1712622712
transform 1 0 1724 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1712622712
transform 1 0 1540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1712622712
transform 1 0 1388 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1712622712
transform 1 0 1340 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1712622712
transform 1 0 1020 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1712622712
transform 1 0 820 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1712622712
transform 1 0 732 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1712622712
transform 1 0 668 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1712622712
transform 1 0 1356 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1712622712
transform 1 0 1340 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1712622712
transform 1 0 1300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1712622712
transform 1 0 1300 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1712622712
transform 1 0 1284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1712622712
transform 1 0 1276 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1712622712
transform 1 0 1260 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1712622712
transform 1 0 1260 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1712622712
transform 1 0 1148 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1712622712
transform 1 0 980 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1712622712
transform 1 0 964 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1712622712
transform 1 0 956 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1712622712
transform 1 0 948 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1712622712
transform 1 0 940 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1712622712
transform 1 0 892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1712622712
transform 1 0 844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1712622712
transform 1 0 788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1712622712
transform 1 0 692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1712622712
transform 1 0 628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1712622712
transform 1 0 596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1712622712
transform 1 0 596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1712622712
transform 1 0 588 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1712622712
transform 1 0 556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1712622712
transform 1 0 340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1712622712
transform 1 0 228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1712622712
transform 1 0 156 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1712622712
transform 1 0 1660 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1712622712
transform 1 0 1628 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1712622712
transform 1 0 1412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1712622712
transform 1 0 1236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1712622712
transform 1 0 724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1712622712
transform 1 0 324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1712622712
transform 1 0 324 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1712622712
transform 1 0 316 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1712622712
transform 1 0 284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1712622712
transform 1 0 252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1712622712
transform 1 0 188 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1712622712
transform 1 0 908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1712622712
transform 1 0 828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1712622712
transform 1 0 788 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1712622712
transform 1 0 620 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1712622712
transform 1 0 500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1712622712
transform 1 0 444 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1712622712
transform 1 0 340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1712622712
transform 1 0 292 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1712622712
transform 1 0 292 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1712622712
transform 1 0 124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1712622712
transform 1 0 1228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1712622712
transform 1 0 1228 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1712622712
transform 1 0 700 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1712622712
transform 1 0 668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1712622712
transform 1 0 652 0 1 1755
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1712622712
transform 1 0 644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1712622712
transform 1 0 396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1712622712
transform 1 0 356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1712622712
transform 1 0 324 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1712622712
transform 1 0 308 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1712622712
transform 1 0 292 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1712622712
transform 1 0 276 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1712622712
transform 1 0 1324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1712622712
transform 1 0 1324 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1712622712
transform 1 0 1292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1712622712
transform 1 0 1292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1712622712
transform 1 0 1292 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1712622712
transform 1 0 1244 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1712622712
transform 1 0 1212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1712622712
transform 1 0 1148 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1712622712
transform 1 0 1148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1712622712
transform 1 0 1148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1712622712
transform 1 0 1044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1712622712
transform 1 0 1028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1712622712
transform 1 0 980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1712622712
transform 1 0 948 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1712622712
transform 1 0 892 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1712622712
transform 1 0 860 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1712622712
transform 1 0 820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1712622712
transform 1 0 764 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1712622712
transform 1 0 668 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1712622712
transform 1 0 628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1712622712
transform 1 0 3436 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1712622712
transform 1 0 3436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1712622712
transform 1 0 3420 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1712622712
transform 1 0 3380 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1712622712
transform 1 0 3372 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1712622712
transform 1 0 3276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1712622712
transform 1 0 3260 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1712622712
transform 1 0 3260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1712622712
transform 1 0 3236 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1712622712
transform 1 0 3172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1712622712
transform 1 0 3036 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1712622712
transform 1 0 3396 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1712622712
transform 1 0 3204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1712622712
transform 1 0 3148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1712622712
transform 1 0 3076 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1712622712
transform 1 0 3364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1712622712
transform 1 0 2916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1712622712
transform 1 0 2692 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1712622712
transform 1 0 1748 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1712622712
transform 1 0 3284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1712622712
transform 1 0 3132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1712622712
transform 1 0 2692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1712622712
transform 1 0 2676 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1712622712
transform 1 0 2676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1712622712
transform 1 0 2660 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1712622712
transform 1 0 2628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1712622712
transform 1 0 2628 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1712622712
transform 1 0 2620 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1712622712
transform 1 0 2620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1712622712
transform 1 0 1684 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1712622712
transform 1 0 1636 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1712622712
transform 1 0 1620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1712622712
transform 1 0 1564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1712622712
transform 1 0 1444 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1712622712
transform 1 0 1068 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1712622712
transform 1 0 1404 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1712622712
transform 1 0 1356 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1712622712
transform 1 0 1268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1712622712
transform 1 0 1260 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1712622712
transform 1 0 1188 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1712622712
transform 1 0 2996 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1712622712
transform 1 0 2980 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1712622712
transform 1 0 2916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1712622712
transform 1 0 2836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1712622712
transform 1 0 2716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1712622712
transform 1 0 2348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1712622712
transform 1 0 1604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1712622712
transform 1 0 1580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1712622712
transform 1 0 1460 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1712622712
transform 1 0 1332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1712622712
transform 1 0 3276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1712622712
transform 1 0 3212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1712622712
transform 1 0 3172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1712622712
transform 1 0 3052 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1712622712
transform 1 0 3004 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1712622712
transform 1 0 3244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1712622712
transform 1 0 2796 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1712622712
transform 1 0 1620 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1712622712
transform 1 0 3332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1712622712
transform 1 0 3228 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1712622712
transform 1 0 3228 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1712622712
transform 1 0 3180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1712622712
transform 1 0 3196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1712622712
transform 1 0 2364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1712622712
transform 1 0 2892 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1712622712
transform 1 0 2860 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1712622712
transform 1 0 3404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1712622712
transform 1 0 3396 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1712622712
transform 1 0 3396 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1712622712
transform 1 0 3324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1712622712
transform 1 0 1444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1712622712
transform 1 0 1316 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1712622712
transform 1 0 1276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1712622712
transform 1 0 1188 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1712622712
transform 1 0 1148 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1712622712
transform 1 0 1428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1712622712
transform 1 0 1308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1712622712
transform 1 0 836 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1712622712
transform 1 0 708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1712622712
transform 1 0 700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1712622712
transform 1 0 676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1712622712
transform 1 0 1388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1712622712
transform 1 0 1308 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1712622712
transform 1 0 1236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1712622712
transform 1 0 1068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1712622712
transform 1 0 964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1712622712
transform 1 0 836 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1712622712
transform 1 0 2300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1712622712
transform 1 0 2300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1712622712
transform 1 0 2284 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1712622712
transform 1 0 2268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1712622712
transform 1 0 2260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1712622712
transform 1 0 2044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1712622712
transform 1 0 1964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1712622712
transform 1 0 1948 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1712622712
transform 1 0 1580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1712622712
transform 1 0 1564 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1712622712
transform 1 0 1564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1712622712
transform 1 0 1444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1712622712
transform 1 0 1372 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1712622712
transform 1 0 908 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1712622712
transform 1 0 740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1712622712
transform 1 0 1084 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1712622712
transform 1 0 700 0 1 1685
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1712622712
transform 1 0 540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1712622712
transform 1 0 524 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1712622712
transform 1 0 476 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1712622712
transform 1 0 476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1712622712
transform 1 0 244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1712622712
transform 1 0 212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1712622712
transform 1 0 3084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1712622712
transform 1 0 3044 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1712622712
transform 1 0 3028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1712622712
transform 1 0 2740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1712622712
transform 1 0 2684 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1712622712
transform 1 0 2164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1712622712
transform 1 0 2084 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1712622712
transform 1 0 1108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1712622712
transform 1 0 900 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1712622712
transform 1 0 596 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1712622712
transform 1 0 540 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1712622712
transform 1 0 316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1712622712
transform 1 0 220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1712622712
transform 1 0 212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1712622712
transform 1 0 2652 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1712622712
transform 1 0 2564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1712622712
transform 1 0 2540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1712622712
transform 1 0 2500 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1712622712
transform 1 0 2348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1712622712
transform 1 0 2340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1712622712
transform 1 0 2316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1712622712
transform 1 0 2148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1712622712
transform 1 0 2060 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1712622712
transform 1 0 2052 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1712622712
transform 1 0 1868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1712622712
transform 1 0 1852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1712622712
transform 1 0 1748 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1712622712
transform 1 0 1636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1712622712
transform 1 0 1340 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1712622712
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1712622712
transform 1 0 1164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1712622712
transform 1 0 892 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1712622712
transform 1 0 724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1712622712
transform 1 0 684 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1712622712
transform 1 0 516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1712622712
transform 1 0 484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1712622712
transform 1 0 436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1712622712
transform 1 0 436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1712622712
transform 1 0 420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1712622712
transform 1 0 420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1712622712
transform 1 0 420 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1712622712
transform 1 0 412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1712622712
transform 1 0 412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1712622712
transform 1 0 380 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1712622712
transform 1 0 372 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1712622712
transform 1 0 2724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1712622712
transform 1 0 2716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1712622712
transform 1 0 2692 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1712622712
transform 1 0 2580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1712622712
transform 1 0 2204 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1712622712
transform 1 0 2188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1712622712
transform 1 0 2180 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1712622712
transform 1 0 3420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1712622712
transform 1 0 3364 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1712622712
transform 1 0 3260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1712622712
transform 1 0 3260 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1712622712
transform 1 0 3188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1712622712
transform 1 0 3076 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1712622712
transform 1 0 3068 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1712622712
transform 1 0 2972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1712622712
transform 1 0 3340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1712622712
transform 1 0 3284 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1712622712
transform 1 0 3148 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1712622712
transform 1 0 3148 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1712622712
transform 1 0 3004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1712622712
transform 1 0 2964 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1712622712
transform 1 0 2948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1712622712
transform 1 0 2940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1712622712
transform 1 0 3436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1712622712
transform 1 0 3388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1712622712
transform 1 0 3300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1712622712
transform 1 0 3244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1712622712
transform 1 0 3092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1712622712
transform 1 0 3084 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1712622712
transform 1 0 2980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1712622712
transform 1 0 2980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1712622712
transform 1 0 2892 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1712622712
transform 1 0 2860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1712622712
transform 1 0 3388 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1712622712
transform 1 0 3356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1712622712
transform 1 0 3364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1712622712
transform 1 0 3348 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1712622712
transform 1 0 3420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1712622712
transform 1 0 3372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1712622712
transform 1 0 3356 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1712622712
transform 1 0 2980 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1712622712
transform 1 0 2908 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1712622712
transform 1 0 2812 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1712622712
transform 1 0 2748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1712622712
transform 1 0 3348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1712622712
transform 1 0 3300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1712622712
transform 1 0 2732 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1712622712
transform 1 0 2652 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1712622712
transform 1 0 2652 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1712622712
transform 1 0 2620 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1712622712
transform 1 0 2548 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1712622712
transform 1 0 3220 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1712622712
transform 1 0 2748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1712622712
transform 1 0 2628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1712622712
transform 1 0 2628 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1712622712
transform 1 0 2580 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1712622712
transform 1 0 2572 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1712622712
transform 1 0 2532 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1712622712
transform 1 0 2532 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1712622712
transform 1 0 3220 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1712622712
transform 1 0 3124 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1712622712
transform 1 0 2700 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1712622712
transform 1 0 2660 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1712622712
transform 1 0 2636 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1712622712
transform 1 0 2628 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1712622712
transform 1 0 2612 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1712622712
transform 1 0 2612 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1712622712
transform 1 0 2612 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1712622712
transform 1 0 2924 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1712622712
transform 1 0 2724 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1712622712
transform 1 0 2668 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1712622712
transform 1 0 2660 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1712622712
transform 1 0 2780 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1712622712
transform 1 0 2772 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1712622712
transform 1 0 2716 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1712622712
transform 1 0 2692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1712622712
transform 1 0 2668 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1712622712
transform 1 0 3388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1712622712
transform 1 0 3388 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1712622712
transform 1 0 3260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1712622712
transform 1 0 3132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1712622712
transform 1 0 3220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1712622712
transform 1 0 3164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1712622712
transform 1 0 3012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1712622712
transform 1 0 3004 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1712622712
transform 1 0 2796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1712622712
transform 1 0 2772 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1712622712
transform 1 0 3396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1712622712
transform 1 0 3300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1712622712
transform 1 0 3260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1712622712
transform 1 0 3172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1712622712
transform 1 0 2724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1712622712
transform 1 0 2724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1712622712
transform 1 0 2924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1712622712
transform 1 0 2916 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1712622712
transform 1 0 3012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1712622712
transform 1 0 3012 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1712622712
transform 1 0 2860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1712622712
transform 1 0 2820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1712622712
transform 1 0 2628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1712622712
transform 1 0 2620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1712622712
transform 1 0 2508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1712622712
transform 1 0 2508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1712622712
transform 1 0 2404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1712622712
transform 1 0 2396 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1712622712
transform 1 0 2132 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1712622712
transform 1 0 2132 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1712622712
transform 1 0 1940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1712622712
transform 1 0 1932 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1712622712
transform 1 0 2260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1712622712
transform 1 0 2228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1712622712
transform 1 0 2324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1712622712
transform 1 0 2324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1712622712
transform 1 0 2068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1712622712
transform 1 0 2028 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1712622712
transform 1 0 1876 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1712622712
transform 1 0 1828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1712622712
transform 1 0 1812 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1712622712
transform 1 0 1692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1712622712
transform 1 0 1684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1712622712
transform 1 0 1580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1712622712
transform 1 0 1500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1712622712
transform 1 0 1500 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1712622712
transform 1 0 1436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1712622712
transform 1 0 1420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1712622712
transform 1 0 1316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1712622712
transform 1 0 1308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1712622712
transform 1 0 1124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1712622712
transform 1 0 1084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1712622712
transform 1 0 1004 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1712622712
transform 1 0 988 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1712622712
transform 1 0 572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1712622712
transform 1 0 572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1712622712
transform 1 0 172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1712622712
transform 1 0 148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1712622712
transform 1 0 116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1712622712
transform 1 0 116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1712622712
transform 1 0 244 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1712622712
transform 1 0 188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1712622712
transform 1 0 292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1712622712
transform 1 0 244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1712622712
transform 1 0 340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1712622712
transform 1 0 244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1712622712
transform 1 0 420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1712622712
transform 1 0 364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1712622712
transform 1 0 484 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1712622712
transform 1 0 476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1712622712
transform 1 0 684 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1712622712
transform 1 0 684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1712622712
transform 1 0 780 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1712622712
transform 1 0 780 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1712622712
transform 1 0 924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1712622712
transform 1 0 916 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1712622712
transform 1 0 1364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1712622712
transform 1 0 1212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1712622712
transform 1 0 2932 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1712622712
transform 1 0 2932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1712622712
transform 1 0 2092 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1712622712
transform 1 0 1732 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1712622712
transform 1 0 2564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1712622712
transform 1 0 2548 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1712622712
transform 1 0 3420 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1712622712
transform 1 0 3380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1712622712
transform 1 0 3228 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1712622712
transform 1 0 3044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1712622712
transform 1 0 2924 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1712622712
transform 1 0 2868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1712622712
transform 1 0 3252 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1712622712
transform 1 0 3244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1712622712
transform 1 0 3212 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1712622712
transform 1 0 2772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1712622712
transform 1 0 2724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1712622712
transform 1 0 2612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1712622712
transform 1 0 3372 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1712622712
transform 1 0 3340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1712622712
transform 1 0 3308 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1712622712
transform 1 0 3404 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1712622712
transform 1 0 3308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1712622712
transform 1 0 3284 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1712622712
transform 1 0 2940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1712622712
transform 1 0 1756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1712622712
transform 1 0 1724 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1712622712
transform 1 0 1668 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1712622712
transform 1 0 1740 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1712622712
transform 1 0 1580 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1712622712
transform 1 0 1556 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1712622712
transform 1 0 1532 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1712622712
transform 1 0 1532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1712622712
transform 1 0 1468 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1712622712
transform 1 0 1508 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1712622712
transform 1 0 1484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1712622712
transform 1 0 1540 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1712622712
transform 1 0 1476 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1712622712
transform 1 0 1492 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1712622712
transform 1 0 1492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1712622712
transform 1 0 1460 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1712622712
transform 1 0 1452 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1712622712
transform 1 0 2068 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1712622712
transform 1 0 1452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1712622712
transform 1 0 1460 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1712622712
transform 1 0 980 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1712622712
transform 1 0 924 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1712622712
transform 1 0 276 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1712622712
transform 1 0 988 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1712622712
transform 1 0 988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1712622712
transform 1 0 1100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1712622712
transform 1 0 956 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1712622712
transform 1 0 972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1712622712
transform 1 0 684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1712622712
transform 1 0 1004 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1712622712
transform 1 0 964 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1712622712
transform 1 0 1684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1712622712
transform 1 0 996 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1712622712
transform 1 0 780 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1712622712
transform 1 0 1068 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1712622712
transform 1 0 1020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1712622712
transform 1 0 1540 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1712622712
transform 1 0 1436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1712622712
transform 1 0 1372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1712622712
transform 1 0 1052 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1712622712
transform 1 0 1244 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1712622712
transform 1 0 1172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1712622712
transform 1 0 1084 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1712622712
transform 1 0 1084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1712622712
transform 1 0 652 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1712622712
transform 1 0 548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1712622712
transform 1 0 388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1712622712
transform 1 0 692 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1712622712
transform 1 0 644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1712622712
transform 1 0 1148 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1712622712
transform 1 0 1084 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1712622712
transform 1 0 1044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1712622712
transform 1 0 900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1712622712
transform 1 0 836 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1712622712
transform 1 0 1372 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1712622712
transform 1 0 1164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1712622712
transform 1 0 1116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1712622712
transform 1 0 1116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1712622712
transform 1 0 204 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1712622712
transform 1 0 204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1712622712
transform 1 0 244 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1712622712
transform 1 0 236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1712622712
transform 1 0 236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1712622712
transform 1 0 220 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1712622712
transform 1 0 268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1712622712
transform 1 0 204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1712622712
transform 1 0 196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1712622712
transform 1 0 220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1712622712
transform 1 0 172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1712622712
transform 1 0 308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1712622712
transform 1 0 252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1712622712
transform 1 0 204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1712622712
transform 1 0 532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1712622712
transform 1 0 260 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1712622712
transform 1 0 252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1712622712
transform 1 0 268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1712622712
transform 1 0 236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1712622712
transform 1 0 228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1712622712
transform 1 0 316 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1712622712
transform 1 0 276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1712622712
transform 1 0 212 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1712622712
transform 1 0 516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1712622712
transform 1 0 172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1712622712
transform 1 0 172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1712622712
transform 1 0 212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1712622712
transform 1 0 212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1712622712
transform 1 0 2108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1712622712
transform 1 0 2108 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1712622712
transform 1 0 2212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1712622712
transform 1 0 2132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1712622712
transform 1 0 2252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1712622712
transform 1 0 2212 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1712622712
transform 1 0 2212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1712622712
transform 1 0 1788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1712622712
transform 1 0 1764 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1712622712
transform 1 0 1764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1712622712
transform 1 0 2300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1712622712
transform 1 0 2292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1712622712
transform 1 0 2236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1712622712
transform 1 0 2236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1712622712
transform 1 0 2324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1712622712
transform 1 0 2204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1712622712
transform 1 0 2196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1712622712
transform 1 0 2092 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1712622712
transform 1 0 2092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1712622712
transform 1 0 2364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1712622712
transform 1 0 2132 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1712622712
transform 1 0 2364 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1712622712
transform 1 0 2356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1712622712
transform 1 0 2340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1712622712
transform 1 0 2332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1712622712
transform 1 0 2324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1712622712
transform 1 0 2388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1712622712
transform 1 0 2388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1712622712
transform 1 0 2340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1712622712
transform 1 0 2340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1712622712
transform 1 0 2100 0 1 1885
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1712622712
transform 1 0 2084 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1712622712
transform 1 0 2100 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1712622712
transform 1 0 1956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1712622712
transform 1 0 1924 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1712622712
transform 1 0 1452 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1712622712
transform 1 0 1428 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1712622712
transform 1 0 1444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1712622712
transform 1 0 1076 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1712622712
transform 1 0 1044 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1712622712
transform 1 0 964 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1712622712
transform 1 0 1068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1712622712
transform 1 0 1052 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1712622712
transform 1 0 956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1712622712
transform 1 0 972 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1712622712
transform 1 0 876 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1712622712
transform 1 0 876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1712622712
transform 1 0 428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1712622712
transform 1 0 428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1712622712
transform 1 0 332 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1712622712
transform 1 0 1572 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1712622712
transform 1 0 1492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1712622712
transform 1 0 2244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1712622712
transform 1 0 1516 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1712622712
transform 1 0 2428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1712622712
transform 1 0 2308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1712622712
transform 1 0 2204 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1712622712
transform 1 0 2260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1712622712
transform 1 0 2252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1712622712
transform 1 0 2148 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1712622712
transform 1 0 1700 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1712622712
transform 1 0 1596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1712622712
transform 1 0 1564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1712622712
transform 1 0 1580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1712622712
transform 1 0 1444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1712622712
transform 1 0 1284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1712622712
transform 1 0 1908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1712622712
transform 1 0 1508 0 1 1695
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1712622712
transform 1 0 1708 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1712622712
transform 1 0 1524 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1712622712
transform 1 0 1524 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1712622712
transform 1 0 396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1712622712
transform 1 0 460 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1712622712
transform 1 0 396 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1712622712
transform 1 0 380 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1712622712
transform 1 0 380 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1712622712
transform 1 0 436 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1712622712
transform 1 0 404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1712622712
transform 1 0 428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1712622712
transform 1 0 420 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1712622712
transform 1 0 428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1712622712
transform 1 0 420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1712622712
transform 1 0 772 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1712622712
transform 1 0 412 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1712622712
transform 1 0 875 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1712622712
transform 1 0 804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1712622712
transform 1 0 924 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1712622712
transform 1 0 820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1712622712
transform 1 0 820 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1712622712
transform 1 0 892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1712622712
transform 1 0 748 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1712622712
transform 1 0 748 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1712622712
transform 1 0 2980 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1712622712
transform 1 0 2868 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1712622712
transform 1 0 2588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1712622712
transform 1 0 2588 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1712622712
transform 1 0 2508 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1712622712
transform 1 0 1668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1712622712
transform 1 0 1652 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1712622712
transform 1 0 1644 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1712622712
transform 1 0 1620 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1712622712
transform 1 0 2652 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1712622712
transform 1 0 2604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1712622712
transform 1 0 1652 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1712622712
transform 1 0 492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1712622712
transform 1 0 444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1712622712
transform 1 0 420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1712622712
transform 1 0 444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1712622712
transform 1 0 436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1712622712
transform 1 0 380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1712622712
transform 1 0 396 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1712622712
transform 1 0 396 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1712622712
transform 1 0 476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1712622712
transform 1 0 476 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1712622712
transform 1 0 452 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1712622712
transform 1 0 444 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1712622712
transform 1 0 484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1712622712
transform 1 0 412 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1712622712
transform 1 0 980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1712622712
transform 1 0 412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1712622712
transform 1 0 444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1712622712
transform 1 0 420 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1712622712
transform 1 0 500 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1712622712
transform 1 0 420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1712622712
transform 1 0 420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1712622712
transform 1 0 460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1712622712
transform 1 0 444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1712622712
transform 1 0 460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1712622712
transform 1 0 444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1712622712
transform 1 0 436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1712622712
transform 1 0 436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1712622712
transform 1 0 508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1712622712
transform 1 0 476 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1712622712
transform 1 0 476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1712622712
transform 1 0 1188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1712622712
transform 1 0 1004 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1712622712
transform 1 0 956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1712622712
transform 1 0 988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1712622712
transform 1 0 948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1712622712
transform 1 0 884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1712622712
transform 1 0 540 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1712622712
transform 1 0 476 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1712622712
transform 1 0 492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1712622712
transform 1 0 460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1712622712
transform 1 0 388 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1712622712
transform 1 0 1772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1712622712
transform 1 0 1684 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1712622712
transform 1 0 1772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1712622712
transform 1 0 1740 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1712622712
transform 1 0 1628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1712622712
transform 1 0 1652 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1712622712
transform 1 0 1572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1712622712
transform 1 0 1524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1712622712
transform 1 0 956 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1712622712
transform 1 0 812 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1712622712
transform 1 0 644 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1712622712
transform 1 0 1532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1712622712
transform 1 0 1308 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1712622712
transform 1 0 1308 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1712622712
transform 1 0 1588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1712622712
transform 1 0 1492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1712622712
transform 1 0 1492 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1712622712
transform 1 0 932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1712622712
transform 1 0 628 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1712622712
transform 1 0 148 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1712622712
transform 1 0 92 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1712622712
transform 1 0 1580 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1712622712
transform 1 0 1580 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1712622712
transform 1 0 1572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1712622712
transform 1 0 1764 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1712622712
transform 1 0 1740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1712622712
transform 1 0 2244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1712622712
transform 1 0 1836 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1712622712
transform 1 0 2492 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1712622712
transform 1 0 2372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1712622712
transform 1 0 2268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1712622712
transform 1 0 2196 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1712622712
transform 1 0 2188 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1712622712
transform 1 0 2364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1712622712
transform 1 0 2236 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1712622712
transform 1 0 2500 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1712622712
transform 1 0 2276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1712622712
transform 1 0 2276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1712622712
transform 1 0 2236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1712622712
transform 1 0 2236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1712622712
transform 1 0 2260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1712622712
transform 1 0 2172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1712622712
transform 1 0 2164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1712622712
transform 1 0 2444 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1712622712
transform 1 0 2228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1712622712
transform 1 0 1868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1712622712
transform 1 0 1868 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1712622712
transform 1 0 1804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1712622712
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1712622712
transform 1 0 1940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1712622712
transform 1 0 1940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1712622712
transform 1 0 1732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1712622712
transform 1 0 1652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1712622712
transform 1 0 1388 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1712622712
transform 1 0 1388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1712622712
transform 1 0 2588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1712622712
transform 1 0 1900 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1712622712
transform 1 0 1916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1712622712
transform 1 0 1908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1712622712
transform 1 0 1844 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1712622712
transform 1 0 1292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1712622712
transform 1 0 1268 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1712622712
transform 1 0 2204 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1712622712
transform 1 0 2156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1712622712
transform 1 0 1844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1712622712
transform 1 0 1828 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1712622712
transform 1 0 1796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1712622712
transform 1 0 1748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1712622712
transform 1 0 1540 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1712622712
transform 1 0 1940 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1712622712
transform 1 0 1940 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1712622712
transform 1 0 2116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1712622712
transform 1 0 2116 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1712622712
transform 1 0 1932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1712622712
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1712622712
transform 1 0 1876 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1712622712
transform 1 0 1764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1712622712
transform 1 0 2636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1712622712
transform 1 0 2596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1712622712
transform 1 0 2660 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1712622712
transform 1 0 2580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1712622712
transform 1 0 2588 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1712622712
transform 1 0 2572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1712622712
transform 1 0 2572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1712622712
transform 1 0 2588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1712622712
transform 1 0 2524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1712622712
transform 1 0 2492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1712622712
transform 1 0 2564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1712622712
transform 1 0 2556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1712622712
transform 1 0 2652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1712622712
transform 1 0 2452 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1712622712
transform 1 0 2452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1712622712
transform 1 0 1652 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1712622712
transform 1 0 1404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1712622712
transform 1 0 1412 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1712622712
transform 1 0 884 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1712622712
transform 1 0 836 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1712622712
transform 1 0 580 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1712622712
transform 1 0 876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1712622712
transform 1 0 868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1712622712
transform 1 0 860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1712622712
transform 1 0 860 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1712622712
transform 1 0 852 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1712622712
transform 1 0 652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1712622712
transform 1 0 1668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1712622712
transform 1 0 892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1712622712
transform 1 0 1668 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1712622712
transform 1 0 1068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1712622712
transform 1 0 1140 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1712622712
transform 1 0 1044 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1712622712
transform 1 0 924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1712622712
transform 1 0 1204 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1712622712
transform 1 0 1084 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1712622712
transform 1 0 988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1712622712
transform 1 0 2596 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1712622712
transform 1 0 2572 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1712622712
transform 1 0 1684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1712622712
transform 1 0 596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1712622712
transform 1 0 508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1712622712
transform 1 0 652 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1712622712
transform 1 0 540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1712622712
transform 1 0 644 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1712622712
transform 1 0 516 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1712622712
transform 1 0 508 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1712622712
transform 1 0 620 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1712622712
transform 1 0 556 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1712622712
transform 1 0 556 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1712622712
transform 1 0 668 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1712622712
transform 1 0 572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1712622712
transform 1 0 524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1712622712
transform 1 0 492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1712622712
transform 1 0 724 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1712622712
transform 1 0 652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1712622712
transform 1 0 556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1712622712
transform 1 0 1044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1712622712
transform 1 0 852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1712622712
transform 1 0 860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1712622712
transform 1 0 756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1712622712
transform 1 0 772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1712622712
transform 1 0 756 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1712622712
transform 1 0 748 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1712622712
transform 1 0 772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1712622712
transform 1 0 756 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1712622712
transform 1 0 676 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1712622712
transform 1 0 1004 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1712622712
transform 1 0 996 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1712622712
transform 1 0 964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1712622712
transform 1 0 1108 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1712622712
transform 1 0 1060 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1712622712
transform 1 0 1060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1712622712
transform 1 0 2100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1712622712
transform 1 0 2084 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1712622712
transform 1 0 2084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1712622712
transform 1 0 2044 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1712622712
transform 1 0 1820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1712622712
transform 1 0 1316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1712622712
transform 1 0 1292 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1712622712
transform 1 0 1228 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1712622712
transform 1 0 1196 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1712622712
transform 1 0 652 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1712622712
transform 1 0 516 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1712622712
transform 1 0 516 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1712622712
transform 1 0 524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1712622712
transform 1 0 508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1712622712
transform 1 0 500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1712622712
transform 1 0 500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1712622712
transform 1 0 668 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1712622712
transform 1 0 564 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1712622712
transform 1 0 2308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1712622712
transform 1 0 1636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1712622712
transform 1 0 1756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1712622712
transform 1 0 1644 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1712622712
transform 1 0 2308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1712622712
transform 1 0 1780 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1712622712
transform 1 0 1836 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1712622712
transform 1 0 1804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1712622712
transform 1 0 1876 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1712622712
transform 1 0 1852 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1712622712
transform 1 0 1884 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1712622712
transform 1 0 1860 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1712622712
transform 1 0 1892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1712622712
transform 1 0 1788 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1712622712
transform 1 0 1788 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1712622712
transform 1 0 2292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1712622712
transform 1 0 2292 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1712622712
transform 1 0 2132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1712622712
transform 1 0 2076 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1712622712
transform 1 0 2028 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1712622712
transform 1 0 2004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1712622712
transform 1 0 1956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1712622712
transform 1 0 1956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1712622712
transform 1 0 1916 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1712622712
transform 1 0 1580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1712622712
transform 1 0 1556 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1712622712
transform 1 0 1460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1712622712
transform 1 0 2404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1712622712
transform 1 0 2332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1712622712
transform 1 0 2388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1712622712
transform 1 0 2348 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1712622712
transform 1 0 2436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1712622712
transform 1 0 2372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1712622712
transform 1 0 2100 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1712622712
transform 1 0 2404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1712622712
transform 1 0 2180 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1712622712
transform 1 0 2420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1712622712
transform 1 0 2348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1712622712
transform 1 0 2220 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1712622712
transform 1 0 2420 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1712622712
transform 1 0 2316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1712622712
transform 1 0 2156 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1712622712
transform 1 0 2396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1712622712
transform 1 0 2276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1712622712
transform 1 0 2284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1712622712
transform 1 0 2260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1712622712
transform 1 0 2244 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1712622712
transform 1 0 2212 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1712622712
transform 1 0 2020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1712622712
transform 1 0 2308 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1712622712
transform 1 0 2292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1712622712
transform 1 0 2500 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1712622712
transform 1 0 2436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1712622712
transform 1 0 2380 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1712622712
transform 1 0 1556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1712622712
transform 1 0 1244 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1712622712
transform 1 0 1596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1712622712
transform 1 0 1580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1712622712
transform 1 0 1748 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1712622712
transform 1 0 1708 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1712622712
transform 1 0 1572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1712622712
transform 1 0 1612 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1712622712
transform 1 0 1476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1712622712
transform 1 0 1340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1712622712
transform 1 0 1228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1712622712
transform 1 0 1212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1712622712
transform 1 0 1140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1712622712
transform 1 0 1260 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1712622712
transform 1 0 1228 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1712622712
transform 1 0 1188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1712622712
transform 1 0 1428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1712622712
transform 1 0 1380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1712622712
transform 1 0 1300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1712622712
transform 1 0 468 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1712622712
transform 1 0 444 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1712622712
transform 1 0 196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1712622712
transform 1 0 100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1712622712
transform 1 0 2052 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1712622712
transform 1 0 1532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1712622712
transform 1 0 1540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1712622712
transform 1 0 820 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1712622712
transform 1 0 740 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1712622712
transform 1 0 532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1712622712
transform 1 0 772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1712622712
transform 1 0 764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1712622712
transform 1 0 796 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1712622712
transform 1 0 780 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1712622712
transform 1 0 772 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1712622712
transform 1 0 772 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1712622712
transform 1 0 932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1712622712
transform 1 0 820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1712622712
transform 1 0 1348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1712622712
transform 1 0 1292 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1712622712
transform 1 0 996 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1712622712
transform 1 0 908 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1712622712
transform 1 0 908 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1712622712
transform 1 0 884 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1712622712
transform 1 0 332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1712622712
transform 1 0 308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1712622712
transform 1 0 948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1712622712
transform 1 0 924 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1712622712
transform 1 0 1036 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1712622712
transform 1 0 1036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1712622712
transform 1 0 940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1712622712
transform 1 0 836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1712622712
transform 1 0 996 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1712622712
transform 1 0 956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1712622712
transform 1 0 924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1712622712
transform 1 0 948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1712622712
transform 1 0 788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1712622712
transform 1 0 804 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1712622712
transform 1 0 732 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1712622712
transform 1 0 1052 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1712622712
transform 1 0 980 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1712622712
transform 1 0 916 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1712622712
transform 1 0 684 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1712622712
transform 1 0 588 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1712622712
transform 1 0 588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1712622712
transform 1 0 756 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1712622712
transform 1 0 740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1712622712
transform 1 0 692 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1712622712
transform 1 0 684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1712622712
transform 1 0 668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1712622712
transform 1 0 1076 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1712622712
transform 1 0 1076 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1712622712
transform 1 0 956 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1712622712
transform 1 0 940 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1712622712
transform 1 0 900 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1712622712
transform 1 0 900 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1712622712
transform 1 0 892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1712622712
transform 1 0 1388 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1712622712
transform 1 0 1212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1712622712
transform 1 0 1020 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1712622712
transform 1 0 1020 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1712622712
transform 1 0 956 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1712622712
transform 1 0 812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1712622712
transform 1 0 732 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1712622712
transform 1 0 684 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1712622712
transform 1 0 620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1712622712
transform 1 0 860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1712622712
transform 1 0 804 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1712622712
transform 1 0 636 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1712622712
transform 1 0 588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1712622712
transform 1 0 580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1712622712
transform 1 0 580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1712622712
transform 1 0 988 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1712622712
transform 1 0 900 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1712622712
transform 1 0 788 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1712622712
transform 1 0 684 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1712622712
transform 1 0 636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1712622712
transform 1 0 636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1712622712
transform 1 0 2484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1712622712
transform 1 0 2460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1712622712
transform 1 0 2460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1712622712
transform 1 0 2444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1712622712
transform 1 0 2444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1712622712
transform 1 0 1484 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1712622712
transform 1 0 1140 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1712622712
transform 1 0 1092 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1712622712
transform 1 0 1044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1712622712
transform 1 0 1036 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1712622712
transform 1 0 996 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1712622712
transform 1 0 796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1712622712
transform 1 0 612 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1712622712
transform 1 0 612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1712622712
transform 1 0 1004 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1712622712
transform 1 0 852 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1712622712
transform 1 0 668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1712622712
transform 1 0 588 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1712622712
transform 1 0 500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1712622712
transform 1 0 572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1712622712
transform 1 0 500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1712622712
transform 1 0 828 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1712622712
transform 1 0 812 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1712622712
transform 1 0 748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1712622712
transform 1 0 724 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1712622712
transform 1 0 580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1712622712
transform 1 0 548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1712622712
transform 1 0 796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1712622712
transform 1 0 708 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1712622712
transform 1 0 692 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1712622712
transform 1 0 668 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1712622712
transform 1 0 652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1712622712
transform 1 0 588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1712622712
transform 1 0 588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1712622712
transform 1 0 2060 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1712622712
transform 1 0 2028 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1712622712
transform 1 0 2532 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1712622712
transform 1 0 2028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1712622712
transform 1 0 2028 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1712622712
transform 1 0 2020 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1712622712
transform 1 0 2044 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1712622712
transform 1 0 2020 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1712622712
transform 1 0 2036 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1712622712
transform 1 0 1452 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1712622712
transform 1 0 2316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1712622712
transform 1 0 2284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1712622712
transform 1 0 2260 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1712622712
transform 1 0 2196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1712622712
transform 1 0 1820 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1712622712
transform 1 0 1748 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1712622712
transform 1 0 1732 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1712622712
transform 1 0 1668 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1712622712
transform 1 0 1588 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1712622712
transform 1 0 1436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1712622712
transform 1 0 1412 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1712622712
transform 1 0 1460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1712622712
transform 1 0 1412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1712622712
transform 1 0 1492 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1712622712
transform 1 0 1484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1712622712
transform 1 0 1404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1712622712
transform 1 0 1364 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1712622712
transform 1 0 1364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1712622712
transform 1 0 1236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1712622712
transform 1 0 1476 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1712622712
transform 1 0 1420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1712622712
transform 1 0 1180 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1712622712
transform 1 0 1172 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1712622712
transform 1 0 1172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1712622712
transform 1 0 1156 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1712622712
transform 1 0 2044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1712622712
transform 1 0 1996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1712622712
transform 1 0 2252 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1712622712
transform 1 0 2092 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1712622712
transform 1 0 2524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1712622712
transform 1 0 2516 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1712622712
transform 1 0 2196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1712622712
transform 1 0 2012 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1712622712
transform 1 0 1612 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1712622712
transform 1 0 1596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1712622712
transform 1 0 2332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1712622712
transform 1 0 2308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1712622712
transform 1 0 2260 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1712622712
transform 1 0 2252 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1712622712
transform 1 0 1900 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1712622712
transform 1 0 1892 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1712622712
transform 1 0 1820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1712622712
transform 1 0 1940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1712622712
transform 1 0 1924 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1712622712
transform 1 0 1916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1712622712
transform 1 0 1876 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1712622712
transform 1 0 1852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1712622712
transform 1 0 2004 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1712622712
transform 1 0 1820 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1712622712
transform 1 0 1724 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1712622712
transform 1 0 1724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1712622712
transform 1 0 1628 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1712622712
transform 1 0 1604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1712622712
transform 1 0 2612 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1712622712
transform 1 0 2508 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1712622712
transform 1 0 2460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1712622712
transform 1 0 2436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1712622712
transform 1 0 2428 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1712622712
transform 1 0 2428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1712622712
transform 1 0 2412 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1712622712
transform 1 0 2388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1712622712
transform 1 0 2388 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1712622712
transform 1 0 2348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1712622712
transform 1 0 2340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1712622712
transform 1 0 2652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1712622712
transform 1 0 2548 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1712622712
transform 1 0 2548 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1712622712
transform 1 0 2524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1712622712
transform 1 0 2516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1712622712
transform 1 0 2476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1712622712
transform 1 0 2132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1712622712
transform 1 0 2100 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1712622712
transform 1 0 3108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1712622712
transform 1 0 3028 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1712622712
transform 1 0 2972 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1712622712
transform 1 0 2908 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1712622712
transform 1 0 2548 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1712622712
transform 1 0 2500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1712622712
transform 1 0 2276 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1712622712
transform 1 0 2260 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1712622712
transform 1 0 2244 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1712622712
transform 1 0 2148 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1712622712
transform 1 0 2148 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1712622712
transform 1 0 2140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1712622712
transform 1 0 2052 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1712622712
transform 1 0 2028 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1712622712
transform 1 0 2060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1712622712
transform 1 0 2004 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1712622712
transform 1 0 1916 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1712622712
transform 1 0 1868 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1712622712
transform 1 0 1788 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1712622712
transform 1 0 1732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1712622712
transform 1 0 2260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1712622712
transform 1 0 2132 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1712622712
transform 1 0 2116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1712622712
transform 1 0 2076 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1712622712
transform 1 0 2052 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1712622712
transform 1 0 1980 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1712622712
transform 1 0 1668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1712622712
transform 1 0 1628 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1712622712
transform 1 0 1652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1712622712
transform 1 0 1652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1712622712
transform 1 0 1628 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1712622712
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1712622712
transform 1 0 3308 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1712622712
transform 1 0 1932 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1712622712
transform 1 0 1636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1712622712
transform 1 0 1588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1712622712
transform 1 0 1564 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1712622712
transform 1 0 1348 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1712622712
transform 1 0 1620 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1712622712
transform 1 0 1620 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1712622712
transform 1 0 1564 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1712622712
transform 1 0 1548 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1712622712
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1712622712
transform 1 0 1604 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1712622712
transform 1 0 1612 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1712622712
transform 1 0 1524 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1712622712
transform 1 0 1508 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1712622712
transform 1 0 372 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1712622712
transform 1 0 1572 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1712622712
transform 1 0 1524 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1712622712
transform 1 0 1540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1712622712
transform 1 0 1524 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1712622712
transform 1 0 1532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1712622712
transform 1 0 1508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1712622712
transform 1 0 1468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1712622712
transform 1 0 1452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1712622712
transform 1 0 1540 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1712622712
transform 1 0 804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1712622712
transform 1 0 764 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1712622712
transform 1 0 724 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1712622712
transform 1 0 724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1712622712
transform 1 0 572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1712622712
transform 1 0 516 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1712622712
transform 1 0 524 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1712622712
transform 1 0 476 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1712622712
transform 1 0 460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1712622712
transform 1 0 524 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1712622712
transform 1 0 380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1712622712
transform 1 0 1524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1712622712
transform 1 0 1340 0 1 1934
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1712622712
transform 1 0 1300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1712622712
transform 1 0 2068 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1712622712
transform 1 0 2044 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1712622712
transform 1 0 1900 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1712622712
transform 1 0 1884 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1712622712
transform 1 0 1580 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1712622712
transform 1 0 356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1712622712
transform 1 0 340 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1712622712
transform 1 0 380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1712622712
transform 1 0 356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1712622712
transform 1 0 428 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1712622712
transform 1 0 356 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1712622712
transform 1 0 404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1712622712
transform 1 0 404 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1712622712
transform 1 0 388 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1712622712
transform 1 0 388 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1712622712
transform 1 0 388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1712622712
transform 1 0 372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1712622712
transform 1 0 428 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1712622712
transform 1 0 364 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1712622712
transform 1 0 364 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1712622712
transform 1 0 340 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1712622712
transform 1 0 340 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1712622712
transform 1 0 452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1712622712
transform 1 0 444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1712622712
transform 1 0 412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1712622712
transform 1 0 332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1712622712
transform 1 0 476 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1712622712
transform 1 0 412 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1712622712
transform 1 0 364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1712622712
transform 1 0 396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1712622712
transform 1 0 356 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1712622712
transform 1 0 452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1712622712
transform 1 0 420 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1712622712
transform 1 0 340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1712622712
transform 1 0 372 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1712622712
transform 1 0 332 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1712622712
transform 1 0 1916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1712622712
transform 1 0 1852 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1712622712
transform 1 0 2724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1712622712
transform 1 0 1868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1712622712
transform 1 0 2828 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1712622712
transform 1 0 2692 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1712622712
transform 1 0 2692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1712622712
transform 1 0 2676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1712622712
transform 1 0 2724 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1712622712
transform 1 0 2652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1712622712
transform 1 0 2612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1712622712
transform 1 0 2540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1712622712
transform 1 0 2236 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1712622712
transform 1 0 2668 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1712622712
transform 1 0 2468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1712622712
transform 1 0 2332 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1712622712
transform 1 0 2724 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1712622712
transform 1 0 2548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1712622712
transform 1 0 2492 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1712622712
transform 1 0 1900 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1712622712
transform 1 0 1876 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1712622712
transform 1 0 2196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1712622712
transform 1 0 1956 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1712622712
transform 1 0 2412 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1712622712
transform 1 0 2316 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1712622712
transform 1 0 2180 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1712622712
transform 1 0 2212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1712622712
transform 1 0 2164 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1712622712
transform 1 0 2156 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1712622712
transform 1 0 1988 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1712622712
transform 1 0 1924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1712622712
transform 1 0 1860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1712622712
transform 1 0 1908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1712622712
transform 1 0 1828 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1712622712
transform 1 0 1748 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1712622712
transform 1 0 1996 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1712622712
transform 1 0 1532 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1712622712
transform 1 0 1556 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1712622712
transform 1 0 1284 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1712622712
transform 1 0 1260 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1712622712
transform 1 0 1220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1712622712
transform 1 0 1372 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1712622712
transform 1 0 1292 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1712622712
transform 1 0 1196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1712622712
transform 1 0 1244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1712622712
transform 1 0 1172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1712622712
transform 1 0 1124 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1712622712
transform 1 0 932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1712622712
transform 1 0 932 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1712622712
transform 1 0 2460 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1712622712
transform 1 0 2036 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1712622712
transform 1 0 2428 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1712622712
transform 1 0 2420 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1712622712
transform 1 0 2388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1712622712
transform 1 0 2476 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1712622712
transform 1 0 2180 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1712622712
transform 1 0 2092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1712622712
transform 1 0 1860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1712622712
transform 1 0 1860 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1712622712
transform 1 0 1660 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1712622712
transform 1 0 1300 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1712622712
transform 1 0 196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1712622712
transform 1 0 1316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1712622712
transform 1 0 668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1712622712
transform 1 0 1684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1712622712
transform 1 0 1324 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1712622712
transform 1 0 2012 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1712622712
transform 1 0 1708 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1712622712
transform 1 0 1732 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1712622712
transform 1 0 1732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1712622712
transform 1 0 2172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1712622712
transform 1 0 1700 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1712622712
transform 1 0 1684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1712622712
transform 1 0 1652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1712622712
transform 1 0 1620 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1712622712
transform 1 0 1612 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1712622712
transform 1 0 1740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1712622712
transform 1 0 1636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1712622712
transform 1 0 1604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1712622712
transform 1 0 1620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1712622712
transform 1 0 1516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1712622712
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1712622712
transform 1 0 1212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1712622712
transform 1 0 1084 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1712622712
transform 1 0 1052 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1712622712
transform 1 0 2116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1712622712
transform 1 0 2116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1712622712
transform 1 0 2212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1712622712
transform 1 0 2188 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1712622712
transform 1 0 2220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1712622712
transform 1 0 2180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1712622712
transform 1 0 2148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1712622712
transform 1 0 2244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1712622712
transform 1 0 2244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1712622712
transform 1 0 2188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1712622712
transform 1 0 2044 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1712622712
transform 1 0 1988 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1712622712
transform 1 0 2220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1712622712
transform 1 0 1988 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1712622712
transform 1 0 2124 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1712622712
transform 1 0 1980 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1712622712
transform 1 0 2108 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1712622712
transform 1 0 2084 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1712622712
transform 1 0 2060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1712622712
transform 1 0 1972 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1712622712
transform 1 0 1964 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1712622712
transform 1 0 2124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1712622712
transform 1 0 2100 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1712622712
transform 1 0 2012 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1712622712
transform 1 0 1956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1712622712
transform 1 0 1988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1712622712
transform 1 0 1852 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1712622712
transform 1 0 1828 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1712622712
transform 1 0 1812 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1712622712
transform 1 0 2396 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1712622712
transform 1 0 2204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1712622712
transform 1 0 2180 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1712622712
transform 1 0 2068 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1712622712
transform 1 0 2332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1712622712
transform 1 0 2236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1712622712
transform 1 0 2172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1712622712
transform 1 0 2124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1712622712
transform 1 0 2028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1712622712
transform 1 0 2052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1712622712
transform 1 0 1908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1712622712
transform 1 0 1868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1712622712
transform 1 0 636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1712622712
transform 1 0 620 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1712622712
transform 1 0 636 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1712622712
transform 1 0 300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1712622712
transform 1 0 244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1712622712
transform 1 0 116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1712622712
transform 1 0 100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1712622712
transform 1 0 268 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1712622712
transform 1 0 212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1712622712
transform 1 0 148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1712622712
transform 1 0 132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1712622712
transform 1 0 228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1712622712
transform 1 0 220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1712622712
transform 1 0 692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1712622712
transform 1 0 676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1712622712
transform 1 0 820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1712622712
transform 1 0 788 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1712622712
transform 1 0 684 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1712622712
transform 1 0 700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1712622712
transform 1 0 556 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1712622712
transform 1 0 556 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1712622712
transform 1 0 460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1712622712
transform 1 0 172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1712622712
transform 1 0 188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1712622712
transform 1 0 188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1712622712
transform 1 0 308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1712622712
transform 1 0 172 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1712622712
transform 1 0 1236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1712622712
transform 1 0 204 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1712622712
transform 1 0 116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1712622712
transform 1 0 292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1712622712
transform 1 0 284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1712622712
transform 1 0 596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1712622712
transform 1 0 492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1712622712
transform 1 0 340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1712622712
transform 1 0 164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1712622712
transform 1 0 148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1712622712
transform 1 0 148 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1712622712
transform 1 0 140 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1712622712
transform 1 0 156 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1712622712
transform 1 0 156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1712622712
transform 1 0 132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1712622712
transform 1 0 132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1712622712
transform 1 0 116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1712622712
transform 1 0 108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1712622712
transform 1 0 84 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1712622712
transform 1 0 84 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1712622712
transform 1 0 1820 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1712622712
transform 1 0 1612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1712622712
transform 1 0 1612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1712622712
transform 1 0 1452 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1712622712
transform 1 0 3204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1712622712
transform 1 0 1700 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1712622712
transform 1 0 1636 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1712622712
transform 1 0 1588 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1712622712
transform 1 0 1508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1712622712
transform 1 0 1420 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1712622712
transform 1 0 1420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1712622712
transform 1 0 900 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1712622712
transform 1 0 1428 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1712622712
transform 1 0 380 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1712622712
transform 1 0 356 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1712622712
transform 1 0 300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1712622712
transform 1 0 372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1712622712
transform 1 0 356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1712622712
transform 1 0 1052 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1712622712
transform 1 0 1012 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1712622712
transform 1 0 492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1712622712
transform 1 0 268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1712622712
transform 1 0 252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1712622712
transform 1 0 396 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1712622712
transform 1 0 340 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1712622712
transform 1 0 332 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1712622712
transform 1 0 292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1712622712
transform 1 0 412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1712622712
transform 1 0 268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1712622712
transform 1 0 268 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1712622712
transform 1 0 1644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1712622712
transform 1 0 1500 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1712622712
transform 1 0 1324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1712622712
transform 1 0 892 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1712622712
transform 1 0 548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1712622712
transform 1 0 1972 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1712622712
transform 1 0 1732 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1712622712
transform 1 0 1660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1712622712
transform 1 0 540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1712622712
transform 1 0 524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1712622712
transform 1 0 324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1712622712
transform 1 0 292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1712622712
transform 1 0 292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1712622712
transform 1 0 348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1712622712
transform 1 0 292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1712622712
transform 1 0 324 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1712622712
transform 1 0 268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1712622712
transform 1 0 356 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1712622712
transform 1 0 356 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1712622712
transform 1 0 252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1712622712
transform 1 0 284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1712622712
transform 1 0 260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1712622712
transform 1 0 252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1712622712
transform 1 0 2172 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1712622712
transform 1 0 2084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1712622712
transform 1 0 2084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1712622712
transform 1 0 668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1712622712
transform 1 0 2140 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1712622712
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1712622712
transform 1 0 1956 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1712622712
transform 1 0 868 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1712622712
transform 1 0 828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1712622712
transform 1 0 772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1712622712
transform 1 0 380 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1712622712
transform 1 0 308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1712622712
transform 1 0 284 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1712622712
transform 1 0 372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1712622712
transform 1 0 308 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1712622712
transform 1 0 228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1712622712
transform 1 0 2148 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1712622712
transform 1 0 2132 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1712622712
transform 1 0 2116 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1712622712
transform 1 0 2116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1712622712
transform 1 0 564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1712622712
transform 1 0 516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1712622712
transform 1 0 500 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3699
timestamp 1712622712
transform 1 0 988 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1712622712
transform 1 0 828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1712622712
transform 1 0 580 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3702
timestamp 1712622712
transform 1 0 540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1712622712
transform 1 0 452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1712622712
transform 1 0 428 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1712622712
transform 1 0 428 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1712622712
transform 1 0 428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3707
timestamp 1712622712
transform 1 0 460 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3708
timestamp 1712622712
transform 1 0 300 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1712622712
transform 1 0 268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1712622712
transform 1 0 996 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1712622712
transform 1 0 972 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1712622712
transform 1 0 956 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1712622712
transform 1 0 956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1712622712
transform 1 0 812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1712622712
transform 1 0 484 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1712622712
transform 1 0 484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1712622712
transform 1 0 724 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1712622712
transform 1 0 716 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1712622712
transform 1 0 708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1712622712
transform 1 0 572 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1712622712
transform 1 0 516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1712622712
transform 1 0 492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1712622712
transform 1 0 732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1712622712
transform 1 0 700 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1712622712
transform 1 0 684 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1712622712
transform 1 0 676 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1712622712
transform 1 0 564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1712622712
transform 1 0 500 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1712622712
transform 1 0 1484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1712622712
transform 1 0 1484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1712622712
transform 1 0 1932 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1712622712
transform 1 0 1724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1712622712
transform 1 0 1468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1712622712
transform 1 0 1508 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1712622712
transform 1 0 1468 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1712622712
transform 1 0 1420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1712622712
transform 1 0 1372 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1712622712
transform 1 0 1028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1712622712
transform 1 0 844 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1712622712
transform 1 0 620 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1712622712
transform 1 0 148 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1712622712
transform 1 0 140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1712622712
transform 1 0 1516 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1712622712
transform 1 0 1508 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1712622712
transform 1 0 1628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1712622712
transform 1 0 1476 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1712622712
transform 1 0 1468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1712622712
transform 1 0 1516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1712622712
transform 1 0 1452 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1712622712
transform 1 0 1380 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1712622712
transform 1 0 1468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1712622712
transform 1 0 1436 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3753
timestamp 1712622712
transform 1 0 1436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1712622712
transform 1 0 2412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1712622712
transform 1 0 1804 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1712622712
transform 1 0 1812 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1712622712
transform 1 0 1812 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1712622712
transform 1 0 1804 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1712622712
transform 1 0 1804 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1712622712
transform 1 0 1852 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1712622712
transform 1 0 1828 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1712622712
transform 1 0 1828 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1712622712
transform 1 0 1812 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1712622712
transform 1 0 1940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1712622712
transform 1 0 1812 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3766
timestamp 1712622712
transform 1 0 1844 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1712622712
transform 1 0 1348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1712622712
transform 1 0 1324 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1712622712
transform 1 0 1292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1712622712
transform 1 0 1484 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1712622712
transform 1 0 1428 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1712622712
transform 1 0 1260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1712622712
transform 1 0 1332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1712622712
transform 1 0 1164 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1712622712
transform 1 0 1156 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1712622712
transform 1 0 1836 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1712622712
transform 1 0 1820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1712622712
transform 1 0 1724 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1712622712
transform 1 0 1572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1712622712
transform 1 0 1308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1712622712
transform 1 0 1180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1712622712
transform 1 0 996 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1712622712
transform 1 0 948 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1712622712
transform 1 0 2380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3785
timestamp 1712622712
transform 1 0 1964 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1712622712
transform 1 0 2476 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1712622712
transform 1 0 2348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1712622712
transform 1 0 2348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1712622712
transform 1 0 2396 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1712622712
transform 1 0 2308 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1712622712
transform 1 0 2276 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1712622712
transform 1 0 2476 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1712622712
transform 1 0 2412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1712622712
transform 1 0 2324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1712622712
transform 1 0 2284 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1712622712
transform 1 0 1932 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1712622712
transform 1 0 2548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1712622712
transform 1 0 2532 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1712622712
transform 1 0 2532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1712622712
transform 1 0 2404 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1712622712
transform 1 0 1836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1712622712
transform 1 0 1764 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1712622712
transform 1 0 1732 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1712622712
transform 1 0 2252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1712622712
transform 1 0 1764 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1712622712
transform 1 0 1828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1712622712
transform 1 0 1772 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3808
timestamp 1712622712
transform 1 0 1860 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1712622712
transform 1 0 1820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1712622712
transform 1 0 1820 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1712622712
transform 1 0 2044 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1712622712
transform 1 0 1940 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1712622712
transform 1 0 1868 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1712622712
transform 1 0 2916 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1712622712
transform 1 0 2852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1712622712
transform 1 0 2596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1712622712
transform 1 0 2556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1712622712
transform 1 0 2436 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1712622712
transform 1 0 2044 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1712622712
transform 1 0 2004 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1712622712
transform 1 0 1908 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1712622712
transform 1 0 3044 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1712622712
transform 1 0 3036 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1712622712
transform 1 0 2900 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1712622712
transform 1 0 2492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3826
timestamp 1712622712
transform 1 0 2484 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1712622712
transform 1 0 2484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1712622712
transform 1 0 2484 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1712622712
transform 1 0 2484 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1712622712
transform 1 0 2740 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1712622712
transform 1 0 2076 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1712622712
transform 1 0 1876 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1712622712
transform 1 0 2276 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1712622712
transform 1 0 2236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1712622712
transform 1 0 2196 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1712622712
transform 1 0 2196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1712622712
transform 1 0 2468 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1712622712
transform 1 0 2356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1712622712
transform 1 0 2260 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1712622712
transform 1 0 3108 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1712622712
transform 1 0 3084 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1712622712
transform 1 0 2644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1712622712
transform 1 0 2620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1712622712
transform 1 0 2508 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1712622712
transform 1 0 2492 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1712622712
transform 1 0 2404 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1712622712
transform 1 0 2388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1712622712
transform 1 0 2364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1712622712
transform 1 0 2364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1712622712
transform 1 0 2412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1712622712
transform 1 0 2396 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1712622712
transform 1 0 2324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1712622712
transform 1 0 2300 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1712622712
transform 1 0 2268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1712622712
transform 1 0 2428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1712622712
transform 1 0 2252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1712622712
transform 1 0 2196 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1712622712
transform 1 0 2772 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1712622712
transform 1 0 2772 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1712622712
transform 1 0 2708 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1712622712
transform 1 0 2652 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1712622712
transform 1 0 3156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1712622712
transform 1 0 3044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1712622712
transform 1 0 3028 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1712622712
transform 1 0 1788 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1712622712
transform 1 0 1636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1712622712
transform 1 0 1628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1712622712
transform 1 0 132 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1712622712
transform 1 0 148 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1712622712
transform 1 0 84 0 1 1495
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1712622712
transform 1 0 132 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1712622712
transform 1 0 84 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1712622712
transform 1 0 140 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1712622712
transform 1 0 116 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1712622712
transform 1 0 716 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1712622712
transform 1 0 132 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1712622712
transform 1 0 148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1712622712
transform 1 0 132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1712622712
transform 1 0 84 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1712622712
transform 1 0 84 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1712622712
transform 1 0 84 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1712622712
transform 1 0 2140 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1712622712
transform 1 0 1676 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1712622712
transform 1 0 1276 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1712622712
transform 1 0 1276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1712622712
transform 1 0 740 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1712622712
transform 1 0 580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1712622712
transform 1 0 372 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1712622712
transform 1 0 332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1712622712
transform 1 0 332 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1712622712
transform 1 0 108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1712622712
transform 1 0 124 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1712622712
transform 1 0 116 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1712622712
transform 1 0 156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1712622712
transform 1 0 116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1712622712
transform 1 0 108 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1712622712
transform 1 0 140 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1712622712
transform 1 0 108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1712622712
transform 1 0 108 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1712622712
transform 1 0 756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1712622712
transform 1 0 732 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1712622712
transform 1 0 1004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1712622712
transform 1 0 996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3904
timestamp 1712622712
transform 1 0 748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1712622712
transform 1 0 796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1712622712
transform 1 0 796 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1712622712
transform 1 0 548 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1712622712
transform 1 0 516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1712622712
transform 1 0 148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3910
timestamp 1712622712
transform 1 0 84 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1712622712
transform 1 0 84 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1712622712
transform 1 0 156 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1712622712
transform 1 0 84 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1712622712
transform 1 0 140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1712622712
transform 1 0 140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3916
timestamp 1712622712
transform 1 0 84 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1712622712
transform 1 0 196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1712622712
transform 1 0 108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1712622712
transform 1 0 100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1712622712
transform 1 0 236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1712622712
transform 1 0 124 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1712622712
transform 1 0 540 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3923
timestamp 1712622712
transform 1 0 228 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1712622712
transform 1 0 220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3925
timestamp 1712622712
transform 1 0 252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3926
timestamp 1712622712
transform 1 0 204 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1712622712
transform 1 0 100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3928
timestamp 1712622712
transform 1 0 1188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1712622712
transform 1 0 1140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1712622712
transform 1 0 1268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1712622712
transform 1 0 1220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1712622712
transform 1 0 1460 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1712622712
transform 1 0 1364 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3934
timestamp 1712622712
transform 1 0 1244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3935
timestamp 1712622712
transform 1 0 1196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1712622712
transform 1 0 1284 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3937
timestamp 1712622712
transform 1 0 1284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1712622712
transform 1 0 1372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3939
timestamp 1712622712
transform 1 0 1372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1712622712
transform 1 0 1348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1712622712
transform 1 0 1308 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3942
timestamp 1712622712
transform 1 0 1244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3943
timestamp 1712622712
transform 1 0 1436 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1712622712
transform 1 0 1348 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1712622712
transform 1 0 1164 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3946
timestamp 1712622712
transform 1 0 1132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3947
timestamp 1712622712
transform 1 0 1620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1712622712
transform 1 0 1508 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1712622712
transform 1 0 1340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1712622712
transform 1 0 1156 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1712622712
transform 1 0 1924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3952
timestamp 1712622712
transform 1 0 1756 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1712622712
transform 1 0 1764 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1712622712
transform 1 0 1764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1712622712
transform 1 0 1908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1712622712
transform 1 0 1764 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1712622712
transform 1 0 2068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1712622712
transform 1 0 1932 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1712622712
transform 1 0 1956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1712622712
transform 1 0 1956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3961
timestamp 1712622712
transform 1 0 1932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1712622712
transform 1 0 1532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1712622712
transform 1 0 1364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3964
timestamp 1712622712
transform 1 0 2508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3965
timestamp 1712622712
transform 1 0 2444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1712622712
transform 1 0 2428 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3967
timestamp 1712622712
transform 1 0 2404 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1712622712
transform 1 0 2108 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1712622712
transform 1 0 1996 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1712622712
transform 1 0 1980 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1712622712
transform 1 0 1956 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1712622712
transform 1 0 1956 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1712622712
transform 1 0 1948 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3974
timestamp 1712622712
transform 1 0 1916 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3975
timestamp 1712622712
transform 1 0 1844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1712622712
transform 1 0 1796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1712622712
transform 1 0 1964 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1712622712
transform 1 0 1964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1712622712
transform 1 0 2108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3980
timestamp 1712622712
transform 1 0 1996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1712622712
transform 1 0 1956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3982
timestamp 1712622712
transform 1 0 1972 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1712622712
transform 1 0 1724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1712622712
transform 1 0 2964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1712622712
transform 1 0 2604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1712622712
transform 1 0 2556 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3987
timestamp 1712622712
transform 1 0 2532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1712622712
transform 1 0 2451 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1712622712
transform 1 0 2196 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1712622712
transform 1 0 2172 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1712622712
transform 1 0 2068 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1712622712
transform 1 0 2052 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1712622712
transform 1 0 2052 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1712622712
transform 1 0 2028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3995
timestamp 1712622712
transform 1 0 2180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1712622712
transform 1 0 2092 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1712622712
transform 1 0 2156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1712622712
transform 1 0 2148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1712622712
transform 1 0 2092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1712622712
transform 1 0 2084 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1712622712
transform 1 0 2188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1712622712
transform 1 0 2188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1712622712
transform 1 0 2156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1712622712
transform 1 0 2052 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1712622712
transform 1 0 2036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4006
timestamp 1712622712
transform 1 0 1724 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1712622712
transform 1 0 1604 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1712622712
transform 1 0 2244 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1712622712
transform 1 0 1740 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4010
timestamp 1712622712
transform 1 0 2220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1712622712
transform 1 0 2148 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4012
timestamp 1712622712
transform 1 0 2260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1712622712
transform 1 0 2260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1712622712
transform 1 0 1956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1712622712
transform 1 0 1740 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1712622712
transform 1 0 1588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1712622712
transform 1 0 1620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1712622712
transform 1 0 1036 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1712622712
transform 1 0 676 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1712622712
transform 1 0 644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1712622712
transform 1 0 2108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4022
timestamp 1712622712
transform 1 0 1940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1712622712
transform 1 0 1908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1712622712
transform 1 0 1948 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1712622712
transform 1 0 1908 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1712622712
transform 1 0 1932 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1712622712
transform 1 0 1804 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4028
timestamp 1712622712
transform 1 0 1804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4029
timestamp 1712622712
transform 1 0 1964 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1712622712
transform 1 0 1884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1712622712
transform 1 0 1884 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1712622712
transform 1 0 1532 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1712622712
transform 1 0 1404 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1712622712
transform 1 0 1596 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1712622712
transform 1 0 1500 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1712622712
transform 1 0 1492 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4037
timestamp 1712622712
transform 1 0 1444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1712622712
transform 1 0 1276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4039
timestamp 1712622712
transform 1 0 1164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4040
timestamp 1712622712
transform 1 0 972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4041
timestamp 1712622712
transform 1 0 956 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1712622712
transform 1 0 940 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1712622712
transform 1 0 892 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1712622712
transform 1 0 804 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1712622712
transform 1 0 540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1712622712
transform 1 0 532 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1712622712
transform 1 0 516 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1712622712
transform 1 0 508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1712622712
transform 1 0 1364 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1712622712
transform 1 0 1340 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1712622712
transform 1 0 1332 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1712622712
transform 1 0 1292 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4053
timestamp 1712622712
transform 1 0 1268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1712622712
transform 1 0 1612 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1712622712
transform 1 0 1612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4056
timestamp 1712622712
transform 1 0 3212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1712622712
transform 1 0 1572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1712622712
transform 1 0 1412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1712622712
transform 1 0 1404 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1712622712
transform 1 0 1732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1712622712
transform 1 0 1636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1712622712
transform 1 0 1300 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1712622712
transform 1 0 1236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1712622712
transform 1 0 1220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1712622712
transform 1 0 1164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1712622712
transform 1 0 1148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1712622712
transform 1 0 1124 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1712622712
transform 1 0 1268 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4069
timestamp 1712622712
transform 1 0 1236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1712622712
transform 1 0 1172 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1712622712
transform 1 0 868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1712622712
transform 1 0 1372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1712622712
transform 1 0 1332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1712622712
transform 1 0 1308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1712622712
transform 1 0 1340 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1712622712
transform 1 0 1196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4077
timestamp 1712622712
transform 1 0 1196 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4078
timestamp 1712622712
transform 1 0 1028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4079
timestamp 1712622712
transform 1 0 716 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1712622712
transform 1 0 524 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1712622712
transform 1 0 1292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4082
timestamp 1712622712
transform 1 0 956 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1712622712
transform 1 0 1364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4084
timestamp 1712622712
transform 1 0 1260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4085
timestamp 1712622712
transform 1 0 1236 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1712622712
transform 1 0 1220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4087
timestamp 1712622712
transform 1 0 1116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1712622712
transform 1 0 1100 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1712622712
transform 1 0 812 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4090
timestamp 1712622712
transform 1 0 532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1712622712
transform 1 0 412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1712622712
transform 1 0 332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4093
timestamp 1712622712
transform 1 0 332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4094
timestamp 1712622712
transform 1 0 1164 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1712622712
transform 1 0 1116 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1712622712
transform 1 0 1068 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1712622712
transform 1 0 1044 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1712622712
transform 1 0 1428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1712622712
transform 1 0 1380 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1712622712
transform 1 0 1004 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1712622712
transform 1 0 1004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4102
timestamp 1712622712
transform 1 0 788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1712622712
transform 1 0 788 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1712622712
transform 1 0 1108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1712622712
transform 1 0 780 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4106
timestamp 1712622712
transform 1 0 1412 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1712622712
transform 1 0 1084 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1712622712
transform 1 0 1164 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1712622712
transform 1 0 1092 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1712622712
transform 1 0 1196 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1712622712
transform 1 0 1196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4112
timestamp 1712622712
transform 1 0 1124 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1712622712
transform 1 0 1116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1712622712
transform 1 0 1020 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1712622712
transform 1 0 812 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1712622712
transform 1 0 372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4117
timestamp 1712622712
transform 1 0 308 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1712622712
transform 1 0 284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1712622712
transform 1 0 1180 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4120
timestamp 1712622712
transform 1 0 1172 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1712622712
transform 1 0 1116 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1712622712
transform 1 0 1068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1712622712
transform 1 0 1452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4124
timestamp 1712622712
transform 1 0 1444 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4125
timestamp 1712622712
transform 1 0 3260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4126
timestamp 1712622712
transform 1 0 3140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1712622712
transform 1 0 3068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4128
timestamp 1712622712
transform 1 0 3004 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4129
timestamp 1712622712
transform 1 0 2972 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1712622712
transform 1 0 868 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4131
timestamp 1712622712
transform 1 0 716 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4132
timestamp 1712622712
transform 1 0 1364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4133
timestamp 1712622712
transform 1 0 844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4134
timestamp 1712622712
transform 1 0 860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1712622712
transform 1 0 852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1712622712
transform 1 0 1004 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4137
timestamp 1712622712
transform 1 0 852 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4138
timestamp 1712622712
transform 1 0 868 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4139
timestamp 1712622712
transform 1 0 828 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4140
timestamp 1712622712
transform 1 0 1284 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1712622712
transform 1 0 1276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1712622712
transform 1 0 1132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4143
timestamp 1712622712
transform 1 0 964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4144
timestamp 1712622712
transform 1 0 932 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4145
timestamp 1712622712
transform 1 0 932 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4146
timestamp 1712622712
transform 1 0 860 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4147
timestamp 1712622712
transform 1 0 1244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4148
timestamp 1712622712
transform 1 0 1188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1712622712
transform 1 0 1204 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4150
timestamp 1712622712
transform 1 0 1188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4151
timestamp 1712622712
transform 1 0 2876 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4152
timestamp 1712622712
transform 1 0 2852 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1712622712
transform 1 0 2308 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4154
timestamp 1712622712
transform 1 0 1468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4155
timestamp 1712622712
transform 1 0 1340 0 1 1285
box -2 -2 2 2
use M2_M1  M2_M1_4156
timestamp 1712622712
transform 1 0 1316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4157
timestamp 1712622712
transform 1 0 1308 0 1 1285
box -2 -2 2 2
use M2_M1  M2_M1_4158
timestamp 1712622712
transform 1 0 1308 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4159
timestamp 1712622712
transform 1 0 1252 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4160
timestamp 1712622712
transform 1 0 1212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4161
timestamp 1712622712
transform 1 0 3004 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1712622712
transform 1 0 2900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4163
timestamp 1712622712
transform 1 0 1660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4164
timestamp 1712622712
transform 1 0 1348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4165
timestamp 1712622712
transform 1 0 1324 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4166
timestamp 1712622712
transform 1 0 1268 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4167
timestamp 1712622712
transform 1 0 1228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4168
timestamp 1712622712
transform 1 0 1220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4169
timestamp 1712622712
transform 1 0 1348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4170
timestamp 1712622712
transform 1 0 1324 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4171
timestamp 1712622712
transform 1 0 1412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4172
timestamp 1712622712
transform 1 0 1404 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4173
timestamp 1712622712
transform 1 0 1420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1712622712
transform 1 0 1348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4175
timestamp 1712622712
transform 1 0 1356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4176
timestamp 1712622712
transform 1 0 1356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4177
timestamp 1712622712
transform 1 0 1132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4178
timestamp 1712622712
transform 1 0 1132 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4179
timestamp 1712622712
transform 1 0 1076 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4180
timestamp 1712622712
transform 1 0 1068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4181
timestamp 1712622712
transform 1 0 996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4182
timestamp 1712622712
transform 1 0 908 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4183
timestamp 1712622712
transform 1 0 1540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4184
timestamp 1712622712
transform 1 0 1436 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4185
timestamp 1712622712
transform 1 0 612 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4186
timestamp 1712622712
transform 1 0 516 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4187
timestamp 1712622712
transform 1 0 588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4188
timestamp 1712622712
transform 1 0 588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4189
timestamp 1712622712
transform 1 0 812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4190
timestamp 1712622712
transform 1 0 596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4191
timestamp 1712622712
transform 1 0 932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4192
timestamp 1712622712
transform 1 0 788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4193
timestamp 1712622712
transform 1 0 804 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1712622712
transform 1 0 740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4195
timestamp 1712622712
transform 1 0 1132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4196
timestamp 1712622712
transform 1 0 1100 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1712622712
transform 1 0 980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1712622712
transform 1 0 940 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4199
timestamp 1712622712
transform 1 0 748 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1712622712
transform 1 0 740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1712622712
transform 1 0 740 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4202
timestamp 1712622712
transform 1 0 308 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4203
timestamp 1712622712
transform 1 0 300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4204
timestamp 1712622712
transform 1 0 236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4205
timestamp 1712622712
transform 1 0 884 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1712622712
transform 1 0 756 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4207
timestamp 1712622712
transform 1 0 756 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4208
timestamp 1712622712
transform 1 0 1244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4209
timestamp 1712622712
transform 1 0 1116 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4210
timestamp 1712622712
transform 1 0 1156 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4211
timestamp 1712622712
transform 1 0 1132 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4212
timestamp 1712622712
transform 1 0 1572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4213
timestamp 1712622712
transform 1 0 1556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1712622712
transform 1 0 1268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4215
timestamp 1712622712
transform 1 0 1196 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4216
timestamp 1712622712
transform 1 0 940 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4217
timestamp 1712622712
transform 1 0 1228 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1712622712
transform 1 0 1188 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4219
timestamp 1712622712
transform 1 0 2820 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4220
timestamp 1712622712
transform 1 0 2788 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4221
timestamp 1712622712
transform 1 0 2708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1712622712
transform 1 0 1684 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1712622712
transform 1 0 1628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4224
timestamp 1712622712
transform 1 0 1364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4225
timestamp 1712622712
transform 1 0 1276 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4226
timestamp 1712622712
transform 1 0 972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1712622712
transform 1 0 588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1712622712
transform 1 0 588 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4229
timestamp 1712622712
transform 1 0 668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1712622712
transform 1 0 628 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4231
timestamp 1712622712
transform 1 0 2964 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1712622712
transform 1 0 2500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4233
timestamp 1712622712
transform 1 0 1196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1712622712
transform 1 0 868 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1712622712
transform 1 0 812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4236
timestamp 1712622712
transform 1 0 1092 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1712622712
transform 1 0 1044 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1712622712
transform 1 0 980 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4239
timestamp 1712622712
transform 1 0 1628 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4240
timestamp 1712622712
transform 1 0 1580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4241
timestamp 1712622712
transform 1 0 1044 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4242
timestamp 1712622712
transform 1 0 916 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4243
timestamp 1712622712
transform 1 0 1268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4244
timestamp 1712622712
transform 1 0 1052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4245
timestamp 1712622712
transform 1 0 436 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4246
timestamp 1712622712
transform 1 0 436 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4247
timestamp 1712622712
transform 1 0 428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1712622712
transform 1 0 396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1712622712
transform 1 0 676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1712622712
transform 1 0 444 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4251
timestamp 1712622712
transform 1 0 476 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4252
timestamp 1712622712
transform 1 0 468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1712622712
transform 1 0 1244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4254
timestamp 1712622712
transform 1 0 700 0 1 1814
box -2 -2 2 2
use M2_M1  M2_M1_4255
timestamp 1712622712
transform 1 0 692 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_4256
timestamp 1712622712
transform 1 0 668 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_4257
timestamp 1712622712
transform 1 0 588 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4258
timestamp 1712622712
transform 1 0 572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4259
timestamp 1712622712
transform 1 0 548 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1712622712
transform 1 0 548 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_4261
timestamp 1712622712
transform 1 0 524 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1712622712
transform 1 0 524 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1712622712
transform 1 0 468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4264
timestamp 1712622712
transform 1 0 452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4265
timestamp 1712622712
transform 1 0 412 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4266
timestamp 1712622712
transform 1 0 316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4267
timestamp 1712622712
transform 1 0 276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4268
timestamp 1712622712
transform 1 0 652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1712622712
transform 1 0 572 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4270
timestamp 1712622712
transform 1 0 468 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4271
timestamp 1712622712
transform 1 0 708 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4272
timestamp 1712622712
transform 1 0 508 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4273
timestamp 1712622712
transform 1 0 508 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4274
timestamp 1712622712
transform 1 0 380 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1712622712
transform 1 0 372 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4276
timestamp 1712622712
transform 1 0 780 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1712622712
transform 1 0 692 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_4278
timestamp 1712622712
transform 1 0 700 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4279
timestamp 1712622712
transform 1 0 668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1712622712
transform 1 0 324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4281
timestamp 1712622712
transform 1 0 196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4282
timestamp 1712622712
transform 1 0 1980 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1712622712
transform 1 0 1300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4284
timestamp 1712622712
transform 1 0 740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4285
timestamp 1712622712
transform 1 0 708 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1712622712
transform 1 0 2892 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4287
timestamp 1712622712
transform 1 0 2836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4288
timestamp 1712622712
transform 1 0 1868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4289
timestamp 1712622712
transform 1 0 1740 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4290
timestamp 1712622712
transform 1 0 1500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4291
timestamp 1712622712
transform 1 0 996 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4292
timestamp 1712622712
transform 1 0 996 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1712622712
transform 1 0 308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4294
timestamp 1712622712
transform 1 0 284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1712622712
transform 1 0 396 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1712622712
transform 1 0 380 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4297
timestamp 1712622712
transform 1 0 2908 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4298
timestamp 1712622712
transform 1 0 2252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4299
timestamp 1712622712
transform 1 0 1252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1712622712
transform 1 0 636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4301
timestamp 1712622712
transform 1 0 604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1712622712
transform 1 0 2036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4303
timestamp 1712622712
transform 1 0 1396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1712622712
transform 1 0 676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1712622712
transform 1 0 652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1712622712
transform 1 0 1100 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4307
timestamp 1712622712
transform 1 0 980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1712622712
transform 1 0 964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4309
timestamp 1712622712
transform 1 0 836 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4310
timestamp 1712622712
transform 1 0 724 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1712622712
transform 1 0 716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4312
timestamp 1712622712
transform 1 0 2748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1712622712
transform 1 0 1356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1712622712
transform 1 0 1356 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1712622712
transform 1 0 1340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4316
timestamp 1712622712
transform 1 0 1284 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1712622712
transform 1 0 1268 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4318
timestamp 1712622712
transform 1 0 1244 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4319
timestamp 1712622712
transform 1 0 1180 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4320
timestamp 1712622712
transform 1 0 1140 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1712622712
transform 1 0 1140 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4322
timestamp 1712622712
transform 1 0 1124 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4323
timestamp 1712622712
transform 1 0 340 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4324
timestamp 1712622712
transform 1 0 340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4325
timestamp 1712622712
transform 1 0 260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4326
timestamp 1712622712
transform 1 0 188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4327
timestamp 1712622712
transform 1 0 332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4328
timestamp 1712622712
transform 1 0 292 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1712622712
transform 1 0 580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1712622712
transform 1 0 356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4331
timestamp 1712622712
transform 1 0 388 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1712622712
transform 1 0 380 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1712622712
transform 1 0 924 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4334
timestamp 1712622712
transform 1 0 372 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1712622712
transform 1 0 356 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1712622712
transform 1 0 996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1712622712
transform 1 0 340 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4338
timestamp 1712622712
transform 1 0 268 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1712622712
transform 1 0 212 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1712622712
transform 1 0 108 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4341
timestamp 1712622712
transform 1 0 1036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4342
timestamp 1712622712
transform 1 0 628 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4343
timestamp 1712622712
transform 1 0 628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4344
timestamp 1712622712
transform 1 0 628 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4345
timestamp 1712622712
transform 1 0 148 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4346
timestamp 1712622712
transform 1 0 68 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4347
timestamp 1712622712
transform 1 0 1988 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4348
timestamp 1712622712
transform 1 0 1556 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4349
timestamp 1712622712
transform 1 0 1020 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1712622712
transform 1 0 1004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4351
timestamp 1712622712
transform 1 0 1068 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4352
timestamp 1712622712
transform 1 0 1036 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4353
timestamp 1712622712
transform 1 0 124 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1712622712
transform 1 0 108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4355
timestamp 1712622712
transform 1 0 228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4356
timestamp 1712622712
transform 1 0 196 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4357
timestamp 1712622712
transform 1 0 2812 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4358
timestamp 1712622712
transform 1 0 2388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4359
timestamp 1712622712
transform 1 0 1580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4360
timestamp 1712622712
transform 1 0 900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4361
timestamp 1712622712
transform 1 0 876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4362
timestamp 1712622712
transform 1 0 1900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4363
timestamp 1712622712
transform 1 0 1700 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4364
timestamp 1712622712
transform 1 0 964 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4365
timestamp 1712622712
transform 1 0 924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4366
timestamp 1712622712
transform 1 0 1068 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4367
timestamp 1712622712
transform 1 0 1044 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4368
timestamp 1712622712
transform 1 0 924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1712622712
transform 1 0 876 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1712622712
transform 1 0 572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1712622712
transform 1 0 556 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_4372
timestamp 1712622712
transform 1 0 292 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1712622712
transform 1 0 276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4374
timestamp 1712622712
transform 1 0 252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4375
timestamp 1712622712
transform 1 0 252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1712622712
transform 1 0 572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1712622712
transform 1 0 292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4378
timestamp 1712622712
transform 1 0 436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4379
timestamp 1712622712
transform 1 0 308 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1712622712
transform 1 0 1228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1712622712
transform 1 0 732 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4382
timestamp 1712622712
transform 1 0 604 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_4383
timestamp 1712622712
transform 1 0 364 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4384
timestamp 1712622712
transform 1 0 364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4385
timestamp 1712622712
transform 1 0 332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4386
timestamp 1712622712
transform 1 0 316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4387
timestamp 1712622712
transform 1 0 316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4388
timestamp 1712622712
transform 1 0 308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4389
timestamp 1712622712
transform 1 0 300 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4390
timestamp 1712622712
transform 1 0 804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4391
timestamp 1712622712
transform 1 0 364 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4392
timestamp 1712622712
transform 1 0 356 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4393
timestamp 1712622712
transform 1 0 1004 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4394
timestamp 1712622712
transform 1 0 356 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_4395
timestamp 1712622712
transform 1 0 268 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1712622712
transform 1 0 188 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_4397
timestamp 1712622712
transform 1 0 132 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4398
timestamp 1712622712
transform 1 0 892 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4399
timestamp 1712622712
transform 1 0 596 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4400
timestamp 1712622712
transform 1 0 620 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1712622712
transform 1 0 572 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1712622712
transform 1 0 132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1712622712
transform 1 0 116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4404
timestamp 1712622712
transform 1 0 900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1712622712
transform 1 0 884 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4406
timestamp 1712622712
transform 1 0 188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4407
timestamp 1712622712
transform 1 0 116 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4408
timestamp 1712622712
transform 1 0 284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4409
timestamp 1712622712
transform 1 0 236 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4410
timestamp 1712622712
transform 1 0 1156 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4411
timestamp 1712622712
transform 1 0 820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4412
timestamp 1712622712
transform 1 0 1172 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4413
timestamp 1712622712
transform 1 0 1148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4414
timestamp 1712622712
transform 1 0 1076 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4415
timestamp 1712622712
transform 1 0 1076 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4416
timestamp 1712622712
transform 1 0 1004 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4417
timestamp 1712622712
transform 1 0 892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4418
timestamp 1712622712
transform 1 0 708 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4419
timestamp 1712622712
transform 1 0 1164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4420
timestamp 1712622712
transform 1 0 980 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4421
timestamp 1712622712
transform 1 0 1124 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1712622712
transform 1 0 980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4423
timestamp 1712622712
transform 1 0 1100 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4424
timestamp 1712622712
transform 1 0 1100 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1712622712
transform 1 0 940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4426
timestamp 1712622712
transform 1 0 916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1712622712
transform 1 0 916 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4428
timestamp 1712622712
transform 1 0 900 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1712622712
transform 1 0 900 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4430
timestamp 1712622712
transform 1 0 876 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4431
timestamp 1712622712
transform 1 0 644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4432
timestamp 1712622712
transform 1 0 1068 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1712622712
transform 1 0 1044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4434
timestamp 1712622712
transform 1 0 1748 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4435
timestamp 1712622712
transform 1 0 1380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4436
timestamp 1712622712
transform 1 0 1244 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1712622712
transform 1 0 1140 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4438
timestamp 1712622712
transform 1 0 268 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4439
timestamp 1712622712
transform 1 0 236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4440
timestamp 1712622712
transform 1 0 212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4441
timestamp 1712622712
transform 1 0 212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4442
timestamp 1712622712
transform 1 0 356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4443
timestamp 1712622712
transform 1 0 220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1712622712
transform 1 0 572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1712622712
transform 1 0 356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4446
timestamp 1712622712
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4447
timestamp 1712622712
transform 1 0 412 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1712622712
transform 1 0 708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4449
timestamp 1712622712
transform 1 0 500 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4450
timestamp 1712622712
transform 1 0 452 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4451
timestamp 1712622712
transform 1 0 1204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1712622712
transform 1 0 692 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_4453
timestamp 1712622712
transform 1 0 620 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1712622712
transform 1 0 420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4455
timestamp 1712622712
transform 1 0 396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1712622712
transform 1 0 324 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4457
timestamp 1712622712
transform 1 0 244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4458
timestamp 1712622712
transform 1 0 228 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4459
timestamp 1712622712
transform 1 0 196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4460
timestamp 1712622712
transform 1 0 724 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4461
timestamp 1712622712
transform 1 0 596 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4462
timestamp 1712622712
transform 1 0 836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1712622712
transform 1 0 772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1712622712
transform 1 0 732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1712622712
transform 1 0 692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4466
timestamp 1712622712
transform 1 0 212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4467
timestamp 1712622712
transform 1 0 116 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4468
timestamp 1712622712
transform 1 0 260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4469
timestamp 1712622712
transform 1 0 236 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4470
timestamp 1712622712
transform 1 0 748 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4471
timestamp 1712622712
transform 1 0 732 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1712622712
transform 1 0 820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1712622712
transform 1 0 308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4474
timestamp 1712622712
transform 1 0 916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1712622712
transform 1 0 796 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4476
timestamp 1712622712
transform 1 0 828 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1712622712
transform 1 0 820 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4478
timestamp 1712622712
transform 1 0 836 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4479
timestamp 1712622712
transform 1 0 820 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_4480
timestamp 1712622712
transform 1 0 908 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1712622712
transform 1 0 900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4482
timestamp 1712622712
transform 1 0 900 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4483
timestamp 1712622712
transform 1 0 852 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1712622712
transform 1 0 628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4485
timestamp 1712622712
transform 1 0 1036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1712622712
transform 1 0 924 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1712622712
transform 1 0 2820 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4488
timestamp 1712622712
transform 1 0 2772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4489
timestamp 1712622712
transform 1 0 1916 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1712622712
transform 1 0 1772 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1712622712
transform 1 0 1564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4492
timestamp 1712622712
transform 1 0 1388 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_4493
timestamp 1712622712
transform 1 0 1276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4494
timestamp 1712622712
transform 1 0 1172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1712622712
transform 1 0 172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1712622712
transform 1 0 132 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4497
timestamp 1712622712
transform 1 0 140 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4498
timestamp 1712622712
transform 1 0 140 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4499
timestamp 1712622712
transform 1 0 420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1712622712
transform 1 0 156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1712622712
transform 1 0 564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4502
timestamp 1712622712
transform 1 0 452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1712622712
transform 1 0 476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4504
timestamp 1712622712
transform 1 0 468 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4505
timestamp 1712622712
transform 1 0 668 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4506
timestamp 1712622712
transform 1 0 628 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4507
timestamp 1712622712
transform 1 0 692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4508
timestamp 1712622712
transform 1 0 660 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4509
timestamp 1712622712
transform 1 0 660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4510
timestamp 1712622712
transform 1 0 620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4511
timestamp 1712622712
transform 1 0 140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4512
timestamp 1712622712
transform 1 0 108 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4513
timestamp 1712622712
transform 1 0 260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1712622712
transform 1 0 188 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4515
timestamp 1712622712
transform 1 0 652 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1712622712
transform 1 0 452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1712622712
transform 1 0 716 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4518
timestamp 1712622712
transform 1 0 684 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4519
timestamp 1712622712
transform 1 0 748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4520
timestamp 1712622712
transform 1 0 172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1712622712
transform 1 0 164 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1712622712
transform 1 0 852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1712622712
transform 1 0 716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4524
timestamp 1712622712
transform 1 0 812 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4525
timestamp 1712622712
transform 1 0 756 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1712622712
transform 1 0 860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1712622712
transform 1 0 804 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1712622712
transform 1 0 956 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4529
timestamp 1712622712
transform 1 0 892 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4530
timestamp 1712622712
transform 1 0 756 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4531
timestamp 1712622712
transform 1 0 756 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1712622712
transform 1 0 756 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1712622712
transform 1 0 748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1712622712
transform 1 0 740 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4535
timestamp 1712622712
transform 1 0 740 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_4536
timestamp 1712622712
transform 1 0 948 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4537
timestamp 1712622712
transform 1 0 852 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_4538
timestamp 1712622712
transform 1 0 180 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4539
timestamp 1712622712
transform 1 0 180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4540
timestamp 1712622712
transform 1 0 140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4541
timestamp 1712622712
transform 1 0 132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1712622712
transform 1 0 276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4543
timestamp 1712622712
transform 1 0 116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4544
timestamp 1712622712
transform 1 0 532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4545
timestamp 1712622712
transform 1 0 292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1712622712
transform 1 0 428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4547
timestamp 1712622712
transform 1 0 324 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4548
timestamp 1712622712
transform 1 0 620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1712622712
transform 1 0 476 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4550
timestamp 1712622712
transform 1 0 388 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1712622712
transform 1 0 1100 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4552
timestamp 1712622712
transform 1 0 1100 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4553
timestamp 1712622712
transform 1 0 1076 0 1 555
box -2 -2 2 2
use M2_M1  M2_M1_4554
timestamp 1712622712
transform 1 0 1004 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4555
timestamp 1712622712
transform 1 0 980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4556
timestamp 1712622712
transform 1 0 900 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4557
timestamp 1712622712
transform 1 0 460 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4558
timestamp 1712622712
transform 1 0 284 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4559
timestamp 1712622712
transform 1 0 276 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4560
timestamp 1712622712
transform 1 0 252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4561
timestamp 1712622712
transform 1 0 724 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4562
timestamp 1712622712
transform 1 0 460 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4563
timestamp 1712622712
transform 1 0 804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1712622712
transform 1 0 732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4565
timestamp 1712622712
transform 1 0 588 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4566
timestamp 1712622712
transform 1 0 588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1712622712
transform 1 0 124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4568
timestamp 1712622712
transform 1 0 100 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1712622712
transform 1 0 204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4570
timestamp 1712622712
transform 1 0 116 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1712622712
transform 1 0 660 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4572
timestamp 1712622712
transform 1 0 644 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1712622712
transform 1 0 852 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4574
timestamp 1712622712
transform 1 0 116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4575
timestamp 1712622712
transform 1 0 116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4576
timestamp 1712622712
transform 1 0 852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4577
timestamp 1712622712
transform 1 0 780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1712622712
transform 1 0 892 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1712622712
transform 1 0 836 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1712622712
transform 1 0 892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1712622712
transform 1 0 868 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4582
timestamp 1712622712
transform 1 0 1324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1712622712
transform 1 0 1236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4584
timestamp 1712622712
transform 1 0 1140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4585
timestamp 1712622712
transform 1 0 1068 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4586
timestamp 1712622712
transform 1 0 1052 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4587
timestamp 1712622712
transform 1 0 1020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4588
timestamp 1712622712
transform 1 0 940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4589
timestamp 1712622712
transform 1 0 868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4590
timestamp 1712622712
transform 1 0 948 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4591
timestamp 1712622712
transform 1 0 868 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1712622712
transform 1 0 2932 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4593
timestamp 1712622712
transform 1 0 2900 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4594
timestamp 1712622712
transform 1 0 2676 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4595
timestamp 1712622712
transform 1 0 2364 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4596
timestamp 1712622712
transform 1 0 2364 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4597
timestamp 1712622712
transform 1 0 2348 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1712622712
transform 1 0 1292 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4599
timestamp 1712622712
transform 1 0 1284 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1712622712
transform 1 0 1124 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4601
timestamp 1712622712
transform 1 0 548 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4602
timestamp 1712622712
transform 1 0 244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4603
timestamp 1712622712
transform 1 0 212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4604
timestamp 1712622712
transform 1 0 188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1712622712
transform 1 0 524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4606
timestamp 1712622712
transform 1 0 228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4607
timestamp 1712622712
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1712622712
transform 1 0 548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4609
timestamp 1712622712
transform 1 0 564 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4610
timestamp 1712622712
transform 1 0 500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1712622712
transform 1 0 1356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4612
timestamp 1712622712
transform 1 0 1356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1712622712
transform 1 0 1148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4614
timestamp 1712622712
transform 1 0 1060 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4615
timestamp 1712622712
transform 1 0 652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4616
timestamp 1712622712
transform 1 0 436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4617
timestamp 1712622712
transform 1 0 404 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1712622712
transform 1 0 396 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4619
timestamp 1712622712
transform 1 0 356 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1712622712
transform 1 0 644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1712622712
transform 1 0 452 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4622
timestamp 1712622712
transform 1 0 380 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4623
timestamp 1712622712
transform 1 0 980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4624
timestamp 1712622712
transform 1 0 380 0 1 695
box -2 -2 2 2
use M2_M1  M2_M1_4625
timestamp 1712622712
transform 1 0 372 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4626
timestamp 1712622712
transform 1 0 372 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_4627
timestamp 1712622712
transform 1 0 348 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_4628
timestamp 1712622712
transform 1 0 156 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1712622712
transform 1 0 140 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4630
timestamp 1712622712
transform 1 0 844 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4631
timestamp 1712622712
transform 1 0 652 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4632
timestamp 1712622712
transform 1 0 860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1712622712
transform 1 0 828 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_4634
timestamp 1712622712
transform 1 0 116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4635
timestamp 1712622712
transform 1 0 116 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4636
timestamp 1712622712
transform 1 0 220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4637
timestamp 1712622712
transform 1 0 196 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1712622712
transform 1 0 1108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4639
timestamp 1712622712
transform 1 0 668 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4640
timestamp 1712622712
transform 1 0 1412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4641
timestamp 1712622712
transform 1 0 1300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4642
timestamp 1712622712
transform 1 0 1148 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_4643
timestamp 1712622712
transform 1 0 1148 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1712622712
transform 1 0 1132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1712622712
transform 1 0 1044 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4646
timestamp 1712622712
transform 1 0 1004 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4647
timestamp 1712622712
transform 1 0 1324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4648
timestamp 1712622712
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4649
timestamp 1712622712
transform 1 0 988 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4650
timestamp 1712622712
transform 1 0 964 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4651
timestamp 1712622712
transform 1 0 1052 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4652
timestamp 1712622712
transform 1 0 972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4653
timestamp 1712622712
transform 1 0 1716 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1712622712
transform 1 0 1556 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1712622712
transform 1 0 1348 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1712622712
transform 1 0 1020 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4657
timestamp 1712622712
transform 1 0 1060 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1712622712
transform 1 0 1052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4659
timestamp 1712622712
transform 1 0 2932 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1712622712
transform 1 0 2916 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4661
timestamp 1712622712
transform 1 0 2876 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4662
timestamp 1712622712
transform 1 0 2436 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4663
timestamp 1712622712
transform 1 0 1716 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4664
timestamp 1712622712
transform 1 0 1412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1712622712
transform 1 0 1356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4666
timestamp 1712622712
transform 1 0 1244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4667
timestamp 1712622712
transform 1 0 1020 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4668
timestamp 1712622712
transform 1 0 2740 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1712622712
transform 1 0 2740 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4670
timestamp 1712622712
transform 1 0 2668 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4671
timestamp 1712622712
transform 1 0 2596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4672
timestamp 1712622712
transform 1 0 1828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1712622712
transform 1 0 1468 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1712622712
transform 1 0 1388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4675
timestamp 1712622712
transform 1 0 988 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4676
timestamp 1712622712
transform 1 0 228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4677
timestamp 1712622712
transform 1 0 180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1712622712
transform 1 0 180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4679
timestamp 1712622712
transform 1 0 228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4680
timestamp 1712622712
transform 1 0 212 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1712622712
transform 1 0 796 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4682
timestamp 1712622712
transform 1 0 244 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4683
timestamp 1712622712
transform 1 0 452 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4684
timestamp 1712622712
transform 1 0 300 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4685
timestamp 1712622712
transform 1 0 828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1712622712
transform 1 0 364 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1712622712
transform 1 0 348 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4688
timestamp 1712622712
transform 1 0 972 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4689
timestamp 1712622712
transform 1 0 516 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1712622712
transform 1 0 276 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_4691
timestamp 1712622712
transform 1 0 196 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4692
timestamp 1712622712
transform 1 0 196 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4693
timestamp 1712622712
transform 1 0 1036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4694
timestamp 1712622712
transform 1 0 980 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4695
timestamp 1712622712
transform 1 0 844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1712622712
transform 1 0 836 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1712622712
transform 1 0 836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1712622712
transform 1 0 964 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4699
timestamp 1712622712
transform 1 0 716 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4700
timestamp 1712622712
transform 1 0 964 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4701
timestamp 1712622712
transform 1 0 940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4702
timestamp 1712622712
transform 1 0 124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4703
timestamp 1712622712
transform 1 0 124 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1712622712
transform 1 0 252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1712622712
transform 1 0 228 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1712622712
transform 1 0 1172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4707
timestamp 1712622712
transform 1 0 956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1712622712
transform 1 0 1172 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4709
timestamp 1712622712
transform 1 0 1140 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1712622712
transform 1 0 2868 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4711
timestamp 1712622712
transform 1 0 2844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4712
timestamp 1712622712
transform 1 0 2524 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1712622712
transform 1 0 2492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1712622712
transform 1 0 2468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1712622712
transform 1 0 1788 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4716
timestamp 1712622712
transform 1 0 1524 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4717
timestamp 1712622712
transform 1 0 1396 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1712622712
transform 1 0 1108 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1712622712
transform 1 0 1124 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4720
timestamp 1712622712
transform 1 0 692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1712622712
transform 1 0 660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1712622712
transform 1 0 436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1712622712
transform 1 0 684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4724
timestamp 1712622712
transform 1 0 644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4725
timestamp 1712622712
transform 1 0 660 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1712622712
transform 1 0 532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1712622712
transform 1 0 628 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1712622712
transform 1 0 620 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1712622712
transform 1 0 596 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1712622712
transform 1 0 500 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4731
timestamp 1712622712
transform 1 0 708 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4732
timestamp 1712622712
transform 1 0 588 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4733
timestamp 1712622712
transform 1 0 588 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1712622712
transform 1 0 364 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4735
timestamp 1712622712
transform 1 0 348 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4736
timestamp 1712622712
transform 1 0 1244 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1712622712
transform 1 0 748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4738
timestamp 1712622712
transform 1 0 692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4739
timestamp 1712622712
transform 1 0 676 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1712622712
transform 1 0 644 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4741
timestamp 1712622712
transform 1 0 740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1712622712
transform 1 0 732 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1712622712
transform 1 0 524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4744
timestamp 1712622712
transform 1 0 412 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4745
timestamp 1712622712
transform 1 0 428 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1712622712
transform 1 0 340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4747
timestamp 1712622712
transform 1 0 1556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4748
timestamp 1712622712
transform 1 0 1548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4749
timestamp 1712622712
transform 1 0 1492 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4750
timestamp 1712622712
transform 1 0 1260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1712622712
transform 1 0 1260 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4752
timestamp 1712622712
transform 1 0 1196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1712622712
transform 1 0 2684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1712622712
transform 1 0 2404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1712622712
transform 1 0 1332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4756
timestamp 1712622712
transform 1 0 1268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4757
timestamp 1712622712
transform 1 0 1220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1712622712
transform 1 0 1204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4759
timestamp 1712622712
transform 1 0 1188 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4760
timestamp 1712622712
transform 1 0 1084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4761
timestamp 1712622712
transform 1 0 1084 0 1 555
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1712622712
transform 1 0 1052 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4763
timestamp 1712622712
transform 1 0 1332 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4764
timestamp 1712622712
transform 1 0 860 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1712622712
transform 1 0 804 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4766
timestamp 1712622712
transform 1 0 804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4767
timestamp 1712622712
transform 1 0 892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4768
timestamp 1712622712
transform 1 0 820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4769
timestamp 1712622712
transform 1 0 980 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4770
timestamp 1712622712
transform 1 0 908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4771
timestamp 1712622712
transform 1 0 940 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1712622712
transform 1 0 940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4773
timestamp 1712622712
transform 1 0 2404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1712622712
transform 1 0 2404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4775
timestamp 1712622712
transform 1 0 2364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4776
timestamp 1712622712
transform 1 0 2236 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4777
timestamp 1712622712
transform 1 0 1476 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1712622712
transform 1 0 988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4779
timestamp 1712622712
transform 1 0 972 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4780
timestamp 1712622712
transform 1 0 900 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4781
timestamp 1712622712
transform 1 0 852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4782
timestamp 1712622712
transform 1 0 588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1712622712
transform 1 0 908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4784
timestamp 1712622712
transform 1 0 900 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1712622712
transform 1 0 892 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4786
timestamp 1712622712
transform 1 0 948 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4787
timestamp 1712622712
transform 1 0 940 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4788
timestamp 1712622712
transform 1 0 908 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1712622712
transform 1 0 836 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4790
timestamp 1712622712
transform 1 0 772 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4791
timestamp 1712622712
transform 1 0 1284 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4792
timestamp 1712622712
transform 1 0 1116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4793
timestamp 1712622712
transform 1 0 988 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1712622712
transform 1 0 948 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4795
timestamp 1712622712
transform 1 0 916 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4796
timestamp 1712622712
transform 1 0 1044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1712622712
transform 1 0 988 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1712622712
transform 1 0 812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4799
timestamp 1712622712
transform 1 0 812 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_4800
timestamp 1712622712
transform 1 0 884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4801
timestamp 1712622712
transform 1 0 860 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4802
timestamp 1712622712
transform 1 0 1852 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4803
timestamp 1712622712
transform 1 0 1692 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_4804
timestamp 1712622712
transform 1 0 1596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4805
timestamp 1712622712
transform 1 0 1332 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4806
timestamp 1712622712
transform 1 0 1332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4807
timestamp 1712622712
transform 1 0 1252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4808
timestamp 1712622712
transform 1 0 1452 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4809
timestamp 1712622712
transform 1 0 1156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4810
timestamp 1712622712
transform 1 0 1124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4811
timestamp 1712622712
transform 1 0 1124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4812
timestamp 1712622712
transform 1 0 1156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4813
timestamp 1712622712
transform 1 0 1140 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4814
timestamp 1712622712
transform 1 0 1164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4815
timestamp 1712622712
transform 1 0 1148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4816
timestamp 1712622712
transform 1 0 1180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1712622712
transform 1 0 1180 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4818
timestamp 1712622712
transform 1 0 1140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4819
timestamp 1712622712
transform 1 0 1060 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1712622712
transform 1 0 1060 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4821
timestamp 1712622712
transform 1 0 1172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4822
timestamp 1712622712
transform 1 0 1132 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4823
timestamp 1712622712
transform 1 0 1124 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4824
timestamp 1712622712
transform 1 0 1076 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4825
timestamp 1712622712
transform 1 0 1076 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_4826
timestamp 1712622712
transform 1 0 1044 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4827
timestamp 1712622712
transform 1 0 1180 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4828
timestamp 1712622712
transform 1 0 1044 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4829
timestamp 1712622712
transform 1 0 1164 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4830
timestamp 1712622712
transform 1 0 1140 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1712622712
transform 1 0 1060 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1712622712
transform 1 0 1044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4833
timestamp 1712622712
transform 1 0 1116 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4834
timestamp 1712622712
transform 1 0 1100 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4835
timestamp 1712622712
transform 1 0 1196 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1712622712
transform 1 0 1156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1712622712
transform 1 0 1724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4838
timestamp 1712622712
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4839
timestamp 1712622712
transform 1 0 1524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4840
timestamp 1712622712
transform 1 0 1428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4841
timestamp 1712622712
transform 1 0 1388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4842
timestamp 1712622712
transform 1 0 1212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4843
timestamp 1712622712
transform 1 0 1196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4844
timestamp 1712622712
transform 1 0 1180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4845
timestamp 1712622712
transform 1 0 1148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4846
timestamp 1712622712
transform 1 0 1220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4847
timestamp 1712622712
transform 1 0 1156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4848
timestamp 1712622712
transform 1 0 2004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4849
timestamp 1712622712
transform 1 0 1908 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4850
timestamp 1712622712
transform 1 0 1724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1712622712
transform 1 0 1708 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4852
timestamp 1712622712
transform 1 0 1668 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4853
timestamp 1712622712
transform 1 0 1668 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4854
timestamp 1712622712
transform 1 0 1492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4855
timestamp 1712622712
transform 1 0 1420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1712622712
transform 1 0 1412 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4857
timestamp 1712622712
transform 1 0 1180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4858
timestamp 1712622712
transform 1 0 1076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1712622712
transform 1 0 1516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4860
timestamp 1712622712
transform 1 0 1484 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1712622712
transform 1 0 1492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4862
timestamp 1712622712
transform 1 0 1492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4863
timestamp 1712622712
transform 1 0 1476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4864
timestamp 1712622712
transform 1 0 1468 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4865
timestamp 1712622712
transform 1 0 1484 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4866
timestamp 1712622712
transform 1 0 1308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4867
timestamp 1712622712
transform 1 0 1348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1712622712
transform 1 0 1284 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1712622712
transform 1 0 1252 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_4870
timestamp 1712622712
transform 1 0 1540 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4871
timestamp 1712622712
transform 1 0 1532 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4872
timestamp 1712622712
transform 1 0 1460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4873
timestamp 1712622712
transform 1 0 1348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4874
timestamp 1712622712
transform 1 0 1284 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_4875
timestamp 1712622712
transform 1 0 1244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4876
timestamp 1712622712
transform 1 0 1508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4877
timestamp 1712622712
transform 1 0 1420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4878
timestamp 1712622712
transform 1 0 1476 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_4879
timestamp 1712622712
transform 1 0 1476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4880
timestamp 1712622712
transform 1 0 1388 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1712622712
transform 1 0 1356 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1712622712
transform 1 0 1388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4883
timestamp 1712622712
transform 1 0 1372 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1712622712
transform 1 0 1420 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4885
timestamp 1712622712
transform 1 0 1404 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4886
timestamp 1712622712
transform 1 0 1492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1712622712
transform 1 0 1412 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1712622712
transform 1 0 1636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4889
timestamp 1712622712
transform 1 0 1636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1712622712
transform 1 0 1572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4891
timestamp 1712622712
transform 1 0 1308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4892
timestamp 1712622712
transform 1 0 1308 0 1 755
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1712622712
transform 1 0 1780 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4894
timestamp 1712622712
transform 1 0 1700 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1712622712
transform 1 0 1756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4896
timestamp 1712622712
transform 1 0 1748 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1712622712
transform 1 0 1788 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4898
timestamp 1712622712
transform 1 0 1756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4899
timestamp 1712622712
transform 1 0 1820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4900
timestamp 1712622712
transform 1 0 1812 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1712622712
transform 1 0 1868 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_4902
timestamp 1712622712
transform 1 0 1868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4903
timestamp 1712622712
transform 1 0 1796 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4904
timestamp 1712622712
transform 1 0 1740 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1712622712
transform 1 0 1724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4906
timestamp 1712622712
transform 1 0 1708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1712622712
transform 1 0 1676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4908
timestamp 1712622712
transform 1 0 1636 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4909
timestamp 1712622712
transform 1 0 1628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4910
timestamp 1712622712
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1712622712
transform 1 0 1732 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1712622712
transform 1 0 1788 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4913
timestamp 1712622712
transform 1 0 1756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1712622712
transform 1 0 1668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4915
timestamp 1712622712
transform 1 0 1668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4916
timestamp 1712622712
transform 1 0 1676 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4917
timestamp 1712622712
transform 1 0 1668 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1712622712
transform 1 0 1724 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4919
timestamp 1712622712
transform 1 0 1684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4920
timestamp 1712622712
transform 1 0 1692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1712622712
transform 1 0 1692 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4922
timestamp 1712622712
transform 1 0 1740 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4923
timestamp 1712622712
transform 1 0 1740 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4924
timestamp 1712622712
transform 1 0 1716 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4925
timestamp 1712622712
transform 1 0 1708 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4926
timestamp 1712622712
transform 1 0 1988 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4927
timestamp 1712622712
transform 1 0 1884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4928
timestamp 1712622712
transform 1 0 1772 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4929
timestamp 1712622712
transform 1 0 1772 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4930
timestamp 1712622712
transform 1 0 1772 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1712622712
transform 1 0 1676 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1712622712
transform 1 0 1396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1712622712
transform 1 0 2124 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_4934
timestamp 1712622712
transform 1 0 2124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1712622712
transform 1 0 2108 0 1 355
box -2 -2 2 2
use M2_M1  M2_M1_4936
timestamp 1712622712
transform 1 0 1812 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1712622712
transform 1 0 1660 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4938
timestamp 1712622712
transform 1 0 1652 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4939
timestamp 1712622712
transform 1 0 1580 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4940
timestamp 1712622712
transform 1 0 1564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4941
timestamp 1712622712
transform 1 0 2164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4942
timestamp 1712622712
transform 1 0 2060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1712622712
transform 1 0 1980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4944
timestamp 1712622712
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4945
timestamp 1712622712
transform 1 0 2108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4946
timestamp 1712622712
transform 1 0 2068 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4947
timestamp 1712622712
transform 1 0 1836 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1712622712
transform 1 0 1836 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4949
timestamp 1712622712
transform 1 0 2052 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4950
timestamp 1712622712
transform 1 0 1852 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_4951
timestamp 1712622712
transform 1 0 908 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_4952
timestamp 1712622712
transform 1 0 604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4953
timestamp 1712622712
transform 1 0 1964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4954
timestamp 1712622712
transform 1 0 1948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4955
timestamp 1712622712
transform 1 0 1868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4956
timestamp 1712622712
transform 1 0 1852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1712622712
transform 1 0 2156 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1712622712
transform 1 0 2156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1712622712
transform 1 0 2300 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4960
timestamp 1712622712
transform 1 0 2220 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1712622712
transform 1 0 2020 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4962
timestamp 1712622712
transform 1 0 2012 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1712622712
transform 1 0 2004 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4964
timestamp 1712622712
transform 1 0 2004 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4965
timestamp 1712622712
transform 1 0 2108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4966
timestamp 1712622712
transform 1 0 2028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4967
timestamp 1712622712
transform 1 0 2012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4968
timestamp 1712622712
transform 1 0 1940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4969
timestamp 1712622712
transform 1 0 1900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1712622712
transform 1 0 1988 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4971
timestamp 1712622712
transform 1 0 1956 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4972
timestamp 1712622712
transform 1 0 1924 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4973
timestamp 1712622712
transform 1 0 1924 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_4974
timestamp 1712622712
transform 1 0 2148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1712622712
transform 1 0 1988 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4976
timestamp 1712622712
transform 1 0 1932 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4977
timestamp 1712622712
transform 1 0 1916 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4978
timestamp 1712622712
transform 1 0 1908 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4979
timestamp 1712622712
transform 1 0 1908 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4980
timestamp 1712622712
transform 1 0 1868 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1712622712
transform 1 0 1868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4982
timestamp 1712622712
transform 1 0 1868 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4983
timestamp 1712622712
transform 1 0 1532 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4984
timestamp 1712622712
transform 1 0 2252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4985
timestamp 1712622712
transform 1 0 1900 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4986
timestamp 1712622712
transform 1 0 2252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4987
timestamp 1712622712
transform 1 0 2228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4988
timestamp 1712622712
transform 1 0 2284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4989
timestamp 1712622712
transform 1 0 2236 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1712622712
transform 1 0 2324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4991
timestamp 1712622712
transform 1 0 2324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4992
timestamp 1712622712
transform 1 0 2396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4993
timestamp 1712622712
transform 1 0 2372 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4994
timestamp 1712622712
transform 1 0 2460 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1712622712
transform 1 0 2388 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4996
timestamp 1712622712
transform 1 0 2236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1712622712
transform 1 0 2444 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4998
timestamp 1712622712
transform 1 0 2412 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4999
timestamp 1712622712
transform 1 0 2148 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5000
timestamp 1712622712
transform 1 0 2068 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5001
timestamp 1712622712
transform 1 0 1892 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1712622712
transform 1 0 2068 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_5003
timestamp 1712622712
transform 1 0 1884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5004
timestamp 1712622712
transform 1 0 1836 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5005
timestamp 1712622712
transform 1 0 1716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5006
timestamp 1712622712
transform 1 0 2260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5007
timestamp 1712622712
transform 1 0 2212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1712622712
transform 1 0 2332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5009
timestamp 1712622712
transform 1 0 2324 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5010
timestamp 1712622712
transform 1 0 2188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5011
timestamp 1712622712
transform 1 0 2044 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5012
timestamp 1712622712
transform 1 0 2428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5013
timestamp 1712622712
transform 1 0 2308 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5014
timestamp 1712622712
transform 1 0 2060 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5015
timestamp 1712622712
transform 1 0 1964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5016
timestamp 1712622712
transform 1 0 1964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5017
timestamp 1712622712
transform 1 0 1964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5018
timestamp 1712622712
transform 1 0 1836 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5019
timestamp 1712622712
transform 1 0 1716 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5020
timestamp 1712622712
transform 1 0 1788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5021
timestamp 1712622712
transform 1 0 1700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5022
timestamp 1712622712
transform 1 0 1796 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5023
timestamp 1712622712
transform 1 0 1580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1712622712
transform 1 0 1804 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5025
timestamp 1712622712
transform 1 0 1700 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5026
timestamp 1712622712
transform 1 0 1692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5027
timestamp 1712622712
transform 1 0 1540 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5028
timestamp 1712622712
transform 1 0 1500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5029
timestamp 1712622712
transform 1 0 2300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1712622712
transform 1 0 2260 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1712622712
transform 1 0 2236 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_5032
timestamp 1712622712
transform 1 0 2084 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1712622712
transform 1 0 2076 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5034
timestamp 1712622712
transform 1 0 2068 0 1 1655
box -2 -2 2 2
use M2_M1  M2_M1_5035
timestamp 1712622712
transform 1 0 2300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5036
timestamp 1712622712
transform 1 0 2276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5037
timestamp 1712622712
transform 1 0 2500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5038
timestamp 1712622712
transform 1 0 2268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5039
timestamp 1712622712
transform 1 0 2476 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1712622712
transform 1 0 2468 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5041
timestamp 1712622712
transform 1 0 2556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1712622712
transform 1 0 2540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1712622712
transform 1 0 2460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5044
timestamp 1712622712
transform 1 0 2420 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5045
timestamp 1712622712
transform 1 0 2348 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5046
timestamp 1712622712
transform 1 0 2308 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5047
timestamp 1712622712
transform 1 0 2164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1712622712
transform 1 0 2148 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5049
timestamp 1712622712
transform 1 0 2148 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5050
timestamp 1712622712
transform 1 0 2068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5051
timestamp 1712622712
transform 1 0 2020 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5052
timestamp 1712622712
transform 1 0 2532 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1712622712
transform 1 0 2516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5054
timestamp 1712622712
transform 1 0 2492 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5055
timestamp 1712622712
transform 1 0 2420 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1712622712
transform 1 0 2388 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1712622712
transform 1 0 2164 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5058
timestamp 1712622712
transform 1 0 2124 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5059
timestamp 1712622712
transform 1 0 1620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5060
timestamp 1712622712
transform 1 0 2140 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5061
timestamp 1712622712
transform 1 0 1660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5062
timestamp 1712622712
transform 1 0 1628 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1712622712
transform 1 0 1620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1712622712
transform 1 0 2308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1712622712
transform 1 0 2212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5066
timestamp 1712622712
transform 1 0 2372 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5067
timestamp 1712622712
transform 1 0 2356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1712622712
transform 1 0 1540 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5069
timestamp 1712622712
transform 1 0 1500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1712622712
transform 1 0 1492 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5071
timestamp 1712622712
transform 1 0 1476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1712622712
transform 1 0 1676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5073
timestamp 1712622712
transform 1 0 1660 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5074
timestamp 1712622712
transform 1 0 1636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1712622712
transform 1 0 1412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5076
timestamp 1712622712
transform 1 0 3084 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1712622712
transform 1 0 2932 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5078
timestamp 1712622712
transform 1 0 2884 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5079
timestamp 1712622712
transform 1 0 2764 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5080
timestamp 1712622712
transform 1 0 2700 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5081
timestamp 1712622712
transform 1 0 2572 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1712622712
transform 1 0 1652 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5083
timestamp 1712622712
transform 1 0 1652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5084
timestamp 1712622712
transform 1 0 1612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5085
timestamp 1712622712
transform 1 0 1604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5086
timestamp 1712622712
transform 1 0 2340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5087
timestamp 1712622712
transform 1 0 2324 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1712622712
transform 1 0 2284 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1712622712
transform 1 0 2180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1712622712
transform 1 0 2492 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1712622712
transform 1 0 2316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1712622712
transform 1 0 2476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5093
timestamp 1712622712
transform 1 0 2460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5094
timestamp 1712622712
transform 1 0 2524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5095
timestamp 1712622712
transform 1 0 2516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1712622712
transform 1 0 2460 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1712622712
transform 1 0 2332 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5098
timestamp 1712622712
transform 1 0 2268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1712622712
transform 1 0 2244 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5100
timestamp 1712622712
transform 1 0 2236 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1712622712
transform 1 0 2124 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1712622712
transform 1 0 2084 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1712622712
transform 1 0 2068 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5104
timestamp 1712622712
transform 1 0 2468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1712622712
transform 1 0 2284 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5106
timestamp 1712622712
transform 1 0 2268 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5107
timestamp 1712622712
transform 1 0 2132 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1712622712
transform 1 0 2100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1712622712
transform 1 0 2108 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1712622712
transform 1 0 2052 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1712622712
transform 1 0 2020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5112
timestamp 1712622712
transform 1 0 2020 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5113
timestamp 1712622712
transform 1 0 2140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1712622712
transform 1 0 2092 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5115
timestamp 1712622712
transform 1 0 2204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5116
timestamp 1712622712
transform 1 0 2180 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5117
timestamp 1712622712
transform 1 0 2564 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5118
timestamp 1712622712
transform 1 0 2444 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5119
timestamp 1712622712
transform 1 0 2428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5120
timestamp 1712622712
transform 1 0 2372 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5121
timestamp 1712622712
transform 1 0 2260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5122
timestamp 1712622712
transform 1 0 2108 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5123
timestamp 1712622712
transform 1 0 1460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5124
timestamp 1712622712
transform 1 0 1380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5125
timestamp 1712622712
transform 1 0 2644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5126
timestamp 1712622712
transform 1 0 1756 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5127
timestamp 1712622712
transform 1 0 1420 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5128
timestamp 1712622712
transform 1 0 1492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5129
timestamp 1712622712
transform 1 0 1492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5130
timestamp 1712622712
transform 1 0 2684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5131
timestamp 1712622712
transform 1 0 2596 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5132
timestamp 1712622712
transform 1 0 2476 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5133
timestamp 1712622712
transform 1 0 2468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5134
timestamp 1712622712
transform 1 0 2460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1712622712
transform 1 0 2308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5136
timestamp 1712622712
transform 1 0 2252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5137
timestamp 1712622712
transform 1 0 1540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5138
timestamp 1712622712
transform 1 0 1396 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5139
timestamp 1712622712
transform 1 0 2340 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5140
timestamp 1712622712
transform 1 0 2268 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5141
timestamp 1712622712
transform 1 0 2260 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5142
timestamp 1712622712
transform 1 0 2220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5143
timestamp 1712622712
transform 1 0 2516 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5144
timestamp 1712622712
transform 1 0 2308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5145
timestamp 1712622712
transform 1 0 2476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5146
timestamp 1712622712
transform 1 0 2460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1712622712
transform 1 0 2580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5148
timestamp 1712622712
transform 1 0 2564 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5149
timestamp 1712622712
transform 1 0 2596 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5150
timestamp 1712622712
transform 1 0 2420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5151
timestamp 1712622712
transform 1 0 2300 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5152
timestamp 1712622712
transform 1 0 2188 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5153
timestamp 1712622712
transform 1 0 2188 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_5154
timestamp 1712622712
transform 1 0 2124 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5155
timestamp 1712622712
transform 1 0 2068 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5156
timestamp 1712622712
transform 1 0 1972 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1712622712
transform 1 0 1972 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5158
timestamp 1712622712
transform 1 0 2468 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5159
timestamp 1712622712
transform 1 0 2404 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5160
timestamp 1712622712
transform 1 0 2364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5161
timestamp 1712622712
transform 1 0 2036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5162
timestamp 1712622712
transform 1 0 1980 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1712622712
transform 1 0 2036 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5164
timestamp 1712622712
transform 1 0 2036 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1712622712
transform 1 0 2020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5166
timestamp 1712622712
transform 1 0 2020 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5167
timestamp 1712622712
transform 1 0 2132 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5168
timestamp 1712622712
transform 1 0 2116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5169
timestamp 1712622712
transform 1 0 2244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5170
timestamp 1712622712
transform 1 0 2220 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5171
timestamp 1712622712
transform 1 0 2508 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5172
timestamp 1712622712
transform 1 0 2468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1712622712
transform 1 0 2460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5174
timestamp 1712622712
transform 1 0 2388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5175
timestamp 1712622712
transform 1 0 2308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5176
timestamp 1712622712
transform 1 0 2612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5177
timestamp 1712622712
transform 1 0 1828 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5178
timestamp 1712622712
transform 1 0 1716 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5179
timestamp 1712622712
transform 1 0 1636 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5180
timestamp 1712622712
transform 1 0 1612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5181
timestamp 1712622712
transform 1 0 1940 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5182
timestamp 1712622712
transform 1 0 1908 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5183
timestamp 1712622712
transform 1 0 1860 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1712622712
transform 1 0 1844 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5185
timestamp 1712622712
transform 1 0 1820 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1712622712
transform 1 0 1820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5187
timestamp 1712622712
transform 1 0 1788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1712622712
transform 1 0 1716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5189
timestamp 1712622712
transform 1 0 1804 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5190
timestamp 1712622712
transform 1 0 1764 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5191
timestamp 1712622712
transform 1 0 1852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5192
timestamp 1712622712
transform 1 0 1804 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5193
timestamp 1712622712
transform 1 0 1788 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5194
timestamp 1712622712
transform 1 0 1844 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5195
timestamp 1712622712
transform 1 0 1836 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5196
timestamp 1712622712
transform 1 0 1836 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5197
timestamp 1712622712
transform 1 0 1820 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5198
timestamp 1712622712
transform 1 0 1820 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5199
timestamp 1712622712
transform 1 0 1932 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1712622712
transform 1 0 1716 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5201
timestamp 1712622712
transform 1 0 1932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5202
timestamp 1712622712
transform 1 0 1924 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5203
timestamp 1712622712
transform 1 0 1836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5204
timestamp 1712622712
transform 1 0 1820 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5205
timestamp 1712622712
transform 1 0 1852 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5206
timestamp 1712622712
transform 1 0 1812 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5207
timestamp 1712622712
transform 1 0 1884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5208
timestamp 1712622712
transform 1 0 1844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5209
timestamp 1712622712
transform 1 0 3004 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1712622712
transform 1 0 2868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5211
timestamp 1712622712
transform 1 0 2868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5212
timestamp 1712622712
transform 1 0 2764 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5213
timestamp 1712622712
transform 1 0 2692 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5214
timestamp 1712622712
transform 1 0 2084 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5215
timestamp 1712622712
transform 1 0 1900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1712622712
transform 1 0 1724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1712622712
transform 1 0 1756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1712622712
transform 1 0 1756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5219
timestamp 1712622712
transform 1 0 2932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5220
timestamp 1712622712
transform 1 0 2708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5221
timestamp 1712622712
transform 1 0 2708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5222
timestamp 1712622712
transform 1 0 2692 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_5223
timestamp 1712622712
transform 1 0 2676 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5224
timestamp 1712622712
transform 1 0 2676 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1712622712
transform 1 0 2524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1712622712
transform 1 0 2524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1712622712
transform 1 0 1988 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1712622712
transform 1 0 1780 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5229
timestamp 1712622712
transform 1 0 1724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5230
timestamp 1712622712
transform 1 0 1444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1712622712
transform 1 0 1356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5232
timestamp 1712622712
transform 1 0 2132 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5233
timestamp 1712622712
transform 1 0 2036 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1712622712
transform 1 0 1964 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5235
timestamp 1712622712
transform 1 0 1924 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5236
timestamp 1712622712
transform 1 0 1980 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1712622712
transform 1 0 1980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5238
timestamp 1712622712
transform 1 0 2028 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1712622712
transform 1 0 1972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1712622712
transform 1 0 1988 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5241
timestamp 1712622712
transform 1 0 1932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1712622712
transform 1 0 2364 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1712622712
transform 1 0 2188 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5244
timestamp 1712622712
transform 1 0 2292 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1712622712
transform 1 0 2188 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5246
timestamp 1712622712
transform 1 0 2036 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5247
timestamp 1712622712
transform 1 0 1988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1712622712
transform 1 0 1908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1712622712
transform 1 0 1892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5250
timestamp 1712622712
transform 1 0 1932 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1712622712
transform 1 0 1932 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1712622712
transform 1 0 2052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5253
timestamp 1712622712
transform 1 0 1972 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5254
timestamp 1712622712
transform 1 0 2172 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1712622712
transform 1 0 2068 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5256
timestamp 1712622712
transform 1 0 2220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5257
timestamp 1712622712
transform 1 0 2148 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5258
timestamp 1712622712
transform 1 0 2220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1712622712
transform 1 0 2188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5260
timestamp 1712622712
transform 1 0 2284 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_5261
timestamp 1712622712
transform 1 0 2236 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5262
timestamp 1712622712
transform 1 0 2436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5263
timestamp 1712622712
transform 1 0 2236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1712622712
transform 1 0 3044 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5265
timestamp 1712622712
transform 1 0 2988 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1712622712
transform 1 0 2764 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1712622712
transform 1 0 2484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5268
timestamp 1712622712
transform 1 0 2396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1712622712
transform 1 0 2220 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5270
timestamp 1712622712
transform 1 0 2132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5271
timestamp 1712622712
transform 1 0 2388 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1712622712
transform 1 0 2228 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5273
timestamp 1712622712
transform 1 0 2180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1712622712
transform 1 0 2172 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5275
timestamp 1712622712
transform 1 0 2276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5276
timestamp 1712622712
transform 1 0 2180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5277
timestamp 1712622712
transform 1 0 2332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5278
timestamp 1712622712
transform 1 0 2284 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1712622712
transform 1 0 2308 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1712622712
transform 1 0 2164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5281
timestamp 1712622712
transform 1 0 2476 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5282
timestamp 1712622712
transform 1 0 2276 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1712622712
transform 1 0 2340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5284
timestamp 1712622712
transform 1 0 2332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5285
timestamp 1712622712
transform 1 0 2308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1712622712
transform 1 0 2172 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5287
timestamp 1712622712
transform 1 0 2156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5288
timestamp 1712622712
transform 1 0 2196 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1712622712
transform 1 0 2188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1712622712
transform 1 0 2364 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1712622712
transform 1 0 2284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5292
timestamp 1712622712
transform 1 0 2428 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5293
timestamp 1712622712
transform 1 0 2372 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5294
timestamp 1712622712
transform 1 0 2340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1712622712
transform 1 0 2244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1712622712
transform 1 0 2460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5297
timestamp 1712622712
transform 1 0 2308 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5298
timestamp 1712622712
transform 1 0 2444 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1712622712
transform 1 0 2348 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5300
timestamp 1712622712
transform 1 0 2508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1712622712
transform 1 0 2436 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_5302
timestamp 1712622712
transform 1 0 2924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5303
timestamp 1712622712
transform 1 0 2796 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5304
timestamp 1712622712
transform 1 0 2564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1712622712
transform 1 0 2548 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1712622712
transform 1 0 2524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5307
timestamp 1712622712
transform 1 0 2524 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1712622712
transform 1 0 2460 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5309
timestamp 1712622712
transform 1 0 2412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5310
timestamp 1712622712
transform 1 0 2508 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5311
timestamp 1712622712
transform 1 0 2476 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5312
timestamp 1712622712
transform 1 0 2404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1712622712
transform 1 0 2348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5314
timestamp 1712622712
transform 1 0 2444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5315
timestamp 1712622712
transform 1 0 2436 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1712622712
transform 1 0 2468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5317
timestamp 1712622712
transform 1 0 2460 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5318
timestamp 1712622712
transform 1 0 2476 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5319
timestamp 1712622712
transform 1 0 2356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5320
timestamp 1712622712
transform 1 0 2988 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5321
timestamp 1712622712
transform 1 0 2932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5322
timestamp 1712622712
transform 1 0 2764 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5323
timestamp 1712622712
transform 1 0 2668 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5324
timestamp 1712622712
transform 1 0 2516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5325
timestamp 1712622712
transform 1 0 2468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5326
timestamp 1712622712
transform 1 0 2452 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5327
timestamp 1712622712
transform 1 0 2452 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5328
timestamp 1712622712
transform 1 0 2436 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5329
timestamp 1712622712
transform 1 0 2396 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5330
timestamp 1712622712
transform 1 0 2612 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5331
timestamp 1712622712
transform 1 0 2460 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1712622712
transform 1 0 2596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5333
timestamp 1712622712
transform 1 0 2556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5334
timestamp 1712622712
transform 1 0 2556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1712622712
transform 1 0 2316 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5336
timestamp 1712622712
transform 1 0 2292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1712622712
transform 1 0 2356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5338
timestamp 1712622712
transform 1 0 2348 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5339
timestamp 1712622712
transform 1 0 2612 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5340
timestamp 1712622712
transform 1 0 2500 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1712622712
transform 1 0 2620 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1712622712
transform 1 0 2580 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5343
timestamp 1712622712
transform 1 0 2596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5344
timestamp 1712622712
transform 1 0 2492 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1712622712
transform 1 0 2596 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1712622712
transform 1 0 2564 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5347
timestamp 1712622712
transform 1 0 2668 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5348
timestamp 1712622712
transform 1 0 2652 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5349
timestamp 1712622712
transform 1 0 2676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5350
timestamp 1712622712
transform 1 0 2660 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1712622712
transform 1 0 2764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1712622712
transform 1 0 2740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5353
timestamp 1712622712
transform 1 0 2724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5354
timestamp 1712622712
transform 1 0 2644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5355
timestamp 1712622712
transform 1 0 2596 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5356
timestamp 1712622712
transform 1 0 2548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5357
timestamp 1712622712
transform 1 0 2628 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5358
timestamp 1712622712
transform 1 0 2596 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5359
timestamp 1712622712
transform 1 0 2516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5360
timestamp 1712622712
transform 1 0 2124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5361
timestamp 1712622712
transform 1 0 2556 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5362
timestamp 1712622712
transform 1 0 2556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5363
timestamp 1712622712
transform 1 0 2572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5364
timestamp 1712622712
transform 1 0 2564 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1712622712
transform 1 0 2668 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1712622712
transform 1 0 2556 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1712622712
transform 1 0 2684 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1712622712
transform 1 0 2676 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5369
timestamp 1712622712
transform 1 0 2668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5370
timestamp 1712622712
transform 1 0 2644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1712622712
transform 1 0 2644 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5372
timestamp 1712622712
transform 1 0 2676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5373
timestamp 1712622712
transform 1 0 2660 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5374
timestamp 1712622712
transform 1 0 2620 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5375
timestamp 1712622712
transform 1 0 2572 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1712622712
transform 1 0 2724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5377
timestamp 1712622712
transform 1 0 2668 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5378
timestamp 1712622712
transform 1 0 2892 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1712622712
transform 1 0 2852 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5380
timestamp 1712622712
transform 1 0 2780 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5381
timestamp 1712622712
transform 1 0 2740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5382
timestamp 1712622712
transform 1 0 2740 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5383
timestamp 1712622712
transform 1 0 2716 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5384
timestamp 1712622712
transform 1 0 2716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5385
timestamp 1712622712
transform 1 0 2676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5386
timestamp 1712622712
transform 1 0 2652 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5387
timestamp 1712622712
transform 1 0 2100 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1712622712
transform 1 0 2100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5389
timestamp 1712622712
transform 1 0 2116 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5390
timestamp 1712622712
transform 1 0 2052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5391
timestamp 1712622712
transform 1 0 3308 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5392
timestamp 1712622712
transform 1 0 3164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5393
timestamp 1712622712
transform 1 0 3116 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5394
timestamp 1712622712
transform 1 0 2612 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1712622712
transform 1 0 2684 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5396
timestamp 1712622712
transform 1 0 2468 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5397
timestamp 1712622712
transform 1 0 2012 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5398
timestamp 1712622712
transform 1 0 1956 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5399
timestamp 1712622712
transform 1 0 1908 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5400
timestamp 1712622712
transform 1 0 1732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5401
timestamp 1712622712
transform 1 0 1716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5402
timestamp 1712622712
transform 1 0 3236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5403
timestamp 1712622712
transform 1 0 3180 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5404
timestamp 1712622712
transform 1 0 3180 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5405
timestamp 1712622712
transform 1 0 3300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5406
timestamp 1712622712
transform 1 0 3284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5407
timestamp 1712622712
transform 1 0 3212 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1712622712
transform 1 0 3180 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1712622712
transform 1 0 2692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1712622712
transform 1 0 2652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1712622712
transform 1 0 2692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5412
timestamp 1712622712
transform 1 0 2660 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5413
timestamp 1712622712
transform 1 0 2764 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_5414
timestamp 1712622712
transform 1 0 2692 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_5415
timestamp 1712622712
transform 1 0 2692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5416
timestamp 1712622712
transform 1 0 2684 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1712622712
transform 1 0 2652 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5418
timestamp 1712622712
transform 1 0 2740 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5419
timestamp 1712622712
transform 1 0 2668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5420
timestamp 1712622712
transform 1 0 2732 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1712622712
transform 1 0 2716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5422
timestamp 1712622712
transform 1 0 2884 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5423
timestamp 1712622712
transform 1 0 2876 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5424
timestamp 1712622712
transform 1 0 2860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5425
timestamp 1712622712
transform 1 0 2860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1712622712
transform 1 0 3004 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5427
timestamp 1712622712
transform 1 0 2868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1712622712
transform 1 0 3060 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5429
timestamp 1712622712
transform 1 0 3020 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5430
timestamp 1712622712
transform 1 0 3060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5431
timestamp 1712622712
transform 1 0 3020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5432
timestamp 1712622712
transform 1 0 3020 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5433
timestamp 1712622712
transform 1 0 2980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5434
timestamp 1712622712
transform 1 0 3236 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5435
timestamp 1712622712
transform 1 0 3140 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5436
timestamp 1712622712
transform 1 0 3124 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5437
timestamp 1712622712
transform 1 0 2996 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5438
timestamp 1712622712
transform 1 0 2996 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5439
timestamp 1712622712
transform 1 0 3060 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5440
timestamp 1712622712
transform 1 0 3044 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5441
timestamp 1712622712
transform 1 0 3068 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1712622712
transform 1 0 3012 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5443
timestamp 1712622712
transform 1 0 2996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5444
timestamp 1712622712
transform 1 0 2924 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5445
timestamp 1712622712
transform 1 0 2908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5446
timestamp 1712622712
transform 1 0 3116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5447
timestamp 1712622712
transform 1 0 3044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5448
timestamp 1712622712
transform 1 0 3060 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1712622712
transform 1 0 2820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1712622712
transform 1 0 2732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5451
timestamp 1712622712
transform 1 0 2724 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5452
timestamp 1712622712
transform 1 0 3116 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1712622712
transform 1 0 2972 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1712622712
transform 1 0 3060 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5455
timestamp 1712622712
transform 1 0 3020 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1712622712
transform 1 0 2996 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1712622712
transform 1 0 2972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5458
timestamp 1712622712
transform 1 0 2916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1712622712
transform 1 0 2892 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1712622712
transform 1 0 3028 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5461
timestamp 1712622712
transform 1 0 2884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5462
timestamp 1712622712
transform 1 0 2988 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5463
timestamp 1712622712
transform 1 0 2932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5464
timestamp 1712622712
transform 1 0 2876 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1712622712
transform 1 0 2876 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5466
timestamp 1712622712
transform 1 0 3060 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1712622712
transform 1 0 3012 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5468
timestamp 1712622712
transform 1 0 3268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1712622712
transform 1 0 3268 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5470
timestamp 1712622712
transform 1 0 3212 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5471
timestamp 1712622712
transform 1 0 2980 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1712622712
transform 1 0 2924 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1712622712
transform 1 0 2836 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5474
timestamp 1712622712
transform 1 0 3060 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1712622712
transform 1 0 3044 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5476
timestamp 1712622712
transform 1 0 3076 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1712622712
transform 1 0 3044 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5478
timestamp 1712622712
transform 1 0 3188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1712622712
transform 1 0 3036 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5480
timestamp 1712622712
transform 1 0 3124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1712622712
transform 1 0 3060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1712622712
transform 1 0 3204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5483
timestamp 1712622712
transform 1 0 3124 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1712622712
transform 1 0 3132 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1712622712
transform 1 0 3132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1712622712
transform 1 0 3132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1712622712
transform 1 0 3108 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1712622712
transform 1 0 2692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1712622712
transform 1 0 2692 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5490
timestamp 1712622712
transform 1 0 2660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5491
timestamp 1712622712
transform 1 0 2620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5492
timestamp 1712622712
transform 1 0 2612 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5493
timestamp 1712622712
transform 1 0 2580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1712622712
transform 1 0 2564 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5495
timestamp 1712622712
transform 1 0 2508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5496
timestamp 1712622712
transform 1 0 2500 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5497
timestamp 1712622712
transform 1 0 2500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1712622712
transform 1 0 2492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1712622712
transform 1 0 2484 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1712622712
transform 1 0 2484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5501
timestamp 1712622712
transform 1 0 2668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5502
timestamp 1712622712
transform 1 0 2660 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1712622712
transform 1 0 3116 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1712622712
transform 1 0 3116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5505
timestamp 1712622712
transform 1 0 3100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5506
timestamp 1712622712
transform 1 0 3044 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5507
timestamp 1712622712
transform 1 0 3084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5508
timestamp 1712622712
transform 1 0 3044 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1712622712
transform 1 0 2972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5510
timestamp 1712622712
transform 1 0 3044 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1712622712
transform 1 0 2748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5512
timestamp 1712622712
transform 1 0 2988 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5513
timestamp 1712622712
transform 1 0 2908 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5514
timestamp 1712622712
transform 1 0 3100 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_5515
timestamp 1712622712
transform 1 0 3076 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5516
timestamp 1712622712
transform 1 0 2924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1712622712
transform 1 0 2924 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5518
timestamp 1712622712
transform 1 0 3188 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5519
timestamp 1712622712
transform 1 0 2980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1712622712
transform 1 0 2988 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5521
timestamp 1712622712
transform 1 0 2948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1712622712
transform 1 0 2580 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5523
timestamp 1712622712
transform 1 0 2516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1712622712
transform 1 0 3092 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1712622712
transform 1 0 2964 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1712622712
transform 1 0 2972 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1712622712
transform 1 0 2924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1712622712
transform 1 0 3100 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1712622712
transform 1 0 3084 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_5530
timestamp 1712622712
transform 1 0 2932 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1712622712
transform 1 0 2924 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5532
timestamp 1712622712
transform 1 0 2892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5533
timestamp 1712622712
transform 1 0 2820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1712622712
transform 1 0 3068 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5535
timestamp 1712622712
transform 1 0 2916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5536
timestamp 1712622712
transform 1 0 3060 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5537
timestamp 1712622712
transform 1 0 3060 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1712622712
transform 1 0 3012 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5539
timestamp 1712622712
transform 1 0 3012 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5540
timestamp 1712622712
transform 1 0 3100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5541
timestamp 1712622712
transform 1 0 3044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5542
timestamp 1712622712
transform 1 0 2636 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1712622712
transform 1 0 2564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5544
timestamp 1712622712
transform 1 0 2996 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5545
timestamp 1712622712
transform 1 0 2972 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1712622712
transform 1 0 2988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5547
timestamp 1712622712
transform 1 0 2940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5548
timestamp 1712622712
transform 1 0 3108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5549
timestamp 1712622712
transform 1 0 2932 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5550
timestamp 1712622712
transform 1 0 2836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5551
timestamp 1712622712
transform 1 0 3228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5552
timestamp 1712622712
transform 1 0 3132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1712622712
transform 1 0 2892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5554
timestamp 1712622712
transform 1 0 2972 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5555
timestamp 1712622712
transform 1 0 2748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5556
timestamp 1712622712
transform 1 0 2908 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5557
timestamp 1712622712
transform 1 0 2828 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5558
timestamp 1712622712
transform 1 0 2876 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_5559
timestamp 1712622712
transform 1 0 2876 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1712622712
transform 1 0 2852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5561
timestamp 1712622712
transform 1 0 2852 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5562
timestamp 1712622712
transform 1 0 2844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5563
timestamp 1712622712
transform 1 0 2868 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5564
timestamp 1712622712
transform 1 0 2828 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5565
timestamp 1712622712
transform 1 0 2868 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5566
timestamp 1712622712
transform 1 0 2852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5567
timestamp 1712622712
transform 1 0 2740 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5568
timestamp 1712622712
transform 1 0 2660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5569
timestamp 1712622712
transform 1 0 2836 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1712622712
transform 1 0 2836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5571
timestamp 1712622712
transform 1 0 2876 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5572
timestamp 1712622712
transform 1 0 2804 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5573
timestamp 1712622712
transform 1 0 2788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5574
timestamp 1712622712
transform 1 0 2756 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5575
timestamp 1712622712
transform 1 0 2796 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5576
timestamp 1712622712
transform 1 0 2764 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1712622712
transform 1 0 2788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5578
timestamp 1712622712
transform 1 0 2772 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5579
timestamp 1712622712
transform 1 0 2908 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5580
timestamp 1712622712
transform 1 0 2788 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5581
timestamp 1712622712
transform 1 0 2916 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5582
timestamp 1712622712
transform 1 0 2884 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5583
timestamp 1712622712
transform 1 0 2980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5584
timestamp 1712622712
transform 1 0 2892 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5585
timestamp 1712622712
transform 1 0 3252 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5586
timestamp 1712622712
transform 1 0 3252 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5587
timestamp 1712622712
transform 1 0 3228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5588
timestamp 1712622712
transform 1 0 3188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1712622712
transform 1 0 2628 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5590
timestamp 1712622712
transform 1 0 2500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5591
timestamp 1712622712
transform 1 0 2916 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5592
timestamp 1712622712
transform 1 0 2796 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5593
timestamp 1712622712
transform 1 0 2796 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5594
timestamp 1712622712
transform 1 0 2780 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5595
timestamp 1712622712
transform 1 0 2812 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5596
timestamp 1712622712
transform 1 0 2700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5597
timestamp 1712622712
transform 1 0 2676 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1712622712
transform 1 0 2668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5599
timestamp 1712622712
transform 1 0 2828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5600
timestamp 1712622712
transform 1 0 2804 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5601
timestamp 1712622712
transform 1 0 2772 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5602
timestamp 1712622712
transform 1 0 2724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5603
timestamp 1712622712
transform 1 0 2868 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5604
timestamp 1712622712
transform 1 0 2836 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1712622712
transform 1 0 2836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5606
timestamp 1712622712
transform 1 0 2796 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5607
timestamp 1712622712
transform 1 0 2780 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5608
timestamp 1712622712
transform 1 0 2796 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5609
timestamp 1712622712
transform 1 0 2788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5610
timestamp 1712622712
transform 1 0 2804 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5611
timestamp 1712622712
transform 1 0 2756 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5612
timestamp 1712622712
transform 1 0 2556 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5613
timestamp 1712622712
transform 1 0 2548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1712622712
transform 1 0 2668 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1712622712
transform 1 0 2516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5616
timestamp 1712622712
transform 1 0 2604 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5617
timestamp 1712622712
transform 1 0 2564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5618
timestamp 1712622712
transform 1 0 3260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5619
timestamp 1712622712
transform 1 0 3228 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5620
timestamp 1712622712
transform 1 0 3228 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5621
timestamp 1712622712
transform 1 0 3188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5622
timestamp 1712622712
transform 1 0 3188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5623
timestamp 1712622712
transform 1 0 3380 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5624
timestamp 1712622712
transform 1 0 3332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1712622712
transform 1 0 2764 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5626
timestamp 1712622712
transform 1 0 2756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1712622712
transform 1 0 2924 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5628
timestamp 1712622712
transform 1 0 2916 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5629
timestamp 1712622712
transform 1 0 3124 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5630
timestamp 1712622712
transform 1 0 3100 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5631
timestamp 1712622712
transform 1 0 3212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1712622712
transform 1 0 3204 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1712622712
transform 1 0 3180 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5634
timestamp 1712622712
transform 1 0 3092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5635
timestamp 1712622712
transform 1 0 3332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5636
timestamp 1712622712
transform 1 0 3196 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_5637
timestamp 1712622712
transform 1 0 3436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5638
timestamp 1712622712
transform 1 0 3324 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_5639
timestamp 1712622712
transform 1 0 3340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1712622712
transform 1 0 3324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1712622712
transform 1 0 3068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5642
timestamp 1712622712
transform 1 0 2892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5643
timestamp 1712622712
transform 1 0 3364 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1712622712
transform 1 0 3364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5645
timestamp 1712622712
transform 1 0 3308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1712622712
transform 1 0 3292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1712622712
transform 1 0 3244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1712622712
transform 1 0 3244 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5649
timestamp 1712622712
transform 1 0 3348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5650
timestamp 1712622712
transform 1 0 3300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1712622712
transform 1 0 3196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1712622712
transform 1 0 3188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5653
timestamp 1712622712
transform 1 0 3396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5654
timestamp 1712622712
transform 1 0 3388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5655
timestamp 1712622712
transform 1 0 3372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5656
timestamp 1712622712
transform 1 0 3340 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1712622712
transform 1 0 3324 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1712622712
transform 1 0 3284 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1712622712
transform 1 0 3404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1712622712
transform 1 0 3372 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5661
timestamp 1712622712
transform 1 0 3420 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1712622712
transform 1 0 3388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5663
timestamp 1712622712
transform 1 0 3364 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5664
timestamp 1712622712
transform 1 0 2932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5665
timestamp 1712622712
transform 1 0 2900 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1712622712
transform 1 0 3348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1712622712
transform 1 0 3308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5668
timestamp 1712622712
transform 1 0 3284 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5669
timestamp 1712622712
transform 1 0 3052 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5670
timestamp 1712622712
transform 1 0 2964 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5671
timestamp 1712622712
transform 1 0 2924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1712622712
transform 1 0 3404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5673
timestamp 1712622712
transform 1 0 3404 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1712622712
transform 1 0 3268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5675
timestamp 1712622712
transform 1 0 3100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1712622712
transform 1 0 2996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5677
timestamp 1712622712
transform 1 0 2940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5678
timestamp 1712622712
transform 1 0 2988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5679
timestamp 1712622712
transform 1 0 2988 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5680
timestamp 1712622712
transform 1 0 3100 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1712622712
transform 1 0 3092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1712622712
transform 1 0 3324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5683
timestamp 1712622712
transform 1 0 3316 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5684
timestamp 1712622712
transform 1 0 3420 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5685
timestamp 1712622712
transform 1 0 3396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5686
timestamp 1712622712
transform 1 0 3316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5687
timestamp 1712622712
transform 1 0 3244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5688
timestamp 1712622712
transform 1 0 3156 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5689
timestamp 1712622712
transform 1 0 3364 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1712622712
transform 1 0 3300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5691
timestamp 1712622712
transform 1 0 3276 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1712622712
transform 1 0 3380 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1712622712
transform 1 0 3308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1712622712
transform 1 0 3292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1712622712
transform 1 0 3356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1712622712
transform 1 0 3260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5697
timestamp 1712622712
transform 1 0 3324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5698
timestamp 1712622712
transform 1 0 3292 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5699
timestamp 1712622712
transform 1 0 3404 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1712622712
transform 1 0 3356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5701
timestamp 1712622712
transform 1 0 3396 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5702
timestamp 1712622712
transform 1 0 3380 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5703
timestamp 1712622712
transform 1 0 3380 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5704
timestamp 1712622712
transform 1 0 3348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5705
timestamp 1712622712
transform 1 0 3292 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5706
timestamp 1712622712
transform 1 0 3228 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1712622712
transform 1 0 3252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5708
timestamp 1712622712
transform 1 0 3252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5709
timestamp 1712622712
transform 1 0 3252 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_5710
timestamp 1712622712
transform 1 0 3188 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5711
timestamp 1712622712
transform 1 0 3132 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1712622712
transform 1 0 3188 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5713
timestamp 1712622712
transform 1 0 3124 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5714
timestamp 1712622712
transform 1 0 3268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5715
timestamp 1712622712
transform 1 0 3164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5716
timestamp 1712622712
transform 1 0 3196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5717
timestamp 1712622712
transform 1 0 3060 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5718
timestamp 1712622712
transform 1 0 3036 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5719
timestamp 1712622712
transform 1 0 2924 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5720
timestamp 1712622712
transform 1 0 2924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1712622712
transform 1 0 2716 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5722
timestamp 1712622712
transform 1 0 2700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5723
timestamp 1712622712
transform 1 0 2940 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5724
timestamp 1712622712
transform 1 0 2932 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5725
timestamp 1712622712
transform 1 0 3076 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5726
timestamp 1712622712
transform 1 0 2988 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5727
timestamp 1712622712
transform 1 0 2804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5728
timestamp 1712622712
transform 1 0 2804 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5729
timestamp 1712622712
transform 1 0 2604 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5730
timestamp 1712622712
transform 1 0 2588 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5731
timestamp 1712622712
transform 1 0 2732 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5732
timestamp 1712622712
transform 1 0 2580 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5733
timestamp 1712622712
transform 1 0 2516 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5734
timestamp 1712622712
transform 1 0 2516 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5735
timestamp 1712622712
transform 1 0 2388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5736
timestamp 1712622712
transform 1 0 2388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5737
timestamp 1712622712
transform 1 0 1996 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5738
timestamp 1712622712
transform 1 0 1956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5739
timestamp 1712622712
transform 1 0 2308 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5740
timestamp 1712622712
transform 1 0 2268 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5741
timestamp 1712622712
transform 1 0 2188 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5742
timestamp 1712622712
transform 1 0 2188 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5743
timestamp 1712622712
transform 1 0 2068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5744
timestamp 1712622712
transform 1 0 2068 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5745
timestamp 1712622712
transform 1 0 1836 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5746
timestamp 1712622712
transform 1 0 1804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5747
timestamp 1712622712
transform 1 0 1940 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5748
timestamp 1712622712
transform 1 0 1836 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5749
timestamp 1712622712
transform 1 0 1716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5750
timestamp 1712622712
transform 1 0 1668 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5751
timestamp 1712622712
transform 1 0 1604 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5752
timestamp 1712622712
transform 1 0 1604 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5753
timestamp 1712622712
transform 1 0 1452 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5754
timestamp 1712622712
transform 1 0 1412 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5755
timestamp 1712622712
transform 1 0 1356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5756
timestamp 1712622712
transform 1 0 1348 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1712622712
transform 1 0 1252 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5758
timestamp 1712622712
transform 1 0 1252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5759
timestamp 1712622712
transform 1 0 1148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5760
timestamp 1712622712
transform 1 0 1052 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5761
timestamp 1712622712
transform 1 0 924 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5762
timestamp 1712622712
transform 1 0 924 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5763
timestamp 1712622712
transform 1 0 156 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5764
timestamp 1712622712
transform 1 0 148 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5765
timestamp 1712622712
transform 1 0 116 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5766
timestamp 1712622712
transform 1 0 116 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5767
timestamp 1712622712
transform 1 0 228 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5768
timestamp 1712622712
transform 1 0 196 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5769
timestamp 1712622712
transform 1 0 356 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5770
timestamp 1712622712
transform 1 0 292 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5771
timestamp 1712622712
transform 1 0 452 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5772
timestamp 1712622712
transform 1 0 364 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5773
timestamp 1712622712
transform 1 0 412 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5774
timestamp 1712622712
transform 1 0 412 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5775
timestamp 1712622712
transform 1 0 468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5776
timestamp 1712622712
transform 1 0 428 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5777
timestamp 1712622712
transform 1 0 612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5778
timestamp 1712622712
transform 1 0 612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5779
timestamp 1712622712
transform 1 0 708 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5780
timestamp 1712622712
transform 1 0 676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5781
timestamp 1712622712
transform 1 0 908 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5782
timestamp 1712622712
transform 1 0 844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5783
timestamp 1712622712
transform 1 0 1140 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1712622712
transform 1 0 1140 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5785
timestamp 1712622712
transform 1 0 3060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5786
timestamp 1712622712
transform 1 0 3052 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5787
timestamp 1712622712
transform 1 0 3036 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5788
timestamp 1712622712
transform 1 0 2948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5789
timestamp 1712622712
transform 1 0 3076 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1712622712
transform 1 0 3052 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5791
timestamp 1712622712
transform 1 0 3068 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5792
timestamp 1712622712
transform 1 0 3044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5793
timestamp 1712622712
transform 1 0 3164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5794
timestamp 1712622712
transform 1 0 2972 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5795
timestamp 1712622712
transform 1 0 2956 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5796
timestamp 1712622712
transform 1 0 3036 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5797
timestamp 1712622712
transform 1 0 2956 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1712622712
transform 1 0 2908 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5799
timestamp 1712622712
transform 1 0 2828 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5800
timestamp 1712622712
transform 1 0 2948 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5801
timestamp 1712622712
transform 1 0 2916 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1712622712
transform 1 0 2988 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1712622712
transform 1 0 2876 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5804
timestamp 1712622712
transform 1 0 2820 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5805
timestamp 1712622712
transform 1 0 2796 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5806
timestamp 1712622712
transform 1 0 2820 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_5807
timestamp 1712622712
transform 1 0 2676 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5808
timestamp 1712622712
transform 1 0 2660 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5809
timestamp 1712622712
transform 1 0 2612 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5810
timestamp 1712622712
transform 1 0 2276 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5811
timestamp 1712622712
transform 1 0 2172 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1712622712
transform 1 0 2124 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5813
timestamp 1712622712
transform 1 0 1124 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5814
timestamp 1712622712
transform 1 0 2452 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5815
timestamp 1712622712
transform 1 0 2388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1712622712
transform 1 0 2172 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5817
timestamp 1712622712
transform 1 0 1772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5818
timestamp 1712622712
transform 1 0 1652 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5819
timestamp 1712622712
transform 1 0 1332 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5820
timestamp 1712622712
transform 1 0 1228 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5821
timestamp 1712622712
transform 1 0 1076 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5822
timestamp 1712622712
transform 1 0 996 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5823
timestamp 1712622712
transform 1 0 1076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5824
timestamp 1712622712
transform 1 0 932 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5825
timestamp 1712622712
transform 1 0 868 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5826
timestamp 1712622712
transform 1 0 868 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5827
timestamp 1712622712
transform 1 0 860 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5828
timestamp 1712622712
transform 1 0 1148 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5829
timestamp 1712622712
transform 1 0 956 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5830
timestamp 1712622712
transform 1 0 1164 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5831
timestamp 1712622712
transform 1 0 1132 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5832
timestamp 1712622712
transform 1 0 908 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5833
timestamp 1712622712
transform 1 0 788 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5834
timestamp 1712622712
transform 1 0 564 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5835
timestamp 1712622712
transform 1 0 2092 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5836
timestamp 1712622712
transform 1 0 1980 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5837
timestamp 1712622712
transform 1 0 1860 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5838
timestamp 1712622712
transform 1 0 1756 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5839
timestamp 1712622712
transform 1 0 2100 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5840
timestamp 1712622712
transform 1 0 1988 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5841
timestamp 1712622712
transform 1 0 1940 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5842
timestamp 1712622712
transform 1 0 1756 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1712622712
transform 1 0 1564 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5844
timestamp 1712622712
transform 1 0 1484 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5845
timestamp 1712622712
transform 1 0 2116 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5846
timestamp 1712622712
transform 1 0 2092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5847
timestamp 1712622712
transform 1 0 2436 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1712622712
transform 1 0 2412 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5849
timestamp 1712622712
transform 1 0 2084 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5850
timestamp 1712622712
transform 1 0 2068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5851
timestamp 1712622712
transform 1 0 1956 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5852
timestamp 1712622712
transform 1 0 3148 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5853
timestamp 1712622712
transform 1 0 3084 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5854
timestamp 1712622712
transform 1 0 2836 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_5855
timestamp 1712622712
transform 1 0 2660 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1712622712
transform 1 0 2652 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5857
timestamp 1712622712
transform 1 0 2436 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5858
timestamp 1712622712
transform 1 0 2372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5859
timestamp 1712622712
transform 1 0 2868 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5860
timestamp 1712622712
transform 1 0 2828 0 1 2985
box -2 -2 2 2
use M2_M1  M2_M1_5861
timestamp 1712622712
transform 1 0 956 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5862
timestamp 1712622712
transform 1 0 860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5863
timestamp 1712622712
transform 1 0 564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1712622712
transform 1 0 524 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5865
timestamp 1712622712
transform 1 0 436 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5866
timestamp 1712622712
transform 1 0 404 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5867
timestamp 1712622712
transform 1 0 388 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5868
timestamp 1712622712
transform 1 0 372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5869
timestamp 1712622712
transform 1 0 244 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5870
timestamp 1712622712
transform 1 0 220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5871
timestamp 1712622712
transform 1 0 212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5872
timestamp 1712622712
transform 1 0 2940 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5873
timestamp 1712622712
transform 1 0 2852 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5874
timestamp 1712622712
transform 1 0 2780 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5875
timestamp 1712622712
transform 1 0 2740 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5876
timestamp 1712622712
transform 1 0 2556 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5877
timestamp 1712622712
transform 1 0 3092 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1712622712
transform 1 0 3092 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5879
timestamp 1712622712
transform 1 0 3068 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5880
timestamp 1712622712
transform 1 0 3052 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1712622712
transform 1 0 3124 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5882
timestamp 1712622712
transform 1 0 3100 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1712622712
transform 1 0 3036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1712622712
transform 1 0 2972 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1712622712
transform 1 0 3020 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5886
timestamp 1712622712
transform 1 0 2996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1712622712
transform 1 0 2556 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5888
timestamp 1712622712
transform 1 0 2540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5889
timestamp 1712622712
transform 1 0 2556 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5890
timestamp 1712622712
transform 1 0 2524 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5891
timestamp 1712622712
transform 1 0 2596 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5892
timestamp 1712622712
transform 1 0 2580 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5893
timestamp 1712622712
transform 1 0 2548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5894
timestamp 1712622712
transform 1 0 2508 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5895
timestamp 1712622712
transform 1 0 2460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5896
timestamp 1712622712
transform 1 0 2892 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5897
timestamp 1712622712
transform 1 0 2788 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5898
timestamp 1712622712
transform 1 0 2740 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5899
timestamp 1712622712
transform 1 0 2716 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5900
timestamp 1712622712
transform 1 0 2764 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1712622712
transform 1 0 2644 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5902
timestamp 1712622712
transform 1 0 2676 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5903
timestamp 1712622712
transform 1 0 2644 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_5904
timestamp 1712622712
transform 1 0 2652 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5905
timestamp 1712622712
transform 1 0 2612 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5906
timestamp 1712622712
transform 1 0 2628 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5907
timestamp 1712622712
transform 1 0 2580 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5908
timestamp 1712622712
transform 1 0 2468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5909
timestamp 1712622712
transform 1 0 2204 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5910
timestamp 1712622712
transform 1 0 2772 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5911
timestamp 1712622712
transform 1 0 2668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5912
timestamp 1712622712
transform 1 0 2692 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1712622712
transform 1 0 2660 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_5914
timestamp 1712622712
transform 1 0 2676 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5915
timestamp 1712622712
transform 1 0 2620 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1712622712
transform 1 0 2452 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5917
timestamp 1712622712
transform 1 0 2428 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5918
timestamp 1712622712
transform 1 0 2460 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5919
timestamp 1712622712
transform 1 0 2436 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5920
timestamp 1712622712
transform 1 0 2188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5921
timestamp 1712622712
transform 1 0 2116 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5922
timestamp 1712622712
transform 1 0 2012 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5923
timestamp 1712622712
transform 1 0 2372 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5924
timestamp 1712622712
transform 1 0 2332 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1712622712
transform 1 0 2324 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5926
timestamp 1712622712
transform 1 0 2228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1712622712
transform 1 0 2212 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5928
timestamp 1712622712
transform 1 0 2020 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5929
timestamp 1712622712
transform 1 0 2412 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1712622712
transform 1 0 2380 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5931
timestamp 1712622712
transform 1 0 2260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5932
timestamp 1712622712
transform 1 0 2012 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5933
timestamp 1712622712
transform 1 0 2012 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5934
timestamp 1712622712
transform 1 0 2068 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5935
timestamp 1712622712
transform 1 0 2004 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5936
timestamp 1712622712
transform 1 0 2332 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1712622712
transform 1 0 2300 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5938
timestamp 1712622712
transform 1 0 2132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5939
timestamp 1712622712
transform 1 0 2036 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5940
timestamp 1712622712
transform 1 0 1900 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5941
timestamp 1712622712
transform 1 0 2316 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5942
timestamp 1712622712
transform 1 0 2076 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5943
timestamp 1712622712
transform 1 0 2356 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5944
timestamp 1712622712
transform 1 0 2308 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1712622712
transform 1 0 2308 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5946
timestamp 1712622712
transform 1 0 2276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5947
timestamp 1712622712
transform 1 0 2172 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1712622712
transform 1 0 1980 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5949
timestamp 1712622712
transform 1 0 2340 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5950
timestamp 1712622712
transform 1 0 2292 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5951
timestamp 1712622712
transform 1 0 2356 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5952
timestamp 1712622712
transform 1 0 2284 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5953
timestamp 1712622712
transform 1 0 2364 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5954
timestamp 1712622712
transform 1 0 2356 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1712622712
transform 1 0 2212 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5956
timestamp 1712622712
transform 1 0 2204 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5957
timestamp 1712622712
transform 1 0 2324 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5958
timestamp 1712622712
transform 1 0 2196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5959
timestamp 1712622712
transform 1 0 2324 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5960
timestamp 1712622712
transform 1 0 2324 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5961
timestamp 1712622712
transform 1 0 2132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5962
timestamp 1712622712
transform 1 0 2124 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_5963
timestamp 1712622712
transform 1 0 2164 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5964
timestamp 1712622712
transform 1 0 2124 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5965
timestamp 1712622712
transform 1 0 2220 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1712622712
transform 1 0 2196 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5967
timestamp 1712622712
transform 1 0 1972 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5968
timestamp 1712622712
transform 1 0 1956 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5969
timestamp 1712622712
transform 1 0 1916 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5970
timestamp 1712622712
transform 1 0 1788 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5971
timestamp 1712622712
transform 1 0 2028 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5972
timestamp 1712622712
transform 1 0 1836 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5973
timestamp 1712622712
transform 1 0 2268 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5974
timestamp 1712622712
transform 1 0 2036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5975
timestamp 1712622712
transform 1 0 1940 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5976
timestamp 1712622712
transform 1 0 1932 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5977
timestamp 1712622712
transform 1 0 1924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5978
timestamp 1712622712
transform 1 0 1980 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5979
timestamp 1712622712
transform 1 0 1900 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5980
timestamp 1712622712
transform 1 0 1860 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5981
timestamp 1712622712
transform 1 0 1756 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5982
timestamp 1712622712
transform 1 0 1724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5983
timestamp 1712622712
transform 1 0 1692 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5984
timestamp 1712622712
transform 1 0 1812 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1712622712
transform 1 0 1812 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_5986
timestamp 1712622712
transform 1 0 1908 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5987
timestamp 1712622712
transform 1 0 1804 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5988
timestamp 1712622712
transform 1 0 1916 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5989
timestamp 1712622712
transform 1 0 1828 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5990
timestamp 1712622712
transform 1 0 1908 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1712622712
transform 1 0 1852 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5992
timestamp 1712622712
transform 1 0 1788 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5993
timestamp 1712622712
transform 1 0 1732 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5994
timestamp 1712622712
transform 1 0 1668 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5995
timestamp 1712622712
transform 1 0 1652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5996
timestamp 1712622712
transform 1 0 1956 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_5997
timestamp 1712622712
transform 1 0 1940 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1712622712
transform 1 0 1948 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5999
timestamp 1712622712
transform 1 0 1932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6000
timestamp 1712622712
transform 1 0 1948 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6001
timestamp 1712622712
transform 1 0 1884 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6002
timestamp 1712622712
transform 1 0 1708 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6003
timestamp 1712622712
transform 1 0 1676 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6004
timestamp 1712622712
transform 1 0 1772 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6005
timestamp 1712622712
transform 1 0 1700 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6006
timestamp 1712622712
transform 1 0 1772 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6007
timestamp 1712622712
transform 1 0 1764 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6008
timestamp 1712622712
transform 1 0 1636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6009
timestamp 1712622712
transform 1 0 1612 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6010
timestamp 1712622712
transform 1 0 1716 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6011
timestamp 1712622712
transform 1 0 1628 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6012
timestamp 1712622712
transform 1 0 1716 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6013
timestamp 1712622712
transform 1 0 1660 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6014
timestamp 1712622712
transform 1 0 1892 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6015
timestamp 1712622712
transform 1 0 1820 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6016
timestamp 1712622712
transform 1 0 1772 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6017
timestamp 1712622712
transform 1 0 1812 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6018
timestamp 1712622712
transform 1 0 1660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6019
timestamp 1712622712
transform 1 0 1596 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6020
timestamp 1712622712
transform 1 0 1580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6021
timestamp 1712622712
transform 1 0 1556 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6022
timestamp 1712622712
transform 1 0 1540 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6023
timestamp 1712622712
transform 1 0 1756 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6024
timestamp 1712622712
transform 1 0 1644 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6025
timestamp 1712622712
transform 1 0 1588 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6026
timestamp 1712622712
transform 1 0 1564 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6027
timestamp 1712622712
transform 1 0 1548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6028
timestamp 1712622712
transform 1 0 1508 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6029
timestamp 1712622712
transform 1 0 1508 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6030
timestamp 1712622712
transform 1 0 1468 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6031
timestamp 1712622712
transform 1 0 1444 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6032
timestamp 1712622712
transform 1 0 1540 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1712622712
transform 1 0 1436 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6034
timestamp 1712622712
transform 1 0 1684 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6035
timestamp 1712622712
transform 1 0 1468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6036
timestamp 1712622712
transform 1 0 1452 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6037
timestamp 1712622712
transform 1 0 1420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1712622712
transform 1 0 1276 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6039
timestamp 1712622712
transform 1 0 1236 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6040
timestamp 1712622712
transform 1 0 1652 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1712622712
transform 1 0 1548 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1712622712
transform 1 0 1356 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6043
timestamp 1712622712
transform 1 0 1340 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6044
timestamp 1712622712
transform 1 0 1444 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6045
timestamp 1712622712
transform 1 0 1348 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6046
timestamp 1712622712
transform 1 0 1572 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6047
timestamp 1712622712
transform 1 0 1452 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6048
timestamp 1712622712
transform 1 0 1260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6049
timestamp 1712622712
transform 1 0 1236 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6050
timestamp 1712622712
transform 1 0 1308 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6051
timestamp 1712622712
transform 1 0 1252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6052
timestamp 1712622712
transform 1 0 1588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6053
timestamp 1712622712
transform 1 0 1332 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6054
timestamp 1712622712
transform 1 0 1196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6055
timestamp 1712622712
transform 1 0 1188 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6056
timestamp 1712622712
transform 1 0 1268 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6057
timestamp 1712622712
transform 1 0 1188 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6058
timestamp 1712622712
transform 1 0 1532 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6059
timestamp 1712622712
transform 1 0 1276 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6060
timestamp 1712622712
transform 1 0 1596 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1712622712
transform 1 0 1508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6062
timestamp 1712622712
transform 1 0 1476 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6063
timestamp 1712622712
transform 1 0 1476 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6064
timestamp 1712622712
transform 1 0 1364 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6065
timestamp 1712622712
transform 1 0 1356 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6066
timestamp 1712622712
transform 1 0 1252 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6067
timestamp 1712622712
transform 1 0 1148 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6068
timestamp 1712622712
transform 1 0 1036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6069
timestamp 1712622712
transform 1 0 1020 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1712622712
transform 1 0 1180 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6071
timestamp 1712622712
transform 1 0 1140 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6072
timestamp 1712622712
transform 1 0 1332 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6073
timestamp 1712622712
transform 1 0 1132 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6074
timestamp 1712622712
transform 1 0 1356 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6075
timestamp 1712622712
transform 1 0 1332 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6076
timestamp 1712622712
transform 1 0 1460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6077
timestamp 1712622712
transform 1 0 1340 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6078
timestamp 1712622712
transform 1 0 1228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6079
timestamp 1712622712
transform 1 0 1124 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1712622712
transform 1 0 1012 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1712622712
transform 1 0 996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6082
timestamp 1712622712
transform 1 0 964 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6083
timestamp 1712622712
transform 1 0 260 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6084
timestamp 1712622712
transform 1 0 1220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6085
timestamp 1712622712
transform 1 0 932 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6086
timestamp 1712622712
transform 1 0 1244 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6087
timestamp 1712622712
transform 1 0 1220 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6088
timestamp 1712622712
transform 1 0 556 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6089
timestamp 1712622712
transform 1 0 244 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6090
timestamp 1712622712
transform 1 0 1116 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1712622712
transform 1 0 548 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6092
timestamp 1712622712
transform 1 0 1140 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6093
timestamp 1712622712
transform 1 0 1116 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6094
timestamp 1712622712
transform 1 0 660 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6095
timestamp 1712622712
transform 1 0 292 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6096
timestamp 1712622712
transform 1 0 1036 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6097
timestamp 1712622712
transform 1 0 628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6098
timestamp 1712622712
transform 1 0 1036 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6099
timestamp 1712622712
transform 1 0 1028 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6100
timestamp 1712622712
transform 1 0 1020 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6101
timestamp 1712622712
transform 1 0 988 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1712622712
transform 1 0 988 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6103
timestamp 1712622712
transform 1 0 964 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1712622712
transform 1 0 932 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6105
timestamp 1712622712
transform 1 0 1020 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6106
timestamp 1712622712
transform 1 0 852 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6107
timestamp 1712622712
transform 1 0 756 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6108
timestamp 1712622712
transform 1 0 1060 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6109
timestamp 1712622712
transform 1 0 892 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1712622712
transform 1 0 612 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6111
timestamp 1712622712
transform 1 0 580 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6112
timestamp 1712622712
transform 1 0 572 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6113
timestamp 1712622712
transform 1 0 572 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6114
timestamp 1712622712
transform 1 0 532 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6115
timestamp 1712622712
transform 1 0 420 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6116
timestamp 1712622712
transform 1 0 660 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6117
timestamp 1712622712
transform 1 0 524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6118
timestamp 1712622712
transform 1 0 756 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6119
timestamp 1712622712
transform 1 0 660 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6120
timestamp 1712622712
transform 1 0 956 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1712622712
transform 1 0 900 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6122
timestamp 1712622712
transform 1 0 716 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6123
timestamp 1712622712
transform 1 0 692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6124
timestamp 1712622712
transform 1 0 692 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6125
timestamp 1712622712
transform 1 0 644 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6126
timestamp 1712622712
transform 1 0 468 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6127
timestamp 1712622712
transform 1 0 444 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6128
timestamp 1712622712
transform 1 0 604 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6129
timestamp 1712622712
transform 1 0 452 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6130
timestamp 1712622712
transform 1 0 700 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6131
timestamp 1712622712
transform 1 0 628 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1712622712
transform 1 0 460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6133
timestamp 1712622712
transform 1 0 436 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6134
timestamp 1712622712
transform 1 0 596 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6135
timestamp 1712622712
transform 1 0 452 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6136
timestamp 1712622712
transform 1 0 660 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6137
timestamp 1712622712
transform 1 0 636 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6138
timestamp 1712622712
transform 1 0 500 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6139
timestamp 1712622712
transform 1 0 484 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6140
timestamp 1712622712
transform 1 0 604 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1712622712
transform 1 0 492 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6142
timestamp 1712622712
transform 1 0 700 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6143
timestamp 1712622712
transform 1 0 636 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6144
timestamp 1712622712
transform 1 0 916 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6145
timestamp 1712622712
transform 1 0 844 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6146
timestamp 1712622712
transform 1 0 836 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6147
timestamp 1712622712
transform 1 0 852 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6148
timestamp 1712622712
transform 1 0 788 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6149
timestamp 1712622712
transform 1 0 772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6150
timestamp 1712622712
transform 1 0 740 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6151
timestamp 1712622712
transform 1 0 708 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6152
timestamp 1712622712
transform 1 0 676 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1712622712
transform 1 0 892 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6154
timestamp 1712622712
transform 1 0 796 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6155
timestamp 1712622712
transform 1 0 716 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6156
timestamp 1712622712
transform 1 0 700 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6157
timestamp 1712622712
transform 1 0 668 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6158
timestamp 1712622712
transform 1 0 620 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6159
timestamp 1712622712
transform 1 0 604 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6160
timestamp 1712622712
transform 1 0 580 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6161
timestamp 1712622712
transform 1 0 788 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6162
timestamp 1712622712
transform 1 0 596 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6163
timestamp 1712622712
transform 1 0 908 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6164
timestamp 1712622712
transform 1 0 892 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6165
timestamp 1712622712
transform 1 0 780 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6166
timestamp 1712622712
transform 1 0 748 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6167
timestamp 1712622712
transform 1 0 716 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6168
timestamp 1712622712
transform 1 0 788 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6169
timestamp 1712622712
transform 1 0 756 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6170
timestamp 1712622712
transform 1 0 668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1712622712
transform 1 0 620 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6172
timestamp 1712622712
transform 1 0 740 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6173
timestamp 1712622712
transform 1 0 660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6174
timestamp 1712622712
transform 1 0 740 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1712622712
transform 1 0 692 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6176
timestamp 1712622712
transform 1 0 884 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6177
timestamp 1712622712
transform 1 0 852 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6178
timestamp 1712622712
transform 1 0 804 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6179
timestamp 1712622712
transform 1 0 644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6180
timestamp 1712622712
transform 1 0 980 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6181
timestamp 1712622712
transform 1 0 972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6182
timestamp 1712622712
transform 1 0 924 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6183
timestamp 1712622712
transform 1 0 724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6184
timestamp 1712622712
transform 1 0 940 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6185
timestamp 1712622712
transform 1 0 940 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6186
timestamp 1712622712
transform 1 0 900 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6187
timestamp 1712622712
transform 1 0 828 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6188
timestamp 1712622712
transform 1 0 780 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6189
timestamp 1712622712
transform 1 0 772 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6190
timestamp 1712622712
transform 1 0 1676 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6191
timestamp 1712622712
transform 1 0 1668 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6192
timestamp 1712622712
transform 1 0 1796 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6193
timestamp 1712622712
transform 1 0 1780 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6194
timestamp 1712622712
transform 1 0 1892 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6195
timestamp 1712622712
transform 1 0 1796 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6196
timestamp 1712622712
transform 1 0 1692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6197
timestamp 1712622712
transform 1 0 1196 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6198
timestamp 1712622712
transform 1 0 1964 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6199
timestamp 1712622712
transform 1 0 1924 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6200
timestamp 1712622712
transform 1 0 3148 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6201
timestamp 1712622712
transform 1 0 2948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6202
timestamp 1712622712
transform 1 0 2820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6203
timestamp 1712622712
transform 1 0 2796 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6204
timestamp 1712622712
transform 1 0 2772 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6205
timestamp 1712622712
transform 1 0 2396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6206
timestamp 1712622712
transform 1 0 2332 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6207
timestamp 1712622712
transform 1 0 2180 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6208
timestamp 1712622712
transform 1 0 2084 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6209
timestamp 1712622712
transform 1 0 1820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6210
timestamp 1712622712
transform 1 0 1132 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6211
timestamp 1712622712
transform 1 0 916 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6212
timestamp 1712622712
transform 1 0 708 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6213
timestamp 1712622712
transform 1 0 620 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6214
timestamp 1712622712
transform 1 0 492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6215
timestamp 1712622712
transform 1 0 468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6216
timestamp 1712622712
transform 1 0 444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6217
timestamp 1712622712
transform 1 0 3148 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6218
timestamp 1712622712
transform 1 0 3132 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6219
timestamp 1712622712
transform 1 0 3244 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6220
timestamp 1712622712
transform 1 0 3156 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6221
timestamp 1712622712
transform 1 0 3124 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6222
timestamp 1712622712
transform 1 0 3156 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6223
timestamp 1712622712
transform 1 0 3092 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6224
timestamp 1712622712
transform 1 0 3028 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6225
timestamp 1712622712
transform 1 0 2908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6226
timestamp 1712622712
transform 1 0 2620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6227
timestamp 1712622712
transform 1 0 2412 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6228
timestamp 1712622712
transform 1 0 2340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6229
timestamp 1712622712
transform 1 0 1988 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6230
timestamp 1712622712
transform 1 0 1860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6231
timestamp 1712622712
transform 1 0 1684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6232
timestamp 1712622712
transform 1 0 1524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6233
timestamp 1712622712
transform 1 0 1252 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6234
timestamp 1712622712
transform 1 0 2508 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6235
timestamp 1712622712
transform 1 0 2372 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6236
timestamp 1712622712
transform 1 0 1932 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6237
timestamp 1712622712
transform 1 0 1908 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1712622712
transform 1 0 908 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6239
timestamp 1712622712
transform 1 0 852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6240
timestamp 1712622712
transform 1 0 2052 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6241
timestamp 1712622712
transform 1 0 1884 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6242
timestamp 1712622712
transform 1 0 1260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6243
timestamp 1712622712
transform 1 0 1220 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6244
timestamp 1712622712
transform 1 0 1420 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6245
timestamp 1712622712
transform 1 0 1412 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6246
timestamp 1712622712
transform 1 0 2260 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6247
timestamp 1712622712
transform 1 0 2260 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6248
timestamp 1712622712
transform 1 0 3140 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6249
timestamp 1712622712
transform 1 0 3100 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6250
timestamp 1712622712
transform 1 0 2724 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6251
timestamp 1712622712
transform 1 0 2652 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6252
timestamp 1712622712
transform 1 0 3132 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6253
timestamp 1712622712
transform 1 0 3132 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6254
timestamp 1712622712
transform 1 0 2844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6255
timestamp 1712622712
transform 1 0 2764 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6256
timestamp 1712622712
transform 1 0 2636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6257
timestamp 1712622712
transform 1 0 2556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6258
timestamp 1712622712
transform 1 0 2756 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6259
timestamp 1712622712
transform 1 0 2740 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6260
timestamp 1712622712
transform 1 0 2764 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6261
timestamp 1712622712
transform 1 0 2764 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6262
timestamp 1712622712
transform 1 0 2452 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6263
timestamp 1712622712
transform 1 0 2428 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6264
timestamp 1712622712
transform 1 0 2092 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6265
timestamp 1712622712
transform 1 0 2020 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6266
timestamp 1712622712
transform 1 0 2348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1712622712
transform 1 0 2300 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6268
timestamp 1712622712
transform 1 0 2212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6269
timestamp 1712622712
transform 1 0 2204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6270
timestamp 1712622712
transform 1 0 2116 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6271
timestamp 1712622712
transform 1 0 2036 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6272
timestamp 1712622712
transform 1 0 1812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6273
timestamp 1712622712
transform 1 0 1740 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6274
timestamp 1712622712
transform 1 0 1956 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6275
timestamp 1712622712
transform 1 0 1892 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6276
timestamp 1712622712
transform 1 0 1660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6277
timestamp 1712622712
transform 1 0 1580 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1712622712
transform 1 0 1612 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6279
timestamp 1712622712
transform 1 0 1532 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6280
timestamp 1712622712
transform 1 0 1428 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6281
timestamp 1712622712
transform 1 0 1412 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6282
timestamp 1712622712
transform 1 0 1412 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6283
timestamp 1712622712
transform 1 0 1340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6284
timestamp 1712622712
transform 1 0 1236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6285
timestamp 1712622712
transform 1 0 1236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6286
timestamp 1712622712
transform 1 0 1172 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6287
timestamp 1712622712
transform 1 0 1076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6288
timestamp 1712622712
transform 1 0 1180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6289
timestamp 1712622712
transform 1 0 1116 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6290
timestamp 1712622712
transform 1 0 236 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1712622712
transform 1 0 140 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6292
timestamp 1712622712
transform 1 0 244 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6293
timestamp 1712622712
transform 1 0 196 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6294
timestamp 1712622712
transform 1 0 276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6295
timestamp 1712622712
transform 1 0 140 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6296
timestamp 1712622712
transform 1 0 396 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6297
timestamp 1712622712
transform 1 0 260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6298
timestamp 1712622712
transform 1 0 428 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6299
timestamp 1712622712
transform 1 0 324 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6300
timestamp 1712622712
transform 1 0 412 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6301
timestamp 1712622712
transform 1 0 308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6302
timestamp 1712622712
transform 1 0 460 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6303
timestamp 1712622712
transform 1 0 364 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1712622712
transform 1 0 572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1712622712
transform 1 0 524 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6306
timestamp 1712622712
transform 1 0 588 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6307
timestamp 1712622712
transform 1 0 484 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6308
timestamp 1712622712
transform 1 0 884 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6309
timestamp 1712622712
transform 1 0 820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6310
timestamp 1712622712
transform 1 0 988 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6311
timestamp 1712622712
transform 1 0 988 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6312
timestamp 1712622712
transform 1 0 3404 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6313
timestamp 1712622712
transform 1 0 3396 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6314
timestamp 1712622712
transform 1 0 3356 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6315
timestamp 1712622712
transform 1 0 3372 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6316
timestamp 1712622712
transform 1 0 3372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6317
timestamp 1712622712
transform 1 0 3300 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6318
timestamp 1712622712
transform 1 0 3292 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6319
timestamp 1712622712
transform 1 0 3356 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6320
timestamp 1712622712
transform 1 0 3308 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6321
timestamp 1712622712
transform 1 0 3396 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1712622712
transform 1 0 3364 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1712622712
transform 1 0 3372 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6324
timestamp 1712622712
transform 1 0 3372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1712622712
transform 1 0 3372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1712622712
transform 1 0 3332 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6327
timestamp 1712622712
transform 1 0 3092 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6328
timestamp 1712622712
transform 1 0 3092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6329
timestamp 1712622712
transform 1 0 3196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1712622712
transform 1 0 3060 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1712622712
transform 1 0 3164 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6332
timestamp 1712622712
transform 1 0 3068 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6333
timestamp 1712622712
transform 1 0 3196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6334
timestamp 1712622712
transform 1 0 3164 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1712622712
transform 1 0 3316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6336
timestamp 1712622712
transform 1 0 3292 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6337
timestamp 1712622712
transform 1 0 3436 0 1 2655
box -2 -2 2 2
use M2_M1  M2_M1_6338
timestamp 1712622712
transform 1 0 3348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1712622712
transform 1 0 3364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6340
timestamp 1712622712
transform 1 0 3228 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6341
timestamp 1712622712
transform 1 0 3052 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6342
timestamp 1712622712
transform 1 0 3052 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6343
timestamp 1712622712
transform 1 0 3348 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6344
timestamp 1712622712
transform 1 0 3324 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_6345
timestamp 1712622712
transform 1 0 3324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6346
timestamp 1712622712
transform 1 0 3364 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6347
timestamp 1712622712
transform 1 0 3364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6348
timestamp 1712622712
transform 1 0 3324 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6349
timestamp 1712622712
transform 1 0 3324 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_6350
timestamp 1712622712
transform 1 0 3268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6351
timestamp 1712622712
transform 1 0 3428 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6352
timestamp 1712622712
transform 1 0 3428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6353
timestamp 1712622712
transform 1 0 3396 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6354
timestamp 1712622712
transform 1 0 3364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6355
timestamp 1712622712
transform 1 0 3428 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6356
timestamp 1712622712
transform 1 0 3388 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6357
timestamp 1712622712
transform 1 0 3332 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6358
timestamp 1712622712
transform 1 0 3332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6359
timestamp 1712622712
transform 1 0 3300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6360
timestamp 1712622712
transform 1 0 3284 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1712622712
transform 1 0 3356 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6362
timestamp 1712622712
transform 1 0 3300 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6363
timestamp 1712622712
transform 1 0 3380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1712622712
transform 1 0 3348 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6365
timestamp 1712622712
transform 1 0 3324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6366
timestamp 1712622712
transform 1 0 3292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6367
timestamp 1712622712
transform 1 0 3252 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6368
timestamp 1712622712
transform 1 0 3076 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6369
timestamp 1712622712
transform 1 0 2900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6370
timestamp 1712622712
transform 1 0 2868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6371
timestamp 1712622712
transform 1 0 2340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6372
timestamp 1712622712
transform 1 0 2332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6373
timestamp 1712622712
transform 1 0 2300 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_6374
timestamp 1712622712
transform 1 0 2300 0 1 1885
box -2 -2 2 2
use M2_M1  M2_M1_6375
timestamp 1712622712
transform 1 0 2244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6376
timestamp 1712622712
transform 1 0 2236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6377
timestamp 1712622712
transform 1 0 2228 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6378
timestamp 1712622712
transform 1 0 3188 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6379
timestamp 1712622712
transform 1 0 2692 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1712622712
transform 1 0 2532 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6381
timestamp 1712622712
transform 1 0 2436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6382
timestamp 1712622712
transform 1 0 2244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6383
timestamp 1712622712
transform 1 0 2164 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6384
timestamp 1712622712
transform 1 0 2092 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6385
timestamp 1712622712
transform 1 0 1780 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1712622712
transform 1 0 1612 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1712622712
transform 1 0 1468 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6388
timestamp 1712622712
transform 1 0 980 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6389
timestamp 1712622712
transform 1 0 868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6390
timestamp 1712622712
transform 1 0 2044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6391
timestamp 1712622712
transform 1 0 2028 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6392
timestamp 1712622712
transform 1 0 1980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6393
timestamp 1712622712
transform 1 0 1964 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6394
timestamp 1712622712
transform 1 0 1924 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6395
timestamp 1712622712
transform 1 0 2212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1712622712
transform 1 0 2156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6397
timestamp 1712622712
transform 1 0 2116 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6398
timestamp 1712622712
transform 1 0 2092 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1712622712
transform 1 0 2092 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6400
timestamp 1712622712
transform 1 0 1700 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6401
timestamp 1712622712
transform 1 0 2404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6402
timestamp 1712622712
transform 1 0 2380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6403
timestamp 1712622712
transform 1 0 2364 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6404
timestamp 1712622712
transform 1 0 2364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6405
timestamp 1712622712
transform 1 0 1756 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6406
timestamp 1712622712
transform 1 0 2524 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6407
timestamp 1712622712
transform 1 0 2508 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6408
timestamp 1712622712
transform 1 0 2492 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6409
timestamp 1712622712
transform 1 0 2420 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6410
timestamp 1712622712
transform 1 0 2268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6411
timestamp 1712622712
transform 1 0 1932 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6412
timestamp 1712622712
transform 1 0 2636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6413
timestamp 1712622712
transform 1 0 2612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6414
timestamp 1712622712
transform 1 0 2612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6415
timestamp 1712622712
transform 1 0 2444 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6416
timestamp 1712622712
transform 1 0 2244 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6417
timestamp 1712622712
transform 1 0 1892 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6418
timestamp 1712622712
transform 1 0 2900 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6419
timestamp 1712622712
transform 1 0 2836 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6420
timestamp 1712622712
transform 1 0 2796 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_6421
timestamp 1712622712
transform 1 0 2772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6422
timestamp 1712622712
transform 1 0 2764 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6423
timestamp 1712622712
transform 1 0 2484 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6424
timestamp 1712622712
transform 1 0 2420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6425
timestamp 1712622712
transform 1 0 1324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6426
timestamp 1712622712
transform 1 0 1316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6427
timestamp 1712622712
transform 1 0 1308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6428
timestamp 1712622712
transform 1 0 1308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6429
timestamp 1712622712
transform 1 0 1164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6430
timestamp 1712622712
transform 1 0 996 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6431
timestamp 1712622712
transform 1 0 908 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6432
timestamp 1712622712
transform 1 0 892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6433
timestamp 1712622712
transform 1 0 892 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6434
timestamp 1712622712
transform 1 0 876 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6435
timestamp 1712622712
transform 1 0 876 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6436
timestamp 1712622712
transform 1 0 868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6437
timestamp 1712622712
transform 1 0 788 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1712622712
transform 1 0 3028 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_6439
timestamp 1712622712
transform 1 0 3028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6440
timestamp 1712622712
transform 1 0 3012 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_6441
timestamp 1712622712
transform 1 0 2996 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6442
timestamp 1712622712
transform 1 0 2964 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6443
timestamp 1712622712
transform 1 0 2908 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6444
timestamp 1712622712
transform 1 0 2844 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6445
timestamp 1712622712
transform 1 0 2844 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6446
timestamp 1712622712
transform 1 0 844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6447
timestamp 1712622712
transform 1 0 748 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6448
timestamp 1712622712
transform 1 0 732 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1712622712
transform 1 0 732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6450
timestamp 1712622712
transform 1 0 708 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6451
timestamp 1712622712
transform 1 0 708 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6452
timestamp 1712622712
transform 1 0 980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6453
timestamp 1712622712
transform 1 0 796 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_6454
timestamp 1712622712
transform 1 0 756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6455
timestamp 1712622712
transform 1 0 652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6456
timestamp 1712622712
transform 1 0 636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6457
timestamp 1712622712
transform 1 0 620 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6458
timestamp 1712622712
transform 1 0 860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1712622712
transform 1 0 540 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6460
timestamp 1712622712
transform 1 0 516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6461
timestamp 1712622712
transform 1 0 468 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6462
timestamp 1712622712
transform 1 0 692 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6463
timestamp 1712622712
transform 1 0 516 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6464
timestamp 1712622712
transform 1 0 428 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6465
timestamp 1712622712
transform 1 0 388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6466
timestamp 1712622712
transform 1 0 572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6467
timestamp 1712622712
transform 1 0 468 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6468
timestamp 1712622712
transform 1 0 348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6469
timestamp 1712622712
transform 1 0 324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6470
timestamp 1712622712
transform 1 0 652 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6471
timestamp 1712622712
transform 1 0 532 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6472
timestamp 1712622712
transform 1 0 316 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6473
timestamp 1712622712
transform 1 0 276 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6474
timestamp 1712622712
transform 1 0 684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6475
timestamp 1712622712
transform 1 0 668 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6476
timestamp 1712622712
transform 1 0 588 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6477
timestamp 1712622712
transform 1 0 252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6478
timestamp 1712622712
transform 1 0 228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6479
timestamp 1712622712
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6480
timestamp 1712622712
transform 1 0 580 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6481
timestamp 1712622712
transform 1 0 548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6482
timestamp 1712622712
transform 1 0 108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1712622712
transform 1 0 84 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6484
timestamp 1712622712
transform 1 0 804 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6485
timestamp 1712622712
transform 1 0 756 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6486
timestamp 1712622712
transform 1 0 732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6487
timestamp 1712622712
transform 1 0 588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6488
timestamp 1712622712
transform 1 0 172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6489
timestamp 1712622712
transform 1 0 124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6490
timestamp 1712622712
transform 1 0 868 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6491
timestamp 1712622712
transform 1 0 852 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6492
timestamp 1712622712
transform 1 0 820 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6493
timestamp 1712622712
transform 1 0 780 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6494
timestamp 1712622712
transform 1 0 644 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6495
timestamp 1712622712
transform 1 0 532 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6496
timestamp 1712622712
transform 1 0 3076 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6497
timestamp 1712622712
transform 1 0 2988 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6498
timestamp 1712622712
transform 1 0 2908 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1712622712
transform 1 0 2900 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6500
timestamp 1712622712
transform 1 0 2868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6501
timestamp 1712622712
transform 1 0 2644 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6502
timestamp 1712622712
transform 1 0 2540 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6503
timestamp 1712622712
transform 1 0 1220 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6504
timestamp 1712622712
transform 1 0 1044 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6505
timestamp 1712622712
transform 1 0 1020 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6506
timestamp 1712622712
transform 1 0 1012 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6507
timestamp 1712622712
transform 1 0 972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6508
timestamp 1712622712
transform 1 0 964 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6509
timestamp 1712622712
transform 1 0 1268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6510
timestamp 1712622712
transform 1 0 1220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6511
timestamp 1712622712
transform 1 0 1204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6512
timestamp 1712622712
transform 1 0 1108 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6513
timestamp 1712622712
transform 1 0 1100 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6514
timestamp 1712622712
transform 1 0 1084 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6515
timestamp 1712622712
transform 1 0 1460 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6516
timestamp 1712622712
transform 1 0 1404 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6517
timestamp 1712622712
transform 1 0 1300 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6518
timestamp 1712622712
transform 1 0 1292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6519
timestamp 1712622712
transform 1 0 1268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6520
timestamp 1712622712
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6521
timestamp 1712622712
transform 1 0 1244 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6522
timestamp 1712622712
transform 1 0 1204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6523
timestamp 1712622712
transform 1 0 1516 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6524
timestamp 1712622712
transform 1 0 1484 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6525
timestamp 1712622712
transform 1 0 1460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6526
timestamp 1712622712
transform 1 0 1412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6527
timestamp 1712622712
transform 1 0 1316 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6528
timestamp 1712622712
transform 1 0 1316 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6529
timestamp 1712622712
transform 1 0 1292 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6530
timestamp 1712622712
transform 1 0 1276 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6531
timestamp 1712622712
transform 1 0 1604 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6532
timestamp 1712622712
transform 1 0 1548 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6533
timestamp 1712622712
transform 1 0 1468 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6534
timestamp 1712622712
transform 1 0 1468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6535
timestamp 1712622712
transform 1 0 1676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6536
timestamp 1712622712
transform 1 0 1676 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6537
timestamp 1712622712
transform 1 0 1668 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6538
timestamp 1712622712
transform 1 0 1668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1712622712
transform 1 0 1796 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6540
timestamp 1712622712
transform 1 0 1780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6541
timestamp 1712622712
transform 1 0 1772 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6542
timestamp 1712622712
transform 1 0 1756 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1712622712
transform 1 0 1700 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6544
timestamp 1712622712
transform 1 0 1684 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6545
timestamp 1712622712
transform 1 0 1852 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1712622712
transform 1 0 1852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6547
timestamp 1712622712
transform 1 0 1852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6548
timestamp 1712622712
transform 1 0 1844 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1712622712
transform 1 0 2148 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6550
timestamp 1712622712
transform 1 0 2100 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6551
timestamp 1712622712
transform 1 0 2084 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1712622712
transform 1 0 2076 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6553
timestamp 1712622712
transform 1 0 2052 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6554
timestamp 1712622712
transform 1 0 2052 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1712622712
transform 1 0 1980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6556
timestamp 1712622712
transform 1 0 2332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6557
timestamp 1712622712
transform 1 0 2308 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6558
timestamp 1712622712
transform 1 0 2284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6559
timestamp 1712622712
transform 1 0 2268 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6560
timestamp 1712622712
transform 1 0 2260 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1712622712
transform 1 0 2236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1712622712
transform 1 0 2180 0 1 1755
box -2 -2 2 2
use M2_M1  M2_M1_6563
timestamp 1712622712
transform 1 0 2172 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1712622712
transform 1 0 2164 0 1 1755
box -2 -2 2 2
use M2_M1  M2_M1_6565
timestamp 1712622712
transform 1 0 2068 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6566
timestamp 1712622712
transform 1 0 2852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6567
timestamp 1712622712
transform 1 0 2732 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6568
timestamp 1712622712
transform 1 0 2708 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6569
timestamp 1712622712
transform 1 0 2684 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6570
timestamp 1712622712
transform 1 0 2580 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6571
timestamp 1712622712
transform 1 0 2484 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6572
timestamp 1712622712
transform 1 0 2468 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1712622712
transform 1 0 3340 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6574
timestamp 1712622712
transform 1 0 3092 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6575
timestamp 1712622712
transform 1 0 3084 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6576
timestamp 1712622712
transform 1 0 2468 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6577
timestamp 1712622712
transform 1 0 2300 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6578
timestamp 1712622712
transform 1 0 2564 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1712622712
transform 1 0 2548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6580
timestamp 1712622712
transform 1 0 2348 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1712622712
transform 1 0 2812 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1712622712
transform 1 0 2804 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6583
timestamp 1712622712
transform 1 0 2780 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1712622712
transform 1 0 2596 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1712622712
transform 1 0 2364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6586
timestamp 1712622712
transform 1 0 2300 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1712622712
transform 1 0 2388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6588
timestamp 1712622712
transform 1 0 2340 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1712622712
transform 1 0 2204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6590
timestamp 1712622712
transform 1 0 2556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6591
timestamp 1712622712
transform 1 0 2452 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6592
timestamp 1712622712
transform 1 0 2348 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6593
timestamp 1712622712
transform 1 0 2620 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6594
timestamp 1712622712
transform 1 0 2556 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6595
timestamp 1712622712
transform 1 0 2412 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6596
timestamp 1712622712
transform 1 0 2412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6597
timestamp 1712622712
transform 1 0 2588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6598
timestamp 1712622712
transform 1 0 2564 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6599
timestamp 1712622712
transform 1 0 2356 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6600
timestamp 1712622712
transform 1 0 2340 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6601
timestamp 1712622712
transform 1 0 2252 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6602
timestamp 1712622712
transform 1 0 2468 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6603
timestamp 1712622712
transform 1 0 2244 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6604
timestamp 1712622712
transform 1 0 2236 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1712622712
transform 1 0 2220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6606
timestamp 1712622712
transform 1 0 2020 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6607
timestamp 1712622712
transform 1 0 1956 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6608
timestamp 1712622712
transform 1 0 1876 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6609
timestamp 1712622712
transform 1 0 1852 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1712622712
transform 1 0 1844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6611
timestamp 1712622712
transform 1 0 1628 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6612
timestamp 1712622712
transform 1 0 2300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6613
timestamp 1712622712
transform 1 0 2236 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6614
timestamp 1712622712
transform 1 0 1900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6615
timestamp 1712622712
transform 1 0 1868 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6616
timestamp 1712622712
transform 1 0 1556 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6617
timestamp 1712622712
transform 1 0 2220 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6618
timestamp 1712622712
transform 1 0 2180 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6619
timestamp 1712622712
transform 1 0 1780 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6620
timestamp 1712622712
transform 1 0 1572 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6621
timestamp 1712622712
transform 1 0 2140 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6622
timestamp 1712622712
transform 1 0 2068 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6623
timestamp 1712622712
transform 1 0 1676 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6624
timestamp 1712622712
transform 1 0 1516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6625
timestamp 1712622712
transform 1 0 1820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6626
timestamp 1712622712
transform 1 0 1804 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6627
timestamp 1712622712
transform 1 0 1676 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6628
timestamp 1712622712
transform 1 0 1388 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6629
timestamp 1712622712
transform 1 0 1388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6630
timestamp 1712622712
transform 1 0 1948 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6631
timestamp 1712622712
transform 1 0 1868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6632
timestamp 1712622712
transform 1 0 1780 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6633
timestamp 1712622712
transform 1 0 1588 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6634
timestamp 1712622712
transform 1 0 1396 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6635
timestamp 1712622712
transform 1 0 1308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6636
timestamp 1712622712
transform 1 0 1724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1712622712
transform 1 0 1716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6638
timestamp 1712622712
transform 1 0 1716 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_6639
timestamp 1712622712
transform 1 0 1620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6640
timestamp 1712622712
transform 1 0 1428 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6641
timestamp 1712622712
transform 1 0 1196 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6642
timestamp 1712622712
transform 1 0 1644 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6643
timestamp 1712622712
transform 1 0 1644 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6644
timestamp 1712622712
transform 1 0 1628 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6645
timestamp 1712622712
transform 1 0 1564 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6646
timestamp 1712622712
transform 1 0 1556 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6647
timestamp 1712622712
transform 1 0 1420 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6648
timestamp 1712622712
transform 1 0 1044 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6649
timestamp 1712622712
transform 1 0 1476 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6650
timestamp 1712622712
transform 1 0 1300 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6651
timestamp 1712622712
transform 1 0 780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6652
timestamp 1712622712
transform 1 0 1380 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6653
timestamp 1712622712
transform 1 0 1236 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6654
timestamp 1712622712
transform 1 0 716 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6655
timestamp 1712622712
transform 1 0 1300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6656
timestamp 1712622712
transform 1 0 1212 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6657
timestamp 1712622712
transform 1 0 1084 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6658
timestamp 1712622712
transform 1 0 676 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6659
timestamp 1712622712
transform 1 0 1204 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6660
timestamp 1712622712
transform 1 0 1172 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6661
timestamp 1712622712
transform 1 0 1052 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6662
timestamp 1712622712
transform 1 0 716 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6663
timestamp 1712622712
transform 1 0 1340 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6664
timestamp 1712622712
transform 1 0 1148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6665
timestamp 1712622712
transform 1 0 860 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6666
timestamp 1712622712
transform 1 0 764 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1712622712
transform 1 0 1220 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6668
timestamp 1712622712
transform 1 0 972 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6669
timestamp 1712622712
transform 1 0 772 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1712622712
transform 1 0 700 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6671
timestamp 1712622712
transform 1 0 1124 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6672
timestamp 1712622712
transform 1 0 836 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6673
timestamp 1712622712
transform 1 0 652 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6674
timestamp 1712622712
transform 1 0 564 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6675
timestamp 1712622712
transform 1 0 564 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6676
timestamp 1712622712
transform 1 0 1012 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6677
timestamp 1712622712
transform 1 0 820 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6678
timestamp 1712622712
transform 1 0 732 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6679
timestamp 1712622712
transform 1 0 668 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6680
timestamp 1712622712
transform 1 0 668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6681
timestamp 1712622712
transform 1 0 748 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6682
timestamp 1712622712
transform 1 0 724 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6683
timestamp 1712622712
transform 1 0 540 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6684
timestamp 1712622712
transform 1 0 540 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6685
timestamp 1712622712
transform 1 0 500 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6686
timestamp 1712622712
transform 1 0 684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6687
timestamp 1712622712
transform 1 0 684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6688
timestamp 1712622712
transform 1 0 508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6689
timestamp 1712622712
transform 1 0 500 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6690
timestamp 1712622712
transform 1 0 476 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6691
timestamp 1712622712
transform 1 0 644 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6692
timestamp 1712622712
transform 1 0 628 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6693
timestamp 1712622712
transform 1 0 596 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6694
timestamp 1712622712
transform 1 0 548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6695
timestamp 1712622712
transform 1 0 532 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6696
timestamp 1712622712
transform 1 0 492 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6697
timestamp 1712622712
transform 1 0 716 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6698
timestamp 1712622712
transform 1 0 684 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6699
timestamp 1712622712
transform 1 0 564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6700
timestamp 1712622712
transform 1 0 540 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6701
timestamp 1712622712
transform 1 0 540 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6702
timestamp 1712622712
transform 1 0 508 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6703
timestamp 1712622712
transform 1 0 644 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6704
timestamp 1712622712
transform 1 0 644 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6705
timestamp 1712622712
transform 1 0 612 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6706
timestamp 1712622712
transform 1 0 740 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6707
timestamp 1712622712
transform 1 0 700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6708
timestamp 1712622712
transform 1 0 900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6709
timestamp 1712622712
transform 1 0 884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6710
timestamp 1712622712
transform 1 0 868 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6711
timestamp 1712622712
transform 1 0 996 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6712
timestamp 1712622712
transform 1 0 980 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6713
timestamp 1712622712
transform 1 0 892 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6714
timestamp 1712622712
transform 1 0 3412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6715
timestamp 1712622712
transform 1 0 3380 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_6716
timestamp 1712622712
transform 1 0 3300 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6717
timestamp 1712622712
transform 1 0 3260 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1712622712
transform 1 0 3412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6719
timestamp 1712622712
transform 1 0 2092 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6720
timestamp 1712622712
transform 1 0 1916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6721
timestamp 1712622712
transform 1 0 3124 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6722
timestamp 1712622712
transform 1 0 3116 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6723
timestamp 1712622712
transform 1 0 3108 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6724
timestamp 1712622712
transform 1 0 2900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1712622712
transform 1 0 2820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6726
timestamp 1712622712
transform 1 0 2692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6727
timestamp 1712622712
transform 1 0 2612 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6728
timestamp 1712622712
transform 1 0 2604 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1712622712
transform 1 0 3204 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1712622712
transform 1 0 3092 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1712622712
transform 1 0 3108 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1712622712
transform 1 0 2876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1712622712
transform 1 0 3140 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1712622712
transform 1 0 3028 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1712622712
transform 1 0 3028 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1712622712
transform 1 0 2988 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1712622712
transform 1 0 2988 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1712622712
transform 1 0 2916 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1712622712
transform 1 0 2884 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1712622712
transform 1 0 2852 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1712622712
transform 1 0 3140 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1712622712
transform 1 0 2924 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1712622712
transform 1 0 2828 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1712622712
transform 1 0 3060 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1712622712
transform 1 0 2996 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1712622712
transform 1 0 2988 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1712622712
transform 1 0 2964 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1712622712
transform 1 0 2964 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1712622712
transform 1 0 2852 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1712622712
transform 1 0 2812 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1712622712
transform 1 0 2836 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1712622712
transform 1 0 2772 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1712622712
transform 1 0 1412 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1712622712
transform 1 0 1404 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1712622712
transform 1 0 1380 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1712622712
transform 1 0 2892 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1712622712
transform 1 0 2804 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1712622712
transform 1 0 1524 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1712622712
transform 1 0 1420 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1712622712
transform 1 0 1364 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1712622712
transform 1 0 3268 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1712622712
transform 1 0 3268 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1712622712
transform 1 0 3180 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1712622712
transform 1 0 3180 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1712622712
transform 1 0 2980 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1712622712
transform 1 0 2980 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1712622712
transform 1 0 2852 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1712622712
transform 1 0 2852 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1712622712
transform 1 0 2828 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1712622712
transform 1 0 2828 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1712622712
transform 1 0 2748 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1712622712
transform 1 0 2748 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1712622712
transform 1 0 2684 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1712622712
transform 1 0 2676 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1712622712
transform 1 0 2588 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1712622712
transform 1 0 2572 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1712622712
transform 1 0 2564 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1712622712
transform 1 0 2412 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1712622712
transform 1 0 2164 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1712622712
transform 1 0 2164 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1712622712
transform 1 0 1964 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1712622712
transform 1 0 1380 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1712622712
transform 1 0 1364 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1712622712
transform 1 0 1364 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1712622712
transform 1 0 1300 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1712622712
transform 1 0 1292 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1712622712
transform 1 0 1292 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1712622712
transform 1 0 1084 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1712622712
transform 1 0 1076 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1712622712
transform 1 0 1028 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1712622712
transform 1 0 1004 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1712622712
transform 1 0 1004 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1712622712
transform 1 0 748 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1712622712
transform 1 0 716 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1712622712
transform 1 0 708 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1712622712
transform 1 0 700 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1712622712
transform 1 0 684 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1712622712
transform 1 0 668 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1712622712
transform 1 0 668 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1712622712
transform 1 0 644 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1712622712
transform 1 0 596 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1712622712
transform 1 0 596 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1712622712
transform 1 0 3188 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1712622712
transform 1 0 2988 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1712622712
transform 1 0 2964 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1712622712
transform 1 0 2684 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1712622712
transform 1 0 2628 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1712622712
transform 1 0 3100 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1712622712
transform 1 0 2956 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1712622712
transform 1 0 2932 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1712622712
transform 1 0 2868 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1712622712
transform 1 0 3004 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1712622712
transform 1 0 2932 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1712622712
transform 1 0 2876 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1712622712
transform 1 0 2892 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1712622712
transform 1 0 2788 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1712622712
transform 1 0 3404 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1712622712
transform 1 0 3300 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1712622712
transform 1 0 3292 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1712622712
transform 1 0 3260 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1712622712
transform 1 0 3420 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1712622712
transform 1 0 3348 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1712622712
transform 1 0 3348 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1712622712
transform 1 0 3284 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1712622712
transform 1 0 2980 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1712622712
transform 1 0 2916 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1712622712
transform 1 0 2900 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1712622712
transform 1 0 2828 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1712622712
transform 1 0 2692 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1712622712
transform 1 0 2564 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1712622712
transform 1 0 2772 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1712622712
transform 1 0 2724 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1712622712
transform 1 0 2820 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1712622712
transform 1 0 2716 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1712622712
transform 1 0 2508 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1712622712
transform 1 0 2404 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1712622712
transform 1 0 2148 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1712622712
transform 1 0 2028 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1712622712
transform 1 0 2236 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1712622712
transform 1 0 2132 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1712622712
transform 1 0 1924 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1712622712
transform 1 0 1852 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1712622712
transform 1 0 1564 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1712622712
transform 1 0 1500 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1712622712
transform 1 0 1444 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1712622712
transform 1 0 1332 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1712622712
transform 1 0 1468 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1712622712
transform 1 0 1348 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1712622712
transform 1 0 1292 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1712622712
transform 1 0 1228 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1712622712
transform 1 0 1148 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1712622712
transform 1 0 1020 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1712622712
transform 1 0 228 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1712622712
transform 1 0 84 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1712622712
transform 1 0 3284 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1712622712
transform 1 0 3276 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1712622712
transform 1 0 3428 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1712622712
transform 1 0 3292 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1712622712
transform 1 0 3436 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1712622712
transform 1 0 3388 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1712622712
transform 1 0 3404 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1712622712
transform 1 0 3332 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1712622712
transform 1 0 3052 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1712622712
transform 1 0 2836 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1712622712
transform 1 0 3364 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1712622712
transform 1 0 3348 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1712622712
transform 1 0 3324 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1712622712
transform 1 0 3324 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1712622712
transform 1 0 3060 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1712622712
transform 1 0 2980 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1712622712
transform 1 0 2756 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1712622712
transform 1 0 2668 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1712622712
transform 1 0 2948 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1712622712
transform 1 0 2884 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1712622712
transform 1 0 3044 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1712622712
transform 1 0 2828 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1712622712
transform 1 0 2844 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1712622712
transform 1 0 2740 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1712622712
transform 1 0 2652 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1712622712
transform 1 0 2596 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1712622712
transform 1 0 2460 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1712622712
transform 1 0 2388 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1712622712
transform 1 0 2260 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1712622712
transform 1 0 2220 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1712622712
transform 1 0 2060 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1712622712
transform 1 0 2036 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1712622712
transform 1 0 1860 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1712622712
transform 1 0 1836 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1712622712
transform 1 0 1484 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1712622712
transform 1 0 1460 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1712622712
transform 1 0 1444 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1712622712
transform 1 0 1356 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1712622712
transform 1 0 1188 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1712622712
transform 1 0 1140 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1712622712
transform 1 0 1060 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1712622712
transform 1 0 956 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1712622712
transform 1 0 764 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1712622712
transform 1 0 628 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1712622712
transform 1 0 180 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1712622712
transform 1 0 84 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1712622712
transform 1 0 724 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1712622712
transform 1 0 612 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1712622712
transform 1 0 836 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1712622712
transform 1 0 716 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1712622712
transform 1 0 948 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1712622712
transform 1 0 868 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1712622712
transform 1 0 1244 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1712622712
transform 1 0 1148 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1712622712
transform 1 0 2972 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1712622712
transform 1 0 2924 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1712622712
transform 1 0 3036 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1712622712
transform 1 0 2876 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1712622712
transform 1 0 2548 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1712622712
transform 1 0 2444 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1712622712
transform 1 0 2436 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1712622712
transform 1 0 2204 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1712622712
transform 1 0 2308 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1712622712
transform 1 0 2260 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1712622712
transform 1 0 2348 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1712622712
transform 1 0 2268 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1712622712
transform 1 0 1996 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1712622712
transform 1 0 1828 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1712622712
transform 1 0 1772 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1712622712
transform 1 0 1716 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1712622712
transform 1 0 1476 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1712622712
transform 1 0 1436 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1712622712
transform 1 0 1308 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1712622712
transform 1 0 1244 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1712622712
transform 1 0 1084 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1712622712
transform 1 0 1020 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1712622712
transform 1 0 988 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1712622712
transform 1 0 860 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1712622712
transform 1 0 3348 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1712622712
transform 1 0 3196 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1712622712
transform 1 0 3180 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1712622712
transform 1 0 3172 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1712622712
transform 1 0 3124 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1712622712
transform 1 0 3124 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1712622712
transform 1 0 3100 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1712622712
transform 1 0 3244 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1712622712
transform 1 0 3196 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1712622712
transform 1 0 3164 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1712622712
transform 1 0 3148 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1712622712
transform 1 0 3148 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1712622712
transform 1 0 3116 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1712622712
transform 1 0 3108 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1712622712
transform 1 0 3100 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1712622712
transform 1 0 3036 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1712622712
transform 1 0 3012 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1712622712
transform 1 0 3012 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1712622712
transform 1 0 2964 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1712622712
transform 1 0 2908 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1712622712
transform 1 0 2844 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1712622712
transform 1 0 2948 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1712622712
transform 1 0 2876 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1712622712
transform 1 0 2828 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1712622712
transform 1 0 2828 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1712622712
transform 1 0 3396 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1712622712
transform 1 0 3188 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1712622712
transform 1 0 3300 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1712622712
transform 1 0 3252 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1712622712
transform 1 0 3148 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1712622712
transform 1 0 3380 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1712622712
transform 1 0 3340 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1712622712
transform 1 0 3428 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1712622712
transform 1 0 3364 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1712622712
transform 1 0 3420 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1712622712
transform 1 0 3316 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1712622712
transform 1 0 3308 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1712622712
transform 1 0 3212 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1712622712
transform 1 0 3188 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1712622712
transform 1 0 3148 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1712622712
transform 1 0 3068 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1712622712
transform 1 0 3028 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1712622712
transform 1 0 2996 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1712622712
transform 1 0 2892 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1712622712
transform 1 0 3332 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1712622712
transform 1 0 3300 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1712622712
transform 1 0 3172 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1712622712
transform 1 0 3148 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1712622712
transform 1 0 3420 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1712622712
transform 1 0 3300 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1712622712
transform 1 0 3276 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1712622712
transform 1 0 3276 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1712622712
transform 1 0 3164 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1712622712
transform 1 0 3188 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1712622712
transform 1 0 3100 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1712622712
transform 1 0 3036 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1712622712
transform 1 0 3196 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1712622712
transform 1 0 3156 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1712622712
transform 1 0 3252 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1712622712
transform 1 0 3172 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1712622712
transform 1 0 2676 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1712622712
transform 1 0 2604 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1712622712
transform 1 0 2588 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1712622712
transform 1 0 2404 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1712622712
transform 1 0 1668 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1712622712
transform 1 0 1668 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1712622712
transform 1 0 1452 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1712622712
transform 1 0 1444 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1712622712
transform 1 0 1260 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1712622712
transform 1 0 3396 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1712622712
transform 1 0 3276 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1712622712
transform 1 0 3260 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1712622712
transform 1 0 3188 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1712622712
transform 1 0 3180 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1712622712
transform 1 0 3268 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1712622712
transform 1 0 3164 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1712622712
transform 1 0 3068 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1712622712
transform 1 0 3068 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1712622712
transform 1 0 2956 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1712622712
transform 1 0 3284 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1712622712
transform 1 0 3236 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1712622712
transform 1 0 3124 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1712622712
transform 1 0 3068 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1712622712
transform 1 0 3012 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1712622712
transform 1 0 2788 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1712622712
transform 1 0 2756 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1712622712
transform 1 0 2756 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1712622712
transform 1 0 2684 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1712622712
transform 1 0 2644 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1712622712
transform 1 0 2644 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1712622712
transform 1 0 2612 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1712622712
transform 1 0 2612 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1712622712
transform 1 0 2420 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1712622712
transform 1 0 2388 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1712622712
transform 1 0 2388 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1712622712
transform 1 0 2284 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1712622712
transform 1 0 2284 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1712622712
transform 1 0 2252 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1712622712
transform 1 0 2252 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1712622712
transform 1 0 2044 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1712622712
transform 1 0 2044 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1712622712
transform 1 0 1916 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1712622712
transform 1 0 1908 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1712622712
transform 1 0 1820 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1712622712
transform 1 0 1748 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1712622712
transform 1 0 1748 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1712622712
transform 1 0 1684 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1712622712
transform 1 0 1380 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1712622712
transform 1 0 1324 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1712622712
transform 1 0 1164 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1712622712
transform 1 0 1164 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1712622712
transform 1 0 1044 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1712622712
transform 1 0 1028 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1712622712
transform 1 0 852 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1712622712
transform 1 0 828 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1712622712
transform 1 0 796 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1712622712
transform 1 0 2660 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1712622712
transform 1 0 2580 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1712622712
transform 1 0 2540 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1712622712
transform 1 0 2540 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1712622712
transform 1 0 2420 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1712622712
transform 1 0 2340 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1712622712
transform 1 0 2140 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1712622712
transform 1 0 2140 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1712622712
transform 1 0 1588 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1712622712
transform 1 0 1588 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1712622712
transform 1 0 1564 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1712622712
transform 1 0 1556 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1712622712
transform 1 0 1484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1712622712
transform 1 0 1484 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1712622712
transform 1 0 1476 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1712622712
transform 1 0 1452 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1712622712
transform 1 0 1396 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1712622712
transform 1 0 1340 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1712622712
transform 1 0 1300 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1712622712
transform 1 0 1020 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1712622712
transform 1 0 972 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1712622712
transform 1 0 964 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1712622712
transform 1 0 932 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1712622712
transform 1 0 932 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1712622712
transform 1 0 1452 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1712622712
transform 1 0 1156 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1712622712
transform 1 0 2860 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1712622712
transform 1 0 2772 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1712622712
transform 1 0 3028 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1712622712
transform 1 0 2932 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1712622712
transform 1 0 3380 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1712622712
transform 1 0 3332 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1712622712
transform 1 0 2948 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1712622712
transform 1 0 2932 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1712622712
transform 1 0 2868 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1712622712
transform 1 0 2844 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1712622712
transform 1 0 2772 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1712622712
transform 1 0 2748 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1712622712
transform 1 0 1500 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1712622712
transform 1 0 1452 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1712622712
transform 1 0 2540 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1712622712
transform 1 0 2452 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1712622712
transform 1 0 2452 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1712622712
transform 1 0 2420 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1712622712
transform 1 0 2372 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1712622712
transform 1 0 2300 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1712622712
transform 1 0 2300 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1712622712
transform 1 0 2220 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1712622712
transform 1 0 2060 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1712622712
transform 1 0 2060 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1712622712
transform 1 0 1980 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1712622712
transform 1 0 1924 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1712622712
transform 1 0 1892 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1712622712
transform 1 0 1812 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1712622712
transform 1 0 1700 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1712622712
transform 1 0 1628 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1712622712
transform 1 0 2940 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1712622712
transform 1 0 2884 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1712622712
transform 1 0 2948 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1712622712
transform 1 0 2836 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1712622712
transform 1 0 2796 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1712622712
transform 1 0 1020 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1712622712
transform 1 0 924 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1712622712
transform 1 0 868 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1712622712
transform 1 0 1268 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1712622712
transform 1 0 1060 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1712622712
transform 1 0 836 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1712622712
transform 1 0 2004 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1712622712
transform 1 0 1932 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1712622712
transform 1 0 1868 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1712622712
transform 1 0 1740 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1712622712
transform 1 0 2700 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1712622712
transform 1 0 2652 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1712622712
transform 1 0 1476 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1712622712
transform 1 0 1420 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1712622712
transform 1 0 772 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1712622712
transform 1 0 692 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1712622712
transform 1 0 628 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1712622712
transform 1 0 1748 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1712622712
transform 1 0 1644 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1712622712
transform 1 0 3036 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1712622712
transform 1 0 2932 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1712622712
transform 1 0 2844 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1712622712
transform 1 0 2844 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1712622712
transform 1 0 2796 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1712622712
transform 1 0 2620 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1712622712
transform 1 0 2620 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1712622712
transform 1 0 2420 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1712622712
transform 1 0 2404 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1712622712
transform 1 0 2396 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1712622712
transform 1 0 1652 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1712622712
transform 1 0 1556 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1712622712
transform 1 0 1524 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1712622712
transform 1 0 1460 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1712622712
transform 1 0 1900 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1712622712
transform 1 0 1796 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1712622712
transform 1 0 2652 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1712622712
transform 1 0 2564 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1712622712
transform 1 0 2468 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1712622712
transform 1 0 2468 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1712622712
transform 1 0 2764 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1712622712
transform 1 0 2676 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1712622712
transform 1 0 1092 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1712622712
transform 1 0 876 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1712622712
transform 1 0 1396 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1712622712
transform 1 0 1164 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1712622712
transform 1 0 2660 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1712622712
transform 1 0 1564 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1712622712
transform 1 0 1540 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1712622712
transform 1 0 1540 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1712622712
transform 1 0 2980 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1712622712
transform 1 0 2724 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1712622712
transform 1 0 1916 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1712622712
transform 1 0 1524 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1712622712
transform 1 0 1380 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1712622712
transform 1 0 1324 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1712622712
transform 1 0 1324 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1712622712
transform 1 0 1276 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1712622712
transform 1 0 1188 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1712622712
transform 1 0 2980 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1712622712
transform 1 0 2900 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1712622712
transform 1 0 2844 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1712622712
transform 1 0 2804 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1712622712
transform 1 0 740 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1712622712
transform 1 0 708 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1712622712
transform 1 0 1612 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1712622712
transform 1 0 1556 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1712622712
transform 1 0 1524 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1712622712
transform 1 0 2372 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1712622712
transform 1 0 2348 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1712622712
transform 1 0 908 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1712622712
transform 1 0 740 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1712622712
transform 1 0 692 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1712622712
transform 1 0 1588 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1712622712
transform 1 0 1516 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1712622712
transform 1 0 1364 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1712622712
transform 1 0 1364 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1712622712
transform 1 0 1276 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1712622712
transform 1 0 2780 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1712622712
transform 1 0 2740 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1712622712
transform 1 0 1708 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1712622712
transform 1 0 3076 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1712622712
transform 1 0 2996 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1712622712
transform 1 0 2332 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1712622712
transform 1 0 2156 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1712622712
transform 1 0 1420 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1712622712
transform 1 0 1364 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1712622712
transform 1 0 1324 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1712622712
transform 1 0 1244 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1712622712
transform 1 0 1084 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1712622712
transform 1 0 1052 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1712622712
transform 1 0 1092 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1712622712
transform 1 0 1004 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1712622712
transform 1 0 1004 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1712622712
transform 1 0 812 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1712622712
transform 1 0 812 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1712622712
transform 1 0 668 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1712622712
transform 1 0 1956 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1712622712
transform 1 0 1900 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1712622712
transform 1 0 1900 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1712622712
transform 1 0 1852 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1712622712
transform 1 0 1820 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1712622712
transform 1 0 1812 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1712622712
transform 1 0 2868 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1712622712
transform 1 0 2852 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1712622712
transform 1 0 2756 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1712622712
transform 1 0 2748 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1712622712
transform 1 0 2564 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1712622712
transform 1 0 2540 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1712622712
transform 1 0 2540 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1712622712
transform 1 0 1100 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1712622712
transform 1 0 900 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1712622712
transform 1 0 708 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1712622712
transform 1 0 1820 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1712622712
transform 1 0 1740 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1712622712
transform 1 0 1740 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1712622712
transform 1 0 1460 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1712622712
transform 1 0 2700 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1712622712
transform 1 0 2676 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1712622712
transform 1 0 2596 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1712622712
transform 1 0 2740 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1712622712
transform 1 0 2628 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1712622712
transform 1 0 1580 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1712622712
transform 1 0 1524 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1712622712
transform 1 0 3372 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1712622712
transform 1 0 3324 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1712622712
transform 1 0 3252 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1712622712
transform 1 0 3148 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1712622712
transform 1 0 3092 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1712622712
transform 1 0 2924 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1712622712
transform 1 0 2924 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1712622712
transform 1 0 2868 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1712622712
transform 1 0 2740 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1712622712
transform 1 0 2764 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1712622712
transform 1 0 2708 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1712622712
transform 1 0 3020 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1712622712
transform 1 0 2740 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1712622712
transform 1 0 2676 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1712622712
transform 1 0 2692 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1712622712
transform 1 0 2556 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1712622712
transform 1 0 2428 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1712622712
transform 1 0 2396 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1712622712
transform 1 0 3156 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1712622712
transform 1 0 2756 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1712622712
transform 1 0 2676 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1712622712
transform 1 0 2652 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1712622712
transform 1 0 2620 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1712622712
transform 1 0 2580 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1712622712
transform 1 0 2580 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1712622712
transform 1 0 2500 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1712622712
transform 1 0 1596 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1712622712
transform 1 0 1588 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1712622712
transform 1 0 1380 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1712622712
transform 1 0 1372 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1712622712
transform 1 0 1348 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1712622712
transform 1 0 1188 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1712622712
transform 1 0 1156 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1712622712
transform 1 0 1044 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1712622712
transform 1 0 1028 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1712622712
transform 1 0 1028 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1712622712
transform 1 0 1020 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1712622712
transform 1 0 900 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1712622712
transform 1 0 884 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1712622712
transform 1 0 884 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1712622712
transform 1 0 836 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1712622712
transform 1 0 836 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1712622712
transform 1 0 644 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1712622712
transform 1 0 532 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1712622712
transform 1 0 1244 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1712622712
transform 1 0 1012 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1712622712
transform 1 0 1012 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1712622712
transform 1 0 884 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1712622712
transform 1 0 852 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1712622712
transform 1 0 844 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1712622712
transform 1 0 516 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1712622712
transform 1 0 452 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1712622712
transform 1 0 436 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1712622712
transform 1 0 236 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1712622712
transform 1 0 228 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1712622712
transform 1 0 228 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1712622712
transform 1 0 220 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1712622712
transform 1 0 156 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1712622712
transform 1 0 148 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1712622712
transform 1 0 132 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1712622712
transform 1 0 1740 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1712622712
transform 1 0 1628 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1712622712
transform 1 0 1620 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1712622712
transform 1 0 1580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1712622712
transform 1 0 1396 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1712622712
transform 1 0 2092 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1712622712
transform 1 0 2068 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1712622712
transform 1 0 2060 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1712622712
transform 1 0 2036 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1712622712
transform 1 0 2516 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1712622712
transform 1 0 2508 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1712622712
transform 1 0 2492 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1712622712
transform 1 0 2492 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1712622712
transform 1 0 2380 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1712622712
transform 1 0 1108 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1712622712
transform 1 0 1108 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1712622712
transform 1 0 1060 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1712622712
transform 1 0 1372 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1712622712
transform 1 0 1284 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1712622712
transform 1 0 676 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1712622712
transform 1 0 676 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1712622712
transform 1 0 620 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1712622712
transform 1 0 580 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1712622712
transform 1 0 1332 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1712622712
transform 1 0 1012 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1712622712
transform 1 0 884 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1712622712
transform 1 0 772 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1712622712
transform 1 0 668 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1712622712
transform 1 0 3132 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1712622712
transform 1 0 3068 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1712622712
transform 1 0 3068 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1712622712
transform 1 0 2900 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1712622712
transform 1 0 2724 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1712622712
transform 1 0 2276 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1712622712
transform 1 0 1932 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1712622712
transform 1 0 1900 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1712622712
transform 1 0 2652 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1712622712
transform 1 0 2628 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1712622712
transform 1 0 2460 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1712622712
transform 1 0 2452 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1712622712
transform 1 0 2356 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1712622712
transform 1 0 2348 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1712622712
transform 1 0 2284 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1712622712
transform 1 0 1300 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1712622712
transform 1 0 1300 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1712622712
transform 1 0 1244 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1712622712
transform 1 0 1292 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1712622712
transform 1 0 1236 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1712622712
transform 1 0 1196 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1712622712
transform 1 0 1196 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1712622712
transform 1 0 1164 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1712622712
transform 1 0 1140 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1712622712
transform 1 0 980 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1712622712
transform 1 0 964 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1712622712
transform 1 0 900 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1712622712
transform 1 0 708 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1712622712
transform 1 0 708 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1712622712
transform 1 0 604 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1712622712
transform 1 0 596 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1712622712
transform 1 0 548 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1712622712
transform 1 0 532 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1712622712
transform 1 0 500 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1712622712
transform 1 0 3004 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1712622712
transform 1 0 2660 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1712622712
transform 1 0 2436 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1712622712
transform 1 0 2380 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1712622712
transform 1 0 2244 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1712622712
transform 1 0 2676 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1712622712
transform 1 0 2484 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1712622712
transform 1 0 2484 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1712622712
transform 1 0 1236 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1712622712
transform 1 0 1324 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1712622712
transform 1 0 1268 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1712622712
transform 1 0 1196 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1712622712
transform 1 0 1164 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1712622712
transform 1 0 1612 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1712622712
transform 1 0 932 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1712622712
transform 1 0 876 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1712622712
transform 1 0 748 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1712622712
transform 1 0 748 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1712622712
transform 1 0 732 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1712622712
transform 1 0 668 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1712622712
transform 1 0 324 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1712622712
transform 1 0 324 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1712622712
transform 1 0 276 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1712622712
transform 1 0 604 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1712622712
transform 1 0 564 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1712622712
transform 1 0 188 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1712622712
transform 1 0 100 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1712622712
transform 1 0 2516 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1712622712
transform 1 0 2484 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1712622712
transform 1 0 2484 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1712622712
transform 1 0 1092 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1712622712
transform 1 0 1076 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1712622712
transform 1 0 972 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1712622712
transform 1 0 940 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1712622712
transform 1 0 1228 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1712622712
transform 1 0 836 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1712622712
transform 1 0 828 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1712622712
transform 1 0 780 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1712622712
transform 1 0 780 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1712622712
transform 1 0 116 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1712622712
transform 1 0 116 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1712622712
transform 1 0 100 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1712622712
transform 1 0 572 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1712622712
transform 1 0 532 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1712622712
transform 1 0 420 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1712622712
transform 1 0 412 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1712622712
transform 1 0 412 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1712622712
transform 1 0 412 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1712622712
transform 1 0 356 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1712622712
transform 1 0 356 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1712622712
transform 1 0 340 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1712622712
transform 1 0 340 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1712622712
transform 1 0 540 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1712622712
transform 1 0 540 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1712622712
transform 1 0 516 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1712622712
transform 1 0 516 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1712622712
transform 1 0 436 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1712622712
transform 1 0 428 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1712622712
transform 1 0 388 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1712622712
transform 1 0 2052 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1712622712
transform 1 0 2020 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1712622712
transform 1 0 2012 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1712622712
transform 1 0 2004 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1712622712
transform 1 0 1780 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1712622712
transform 1 0 1556 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1712622712
transform 1 0 1500 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1712622712
transform 1 0 1284 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1712622712
transform 1 0 1244 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1712622712
transform 1 0 1212 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1712622712
transform 1 0 2924 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1712622712
transform 1 0 2892 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1712622712
transform 1 0 2404 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1712622712
transform 1 0 2236 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1712622712
transform 1 0 2076 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1712622712
transform 1 0 2020 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1712622712
transform 1 0 2660 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1712622712
transform 1 0 2572 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1712622712
transform 1 0 2548 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1712622712
transform 1 0 2540 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1712622712
transform 1 0 2540 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1712622712
transform 1 0 1404 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1712622712
transform 1 0 1404 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1712622712
transform 1 0 1220 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1712622712
transform 1 0 1212 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1712622712
transform 1 0 1172 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1712622712
transform 1 0 1156 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1712622712
transform 1 0 1148 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1712622712
transform 1 0 1556 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1712622712
transform 1 0 1532 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1712622712
transform 1 0 1260 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1712622712
transform 1 0 1260 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1712622712
transform 1 0 1220 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1712622712
transform 1 0 1180 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1712622712
transform 1 0 1180 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1712622712
transform 1 0 828 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1712622712
transform 1 0 820 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1712622712
transform 1 0 660 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1712622712
transform 1 0 748 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1712622712
transform 1 0 740 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1712622712
transform 1 0 684 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1712622712
transform 1 0 676 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1712622712
transform 1 0 668 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1712622712
transform 1 0 508 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1712622712
transform 1 0 492 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1712622712
transform 1 0 476 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1712622712
transform 1 0 476 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1712622712
transform 1 0 292 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1712622712
transform 1 0 292 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1712622712
transform 1 0 284 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1712622712
transform 1 0 228 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1712622712
transform 1 0 1052 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1712622712
transform 1 0 892 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1712622712
transform 1 0 844 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1712622712
transform 1 0 844 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1712622712
transform 1 0 780 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1712622712
transform 1 0 516 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1712622712
transform 1 0 436 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1712622712
transform 1 0 692 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1712622712
transform 1 0 500 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1712622712
transform 1 0 484 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1712622712
transform 1 0 388 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1712622712
transform 1 0 292 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1712622712
transform 1 0 796 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1712622712
transform 1 0 772 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1712622712
transform 1 0 444 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1712622712
transform 1 0 340 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1712622712
transform 1 0 260 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1712622712
transform 1 0 2644 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1712622712
transform 1 0 2388 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1712622712
transform 1 0 3020 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1712622712
transform 1 0 2660 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1712622712
transform 1 0 2620 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1712622712
transform 1 0 2396 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1712622712
transform 1 0 2372 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1712622712
transform 1 0 2532 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1712622712
transform 1 0 2524 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1712622712
transform 1 0 2516 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1712622712
transform 1 0 2444 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1712622712
transform 1 0 2444 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1712622712
transform 1 0 2428 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1712622712
transform 1 0 2420 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1712622712
transform 1 0 1564 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1712622712
transform 1 0 1124 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1712622712
transform 1 0 1116 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1712622712
transform 1 0 1404 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1712622712
transform 1 0 828 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1712622712
transform 1 0 820 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1712622712
transform 1 0 644 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1712622712
transform 1 0 596 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1712622712
transform 1 0 492 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1712622712
transform 1 0 380 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1712622712
transform 1 0 260 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1712622712
transform 1 0 196 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1712622712
transform 1 0 188 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1712622712
transform 1 0 172 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1712622712
transform 1 0 92 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1712622712
transform 1 0 532 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1712622712
transform 1 0 460 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1712622712
transform 1 0 412 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1712622712
transform 1 0 1300 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1712622712
transform 1 0 1052 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1712622712
transform 1 0 1052 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1712622712
transform 1 0 572 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1712622712
transform 1 0 556 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1712622712
transform 1 0 548 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1712622712
transform 1 0 460 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1712622712
transform 1 0 460 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1712622712
transform 1 0 412 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1712622712
transform 1 0 1196 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1712622712
transform 1 0 996 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1712622712
transform 1 0 1308 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1712622712
transform 1 0 1300 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1712622712
transform 1 0 1228 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1712622712
transform 1 0 1220 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1712622712
transform 1 0 1060 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1712622712
transform 1 0 964 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1712622712
transform 1 0 3036 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1712622712
transform 1 0 3036 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1712622712
transform 1 0 3004 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1712622712
transform 1 0 2972 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1712622712
transform 1 0 2748 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1712622712
transform 1 0 2236 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1712622712
transform 1 0 2124 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1712622712
transform 1 0 2116 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1712622712
transform 1 0 2076 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1712622712
transform 1 0 2020 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1712622712
transform 1 0 2020 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1712622712
transform 1 0 1988 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1712622712
transform 1 0 1940 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1712622712
transform 1 0 2660 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1712622712
transform 1 0 2596 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1712622712
transform 1 0 2540 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1712622712
transform 1 0 2420 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1712622712
transform 1 0 2372 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1712622712
transform 1 0 1860 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1712622712
transform 1 0 1820 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1712622712
transform 1 0 1820 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1712622712
transform 1 0 1620 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1712622712
transform 1 0 1572 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1712622712
transform 1 0 2636 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1712622712
transform 1 0 2604 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1712622712
transform 1 0 2572 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1712622712
transform 1 0 2572 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1712622712
transform 1 0 2540 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1712622712
transform 1 0 2444 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1712622712
transform 1 0 1372 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1712622712
transform 1 0 1764 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1712622712
transform 1 0 1668 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1712622712
transform 1 0 1660 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1712622712
transform 1 0 1364 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1712622712
transform 1 0 1260 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1712622712
transform 1 0 1524 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1712622712
transform 1 0 1068 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1712622712
transform 1 0 852 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1712622712
transform 1 0 612 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1712622712
transform 1 0 580 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1712622712
transform 1 0 508 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1712622712
transform 1 0 260 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1712622712
transform 1 0 164 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1712622712
transform 1 0 2084 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1712622712
transform 1 0 924 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1712622712
transform 1 0 468 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1712622712
transform 1 0 444 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1712622712
transform 1 0 404 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1712622712
transform 1 0 396 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1712622712
transform 1 0 396 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1712622712
transform 1 0 356 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1712622712
transform 1 0 524 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1712622712
transform 1 0 468 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1712622712
transform 1 0 340 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1712622712
transform 1 0 332 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1712622712
transform 1 0 2620 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1712622712
transform 1 0 2612 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1712622712
transform 1 0 2580 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1712622712
transform 1 0 2572 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1712622712
transform 1 0 2380 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1712622712
transform 1 0 2380 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1712622712
transform 1 0 2332 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1712622712
transform 1 0 2300 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1712622712
transform 1 0 2292 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1712622712
transform 1 0 2276 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1712622712
transform 1 0 2260 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1712622712
transform 1 0 2468 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1712622712
transform 1 0 2428 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1712622712
transform 1 0 2388 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1712622712
transform 1 0 2388 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1712622712
transform 1 0 1892 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1712622712
transform 1 0 2652 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1712622712
transform 1 0 2500 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1712622712
transform 1 0 2436 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1712622712
transform 1 0 2412 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1712622712
transform 1 0 2412 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1712622712
transform 1 0 2884 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1712622712
transform 1 0 2204 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1712622712
transform 1 0 1708 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1712622712
transform 1 0 1708 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1712622712
transform 1 0 1588 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1712622712
transform 1 0 1588 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1712622712
transform 1 0 1556 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1712622712
transform 1 0 1476 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1712622712
transform 1 0 1108 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1712622712
transform 1 0 964 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1712622712
transform 1 0 900 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1712622712
transform 1 0 868 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1712622712
transform 1 0 676 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1712622712
transform 1 0 556 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1712622712
transform 1 0 604 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1712622712
transform 1 0 556 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1712622712
transform 1 0 452 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1712622712
transform 1 0 420 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1712622712
transform 1 0 260 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1712622712
transform 1 0 212 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1712622712
transform 1 0 156 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1712622712
transform 1 0 228 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1712622712
transform 1 0 76 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1712622712
transform 1 0 204 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1712622712
transform 1 0 124 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1712622712
transform 1 0 1156 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1712622712
transform 1 0 1012 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1712622712
transform 1 0 1012 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1712622712
transform 1 0 932 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1712622712
transform 1 0 1388 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1712622712
transform 1 0 1348 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1712622712
transform 1 0 1564 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1712622712
transform 1 0 1516 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1712622712
transform 1 0 1940 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1712622712
transform 1 0 1860 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1712622712
transform 1 0 1820 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1712622712
transform 1 0 2028 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1712622712
transform 1 0 1996 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1712622712
transform 1 0 2708 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1712622712
transform 1 0 2532 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1712622712
transform 1 0 2724 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1712622712
transform 1 0 2700 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1712622712
transform 1 0 3188 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1712622712
transform 1 0 3108 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1712622712
transform 1 0 3100 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1712622712
transform 1 0 3036 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1712622712
transform 1 0 3404 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1712622712
transform 1 0 3316 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1712622712
transform 1 0 3284 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1712622712
transform 1 0 3228 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1712622712
transform 1 0 3132 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1712622712
transform 1 0 3124 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1712622712
transform 1 0 3036 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1712622712
transform 1 0 3244 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1712622712
transform 1 0 3092 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1712622712
transform 1 0 3292 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1712622712
transform 1 0 3260 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1712622712
transform 1 0 3164 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1712622712
transform 1 0 3204 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1712622712
transform 1 0 3172 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1712622712
transform 1 0 3420 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1712622712
transform 1 0 3380 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1712622712
transform 1 0 3316 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1712622712
transform 1 0 3260 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1712622712
transform 1 0 3236 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1712622712
transform 1 0 3220 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1712622712
transform 1 0 3116 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1712622712
transform 1 0 3060 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1712622712
transform 1 0 3412 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1712622712
transform 1 0 3404 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1712622712
transform 1 0 3364 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1712622712
transform 1 0 3364 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1712622712
transform 1 0 3364 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1712622712
transform 1 0 3180 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1712622712
transform 1 0 3396 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1712622712
transform 1 0 3396 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1712622712
transform 1 0 3364 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1712622712
transform 1 0 3364 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1712622712
transform 1 0 3316 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1712622712
transform 1 0 3236 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1712622712
transform 1 0 3228 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1712622712
transform 1 0 3204 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1712622712
transform 1 0 3140 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1712622712
transform 1 0 3140 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1712622712
transform 1 0 3268 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1712622712
transform 1 0 3244 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1712622712
transform 1 0 3236 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1712622712
transform 1 0 3204 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1712622712
transform 1 0 3204 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1712622712
transform 1 0 3172 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1712622712
transform 1 0 3124 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1712622712
transform 1 0 3076 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1712622712
transform 1 0 3196 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1712622712
transform 1 0 3188 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1712622712
transform 1 0 3172 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1712622712
transform 1 0 3092 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1712622712
transform 1 0 3092 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1712622712
transform 1 0 3084 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1712622712
transform 1 0 2644 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1712622712
transform 1 0 1716 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1712622712
transform 1 0 3364 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1712622712
transform 1 0 3300 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1712622712
transform 1 0 3172 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1712622712
transform 1 0 2132 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1712622712
transform 1 0 2092 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1712622712
transform 1 0 2124 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1712622712
transform 1 0 1972 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1712622712
transform 1 0 2140 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1712622712
transform 1 0 1980 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1712622712
transform 1 0 1900 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1712622712
transform 1 0 1900 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1712622712
transform 1 0 2276 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1712622712
transform 1 0 2132 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1712622712
transform 1 0 2220 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1712622712
transform 1 0 2220 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1712622712
transform 1 0 2220 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1712622712
transform 1 0 2188 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1712622712
transform 1 0 2188 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1712622712
transform 1 0 2156 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1712622712
transform 1 0 2532 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1712622712
transform 1 0 2428 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1712622712
transform 1 0 2380 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1712622712
transform 1 0 2500 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1712622712
transform 1 0 2460 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1712622712
transform 1 0 2380 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1712622712
transform 1 0 2340 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1712622712
transform 1 0 1660 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1712622712
transform 1 0 1636 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1712622712
transform 1 0 2668 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1712622712
transform 1 0 2628 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1712622712
transform 1 0 2580 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1712622712
transform 1 0 1420 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1712622712
transform 1 0 1348 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1712622712
transform 1 0 1316 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1712622712
transform 1 0 1300 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1712622712
transform 1 0 1244 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1712622712
transform 1 0 908 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1712622712
transform 1 0 1636 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1712622712
transform 1 0 1588 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1712622712
transform 1 0 1156 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1712622712
transform 1 0 1108 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1712622712
transform 1 0 1052 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1712622712
transform 1 0 996 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1712622712
transform 1 0 1116 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1712622712
transform 1 0 1092 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1712622712
transform 1 0 1476 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1712622712
transform 1 0 1444 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1712622712
transform 1 0 1212 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1712622712
transform 1 0 1172 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1712622712
transform 1 0 684 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1712622712
transform 1 0 604 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1712622712
transform 1 0 516 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1712622712
transform 1 0 1196 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1712622712
transform 1 0 1108 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1712622712
transform 1 0 804 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1712622712
transform 1 0 748 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1712622712
transform 1 0 804 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1712622712
transform 1 0 604 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1712622712
transform 1 0 892 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1712622712
transform 1 0 556 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1712622712
transform 1 0 236 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1712622712
transform 1 0 204 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1712622712
transform 1 0 316 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1712622712
transform 1 0 204 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1712622712
transform 1 0 732 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1712622712
transform 1 0 708 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1712622712
transform 1 0 444 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1712622712
transform 1 0 404 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1712622712
transform 1 0 252 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1712622712
transform 1 0 300 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1712622712
transform 1 0 276 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1712622712
transform 1 0 276 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1712622712
transform 1 0 172 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1712622712
transform 1 0 140 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1712622712
transform 1 0 420 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1712622712
transform 1 0 388 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1712622712
transform 1 0 132 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1712622712
transform 1 0 68 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1712622712
transform 1 0 116 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1712622712
transform 1 0 68 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1712622712
transform 1 0 252 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1712622712
transform 1 0 220 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1712622712
transform 1 0 212 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1712622712
transform 1 0 180 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1712622712
transform 1 0 180 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1712622712
transform 1 0 1868 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1712622712
transform 1 0 1692 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1712622712
transform 1 0 1652 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1712622712
transform 1 0 852 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1712622712
transform 1 0 820 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1712622712
transform 1 0 772 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1712622712
transform 1 0 708 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1712622712
transform 1 0 708 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1712622712
transform 1 0 684 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1712622712
transform 1 0 772 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1712622712
transform 1 0 732 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1712622712
transform 1 0 596 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1712622712
transform 1 0 564 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1712622712
transform 1 0 924 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1712622712
transform 1 0 900 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1712622712
transform 1 0 828 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1712622712
transform 1 0 788 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1712622712
transform 1 0 988 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1712622712
transform 1 0 500 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1712622712
transform 1 0 828 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1712622712
transform 1 0 804 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1712622712
transform 1 0 1244 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1712622712
transform 1 0 1188 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1712622712
transform 1 0 1404 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1712622712
transform 1 0 1132 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1712622712
transform 1 0 1508 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1712622712
transform 1 0 1380 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1712622712
transform 1 0 1700 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1712622712
transform 1 0 1580 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1712622712
transform 1 0 1340 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1712622712
transform 1 0 1028 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1712622712
transform 1 0 1556 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1712622712
transform 1 0 1268 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1712622712
transform 1 0 1268 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1712622712
transform 1 0 1156 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1712622712
transform 1 0 1068 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1712622712
transform 1 0 1004 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1712622712
transform 1 0 1588 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1712622712
transform 1 0 1260 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1712622712
transform 1 0 1540 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1712622712
transform 1 0 1500 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1712622712
transform 1 0 1796 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1712622712
transform 1 0 1628 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1712622712
transform 1 0 1948 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1712622712
transform 1 0 1884 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1712622712
transform 1 0 2164 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1712622712
transform 1 0 2124 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1712622712
transform 1 0 2172 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1712622712
transform 1 0 2044 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1712622712
transform 1 0 1852 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1712622712
transform 1 0 1820 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1712622712
transform 1 0 1884 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1712622712
transform 1 0 1836 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1712622712
transform 1 0 1772 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1712622712
transform 1 0 1684 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1712622712
transform 1 0 2028 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1712622712
transform 1 0 1828 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1712622712
transform 1 0 1748 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1712622712
transform 1 0 980 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1712622712
transform 1 0 948 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1712622712
transform 1 0 2604 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1712622712
transform 1 0 2404 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1712622712
transform 1 0 2140 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1712622712
transform 1 0 2076 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1712622712
transform 1 0 2060 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1712622712
transform 1 0 2060 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1712622712
transform 1 0 2852 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1712622712
transform 1 0 2516 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1712622712
transform 1 0 2460 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1712622712
transform 1 0 2460 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1712622712
transform 1 0 2268 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1712622712
transform 1 0 2180 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1712622712
transform 1 0 2020 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1712622712
transform 1 0 2844 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1712622712
transform 1 0 2636 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1712622712
transform 1 0 2292 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1712622712
transform 1 0 2564 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1712622712
transform 1 0 2468 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1712622712
transform 1 0 3412 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1712622712
transform 1 0 3340 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1712622712
transform 1 0 3300 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1712622712
transform 1 0 3412 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1712622712
transform 1 0 3356 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1712622712
transform 1 0 3316 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1712622712
transform 1 0 3252 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1712622712
transform 1 0 3340 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1712622712
transform 1 0 3316 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1712622712
transform 1 0 3292 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1712622712
transform 1 0 3252 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1712622712
transform 1 0 3404 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1712622712
transform 1 0 3356 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1712622712
transform 1 0 3324 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1712622712
transform 1 0 2948 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1712622712
transform 1 0 2900 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1712622712
transform 1 0 2692 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1712622712
transform 1 0 3356 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1712622712
transform 1 0 3268 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1712622712
transform 1 0 3252 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1712622712
transform 1 0 3188 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1712622712
transform 1 0 3132 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1712622712
transform 1 0 2852 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1712622712
transform 1 0 2332 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1712622712
transform 1 0 1452 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1712622712
transform 1 0 1284 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1712622712
transform 1 0 836 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1712622712
transform 1 0 3236 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1712622712
transform 1 0 3196 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1712622712
transform 1 0 3348 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1712622712
transform 1 0 3348 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1712622712
transform 1 0 3316 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1712622712
transform 1 0 2428 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1712622712
transform 1 0 2252 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1712622712
transform 1 0 2156 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1712622712
transform 1 0 2060 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1712622712
transform 1 0 1988 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1712622712
transform 1 0 1844 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1712622712
transform 1 0 1692 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1712622712
transform 1 0 1532 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1712622712
transform 1 0 1484 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1712622712
transform 1 0 1364 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1712622712
transform 1 0 1364 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1712622712
transform 1 0 1212 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1712622712
transform 1 0 1028 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1712622712
transform 1 0 3212 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1712622712
transform 1 0 3076 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1712622712
transform 1 0 3052 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1712622712
transform 1 0 3052 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1712622712
transform 1 0 3004 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1712622712
transform 1 0 3004 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1712622712
transform 1 0 1460 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1712622712
transform 1 0 1460 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1712622712
transform 1 0 1068 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1712622712
transform 1 0 1068 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1712622712
transform 1 0 964 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1712622712
transform 1 0 780 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1712622712
transform 1 0 780 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1712622712
transform 1 0 476 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1712622712
transform 1 0 436 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1712622712
transform 1 0 316 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1712622712
transform 1 0 276 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1712622712
transform 1 0 260 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1712622712
transform 1 0 212 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1712622712
transform 1 0 148 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1712622712
transform 1 0 92 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1712622712
transform 1 0 3412 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1712622712
transform 1 0 3412 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1712622712
transform 1 0 3348 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1712622712
transform 1 0 3340 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1712622712
transform 1 0 3340 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1712622712
transform 1 0 3324 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1712622712
transform 1 0 3220 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1712622712
transform 1 0 3204 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1712622712
transform 1 0 3196 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1712622712
transform 1 0 3196 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1712622712
transform 1 0 3172 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1712622712
transform 1 0 3108 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1712622712
transform 1 0 3060 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1712622712
transform 1 0 3052 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1712622712
transform 1 0 3044 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1712622712
transform 1 0 2980 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1712622712
transform 1 0 2932 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1712622712
transform 1 0 2812 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1712622712
transform 1 0 2812 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1712622712
transform 1 0 2788 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1712622712
transform 1 0 2756 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1712622712
transform 1 0 2740 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1712622712
transform 1 0 3348 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1712622712
transform 1 0 3340 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1712622712
transform 1 0 3308 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1712622712
transform 1 0 3308 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1712622712
transform 1 0 3244 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1712622712
transform 1 0 3236 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1712622712
transform 1 0 3172 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1712622712
transform 1 0 2956 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1712622712
transform 1 0 2956 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1712622712
transform 1 0 2892 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1712622712
transform 1 0 2892 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1712622712
transform 1 0 2764 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1712622712
transform 1 0 2652 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1712622712
transform 1 0 2564 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1712622712
transform 1 0 2532 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1712622712
transform 1 0 2532 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1712622712
transform 1 0 2468 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1712622712
transform 1 0 2356 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1712622712
transform 1 0 2220 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1712622712
transform 1 0 2156 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1712622712
transform 1 0 2156 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1712622712
transform 1 0 2036 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1712622712
transform 1 0 1916 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1712622712
transform 1 0 1804 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1712622712
transform 1 0 1692 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1712622712
transform 1 0 1580 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1712622712
transform 1 0 1428 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1712622712
transform 1 0 1332 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1712622712
transform 1 0 1220 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1712622712
transform 1 0 1004 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1712622712
transform 1 0 900 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1712622712
transform 1 0 3004 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1712622712
transform 1 0 2908 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1712622712
transform 1 0 2316 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1712622712
transform 1 0 1116 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1712622712
transform 1 0 1116 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1712622712
transform 1 0 796 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1712622712
transform 1 0 684 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1712622712
transform 1 0 580 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1712622712
transform 1 0 380 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1712622712
transform 1 0 364 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1712622712
transform 1 0 356 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1712622712
transform 1 0 316 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1712622712
transform 1 0 244 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1712622712
transform 1 0 204 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1712622712
transform 1 0 124 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1712622712
transform 1 0 2972 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1712622712
transform 1 0 2868 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1712622712
transform 1 0 2772 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1712622712
transform 1 0 2676 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1712622712
transform 1 0 2572 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1712622712
transform 1 0 2476 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1712622712
transform 1 0 2380 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1712622712
transform 1 0 2276 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1712622712
transform 1 0 2180 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1712622712
transform 1 0 2084 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1712622712
transform 1 0 1980 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1712622712
transform 1 0 1908 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1712622712
transform 1 0 1884 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1712622712
transform 1 0 1780 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1712622712
transform 1 0 1756 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1712622712
transform 1 0 1644 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1712622712
transform 1 0 1524 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1712622712
transform 1 0 1476 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1712622712
transform 1 0 1372 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1712622712
transform 1 0 1268 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1712622712
transform 1 0 1268 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1712622712
transform 1 0 1036 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1712622712
transform 1 0 1028 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1712622712
transform 1 0 980 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1712622712
transform 1 0 540 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1712622712
transform 1 0 204 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1712622712
transform 1 0 140 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1712622712
transform 1 0 92 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1712622712
transform 1 0 3428 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1712622712
transform 1 0 3420 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1712622712
transform 1 0 3348 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1712622712
transform 1 0 3340 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1712622712
transform 1 0 3236 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1712622712
transform 1 0 3124 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1712622712
transform 1 0 3116 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1712622712
transform 1 0 3092 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1712622712
transform 1 0 3092 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1712622712
transform 1 0 2956 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1712622712
transform 1 0 2748 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1712622712
transform 1 0 1756 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1712622712
transform 1 0 1756 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1712622712
transform 1 0 1164 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1712622712
transform 1 0 868 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1712622712
transform 1 0 756 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1712622712
transform 1 0 644 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1712622712
transform 1 0 428 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1712622712
transform 1 0 316 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1712622712
transform 1 0 2300 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1712622712
transform 1 0 2140 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1712622712
transform 1 0 1924 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1712622712
transform 1 0 1892 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1712622712
transform 1 0 1724 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1712622712
transform 1 0 2444 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1712622712
transform 1 0 2388 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1712622712
transform 1 0 2276 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1712622712
transform 1 0 2124 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1712622712
transform 1 0 2628 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1712622712
transform 1 0 2468 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1712622712
transform 1 0 2292 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1712622712
transform 1 0 2132 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1712622712
transform 1 0 1996 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1712622712
transform 1 0 1996 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1712622712
transform 1 0 1844 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1712622712
transform 1 0 1844 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1712622712
transform 1 0 1764 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1712622712
transform 1 0 1668 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1712622712
transform 1 0 1668 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1712622712
transform 1 0 1564 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1712622712
transform 1 0 1476 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1712622712
transform 1 0 1452 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1712622712
transform 1 0 2852 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1712622712
transform 1 0 2292 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1712622712
transform 1 0 1212 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1712622712
transform 1 0 1204 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1712622712
transform 1 0 916 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1712622712
transform 1 0 748 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1712622712
transform 1 0 188 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1712622712
transform 1 0 132 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1712622712
transform 1 0 100 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1712622712
transform 1 0 2836 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1712622712
transform 1 0 2428 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1712622712
transform 1 0 2428 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1712622712
transform 1 0 724 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1712622712
transform 1 0 724 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1712622712
transform 1 0 628 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1712622712
transform 1 0 508 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1712622712
transform 1 0 372 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1712622712
transform 1 0 308 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1712622712
transform 1 0 2756 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1712622712
transform 1 0 2412 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1712622712
transform 1 0 1116 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1712622712
transform 1 0 892 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1712622712
transform 1 0 2604 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1712622712
transform 1 0 2476 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1712622712
transform 1 0 2468 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1712622712
transform 1 0 2396 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1712622712
transform 1 0 2284 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1712622712
transform 1 0 2148 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1712622712
transform 1 0 1972 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1712622712
transform 1 0 2852 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1712622712
transform 1 0 2772 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1712622712
transform 1 0 2484 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1712622712
transform 1 0 2476 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1712622712
transform 1 0 1172 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1712622712
transform 1 0 900 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1712622712
transform 1 0 740 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1712622712
transform 1 0 644 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1712622712
transform 1 0 524 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1712622712
transform 1 0 436 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1712622712
transform 1 0 356 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1712622712
transform 1 0 324 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1712622712
transform 1 0 260 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1712622712
transform 1 0 180 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1712622712
transform 1 0 116 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1712622712
transform 1 0 3044 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1712622712
transform 1 0 2996 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1712622712
transform 1 0 2924 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1712622712
transform 1 0 3084 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1712622712
transform 1 0 2972 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1712622712
transform 1 0 2724 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1712622712
transform 1 0 2556 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1712622712
transform 1 0 2036 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1712622712
transform 1 0 1844 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1712622712
transform 1 0 1668 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1712622712
transform 1 0 1580 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1712622712
transform 1 0 1364 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1712622712
transform 1 0 1340 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1712622712
transform 1 0 1156 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1712622712
transform 1 0 1156 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1712622712
transform 1 0 948 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1712622712
transform 1 0 948 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1712622712
transform 1 0 364 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1712622712
transform 1 0 164 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1712622712
transform 1 0 140 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1712622712
transform 1 0 3020 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1712622712
transform 1 0 2932 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1712622712
transform 1 0 2932 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1712622712
transform 1 0 2828 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1712622712
transform 1 0 2492 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1712622712
transform 1 0 2524 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1712622712
transform 1 0 2308 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1712622712
transform 1 0 2236 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1712622712
transform 1 0 2148 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1712622712
transform 1 0 2028 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1712622712
transform 1 0 1956 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1712622712
transform 1 0 1956 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1712622712
transform 1 0 1828 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1712622712
transform 1 0 1828 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1712622712
transform 1 0 1732 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1712622712
transform 1 0 1652 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1712622712
transform 1 0 1484 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1712622712
transform 1 0 1372 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1712622712
transform 1 0 1276 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1712622712
transform 1 0 1212 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1712622712
transform 1 0 1156 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1712622712
transform 1 0 988 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1712622712
transform 1 0 988 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1712622712
transform 1 0 868 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1712622712
transform 1 0 868 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1712622712
transform 1 0 684 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1712622712
transform 1 0 676 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1712622712
transform 1 0 620 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1712622712
transform 1 0 572 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1712622712
transform 1 0 572 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1712622712
transform 1 0 548 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1712622712
transform 1 0 516 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1712622712
transform 1 0 516 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1712622712
transform 1 0 516 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1712622712
transform 1 0 484 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1712622712
transform 1 0 3036 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1712622712
transform 1 0 2884 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1712622712
transform 1 0 2788 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1712622712
transform 1 0 2748 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1712622712
transform 1 0 2716 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1712622712
transform 1 0 2708 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1712622712
transform 1 0 2532 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1712622712
transform 1 0 2396 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1712622712
transform 1 0 2316 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1712622712
transform 1 0 2180 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1712622712
transform 1 0 2180 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1712622712
transform 1 0 2092 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1712622712
transform 1 0 1988 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1712622712
transform 1 0 1932 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1712622712
transform 1 0 1788 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1712622712
transform 1 0 1620 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1712622712
transform 1 0 1572 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1712622712
transform 1 0 1396 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1712622712
transform 1 0 1388 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1712622712
transform 1 0 1300 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1712622712
transform 1 0 1148 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1712622712
transform 1 0 2372 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1712622712
transform 1 0 2276 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1712622712
transform 1 0 2196 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1712622712
transform 1 0 2196 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1712622712
transform 1 0 2140 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1712622712
transform 1 0 2140 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1712622712
transform 1 0 2132 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1712622712
transform 1 0 2132 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1712622712
transform 1 0 2124 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1712622712
transform 1 0 2116 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1712622712
transform 1 0 2084 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1712622712
transform 1 0 2044 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1712622712
transform 1 0 1940 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1712622712
transform 1 0 1940 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1712622712
transform 1 0 1860 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1712622712
transform 1 0 1780 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1712622712
transform 1 0 1772 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1712622712
transform 1 0 1772 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1712622712
transform 1 0 1756 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1712622712
transform 1 0 1732 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1712622712
transform 1 0 1732 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1712622712
transform 1 0 1716 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1712622712
transform 1 0 1684 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1712622712
transform 1 0 1484 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1712622712
transform 1 0 1484 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1712622712
transform 1 0 1012 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1712622712
transform 1 0 1012 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1712622712
transform 1 0 796 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1712622712
transform 1 0 788 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1712622712
transform 1 0 684 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1712622712
transform 1 0 644 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1712622712
transform 1 0 604 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1712622712
transform 1 0 508 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1712622712
transform 1 0 236 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1712622712
transform 1 0 236 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1712622712
transform 1 0 156 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1712622712
transform 1 0 156 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1712622712
transform 1 0 108 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1712622712
transform 1 0 108 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1712622712
transform 1 0 108 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1712622712
transform 1 0 92 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1712622712
transform 1 0 68 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1712622712
transform 1 0 68 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1712622712
transform 1 0 68 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1712622712
transform 1 0 2220 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1712622712
transform 1 0 1716 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1712622712
transform 1 0 1452 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1712622712
transform 1 0 1452 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1712622712
transform 1 0 572 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1712622712
transform 1 0 412 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1712622712
transform 1 0 404 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1712622712
transform 1 0 324 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1712622712
transform 1 0 308 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1712622712
transform 1 0 308 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1712622712
transform 1 0 308 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1712622712
transform 1 0 292 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1712622712
transform 1 0 292 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1712622712
transform 1 0 276 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1712622712
transform 1 0 276 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1712622712
transform 1 0 260 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1712622712
transform 1 0 252 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1712622712
transform 1 0 252 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1712622712
transform 1 0 252 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1712622712
transform 1 0 228 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1712622712
transform 1 0 228 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1712622712
transform 1 0 2412 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1712622712
transform 1 0 2396 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1712622712
transform 1 0 2396 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1712622712
transform 1 0 2396 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1712622712
transform 1 0 2364 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1712622712
transform 1 0 2364 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1712622712
transform 1 0 2356 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1712622712
transform 1 0 2268 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1712622712
transform 1 0 2204 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1712622712
transform 1 0 1940 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1712622712
transform 1 0 1844 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1712622712
transform 1 0 1772 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1712622712
transform 1 0 1588 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1712622712
transform 1 0 1484 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1712622712
transform 1 0 1116 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1712622712
transform 1 0 900 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1712622712
transform 1 0 2116 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1712622712
transform 1 0 2068 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1712622712
transform 1 0 2036 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1712622712
transform 1 0 2036 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1712622712
transform 1 0 1964 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1712622712
transform 1 0 1924 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1712622712
transform 1 0 1900 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1712622712
transform 1 0 1900 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1712622712
transform 1 0 1316 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1712622712
transform 1 0 1316 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1712622712
transform 1 0 724 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1712622712
transform 1 0 724 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1712622712
transform 1 0 604 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1712622712
transform 1 0 540 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1712622712
transform 1 0 300 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1712622712
transform 1 0 172 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1712622712
transform 1 0 172 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1712622712
transform 1 0 164 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1712622712
transform 1 0 164 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1712622712
transform 1 0 132 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1712622712
transform 1 0 132 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1712622712
transform 1 0 132 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1712622712
transform 1 0 68 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1712622712
transform 1 0 68 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1712622712
transform 1 0 2308 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1712622712
transform 1 0 2228 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1712622712
transform 1 0 2220 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1712622712
transform 1 0 2172 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1712622712
transform 1 0 2172 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1712622712
transform 1 0 2164 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1712622712
transform 1 0 2164 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1712622712
transform 1 0 2148 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1712622712
transform 1 0 2132 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1712622712
transform 1 0 2012 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1712622712
transform 1 0 2012 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1712622712
transform 1 0 1924 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1712622712
transform 1 0 1908 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1712622712
transform 1 0 1836 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1712622712
transform 1 0 1748 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1712622712
transform 1 0 1692 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1712622712
transform 1 0 1532 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1712622712
transform 1 0 1532 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1712622712
transform 1 0 1060 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1712622712
transform 1 0 868 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1712622712
transform 1 0 2740 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1712622712
transform 1 0 2708 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1712622712
transform 1 0 2972 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1712622712
transform 1 0 2956 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1712622712
transform 1 0 2852 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1712622712
transform 1 0 2636 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1712622712
transform 1 0 2556 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1712622712
transform 1 0 1764 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1712622712
transform 1 0 1404 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1712622712
transform 1 0 1156 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1712622712
transform 1 0 2564 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1712622712
transform 1 0 2492 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1712622712
transform 1 0 2492 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1712622712
transform 1 0 2484 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1712622712
transform 1 0 2476 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1712622712
transform 1 0 2476 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1712622712
transform 1 0 2476 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1712622712
transform 1 0 2436 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1712622712
transform 1 0 2436 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1712622712
transform 1 0 2348 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1712622712
transform 1 0 2332 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1712622712
transform 1 0 2332 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1712622712
transform 1 0 2044 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1712622712
transform 1 0 2044 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1712622712
transform 1 0 1948 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1712622712
transform 1 0 1844 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1712622712
transform 1 0 1732 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1712622712
transform 1 0 1556 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1712622712
transform 1 0 1516 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1712622712
transform 1 0 1516 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1712622712
transform 1 0 1484 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1712622712
transform 1 0 1476 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1712622712
transform 1 0 1476 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1712622712
transform 1 0 1164 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1712622712
transform 1 0 1164 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1712622712
transform 1 0 1036 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1712622712
transform 1 0 1036 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1712622712
transform 1 0 988 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1712622712
transform 1 0 948 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1712622712
transform 1 0 940 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1712622712
transform 1 0 836 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1712622712
transform 1 0 836 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1712622712
transform 1 0 804 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1712622712
transform 1 0 724 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1712622712
transform 1 0 724 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1712622712
transform 1 0 692 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1712622712
transform 1 0 604 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1712622712
transform 1 0 604 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1712622712
transform 1 0 596 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1712622712
transform 1 0 596 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1712622712
transform 1 0 596 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1712622712
transform 1 0 580 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1712622712
transform 1 0 580 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1712622712
transform 1 0 580 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1712622712
transform 1 0 580 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1712622712
transform 1 0 564 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1712622712
transform 1 0 548 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1712622712
transform 1 0 508 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1712622712
transform 1 0 500 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1712622712
transform 1 0 3164 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1712622712
transform 1 0 2844 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1712622712
transform 1 0 3140 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1712622712
transform 1 0 3132 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1712622712
transform 1 0 3092 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1712622712
transform 1 0 3060 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1712622712
transform 1 0 2892 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1712622712
transform 1 0 2588 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1712622712
transform 1 0 3228 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1712622712
transform 1 0 3140 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1712622712
transform 1 0 2836 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1712622712
transform 1 0 2804 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1712622712
transform 1 0 2540 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1712622712
transform 1 0 2492 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1712622712
transform 1 0 2476 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1712622712
transform 1 0 2468 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1712622712
transform 1 0 2468 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1712622712
transform 1 0 2452 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1712622712
transform 1 0 2452 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1712622712
transform 1 0 2444 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1712622712
transform 1 0 2444 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1712622712
transform 1 0 2444 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1712622712
transform 1 0 2444 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1712622712
transform 1 0 2436 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1712622712
transform 1 0 2316 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1712622712
transform 1 0 2308 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1712622712
transform 1 0 2300 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1712622712
transform 1 0 1916 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1712622712
transform 1 0 1812 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1712622712
transform 1 0 1812 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1712622712
transform 1 0 1772 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1712622712
transform 1 0 1772 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1712622712
transform 1 0 1724 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1712622712
transform 1 0 1724 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1712622712
transform 1 0 1700 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1712622712
transform 1 0 1452 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1712622712
transform 1 0 1108 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1712622712
transform 1 0 1108 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1712622712
transform 1 0 940 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1712622712
transform 1 0 764 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1712622712
transform 1 0 700 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1712622712
transform 1 0 660 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1712622712
transform 1 0 2828 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1712622712
transform 1 0 2740 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1712622712
transform 1 0 2596 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1712622712
transform 1 0 2596 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1712622712
transform 1 0 2012 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1712622712
transform 1 0 2012 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1712622712
transform 1 0 1460 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1712622712
transform 1 0 1428 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1712622712
transform 1 0 1316 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1712622712
transform 1 0 1316 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1712622712
transform 1 0 1300 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1712622712
transform 1 0 1236 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1712622712
transform 1 0 1220 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1712622712
transform 1 0 1220 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1712622712
transform 1 0 1100 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1712622712
transform 1 0 1100 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1712622712
transform 1 0 956 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1712622712
transform 1 0 948 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1712622712
transform 1 0 916 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1712622712
transform 1 0 916 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1712622712
transform 1 0 788 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1712622712
transform 1 0 788 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1712622712
transform 1 0 564 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1712622712
transform 1 0 516 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1712622712
transform 1 0 508 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1712622712
transform 1 0 452 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1712622712
transform 1 0 452 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1712622712
transform 1 0 2740 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1712622712
transform 1 0 2484 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1712622712
transform 1 0 3140 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1712622712
transform 1 0 3076 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1712622712
transform 1 0 2996 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1712622712
transform 1 0 2468 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1712622712
transform 1 0 2332 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1712622712
transform 1 0 2308 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1712622712
transform 1 0 2284 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1712622712
transform 1 0 2228 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1712622712
transform 1 0 2196 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1712622712
transform 1 0 2172 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1712622712
transform 1 0 2156 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1712622712
transform 1 0 2132 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1712622712
transform 1 0 2132 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1712622712
transform 1 0 1876 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1712622712
transform 1 0 1788 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1712622712
transform 1 0 1788 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1712622712
transform 1 0 1716 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1712622712
transform 1 0 1708 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1712622712
transform 1 0 1708 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1712622712
transform 1 0 1452 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1712622712
transform 1 0 1084 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1712622712
transform 1 0 1060 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1712622712
transform 1 0 836 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1712622712
transform 1 0 380 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1712622712
transform 1 0 324 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1712622712
transform 1 0 228 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1712622712
transform 1 0 2660 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1712622712
transform 1 0 2564 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1712622712
transform 1 0 2556 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1712622712
transform 1 0 2332 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1712622712
transform 1 0 2332 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1712622712
transform 1 0 2180 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1712622712
transform 1 0 2172 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1712622712
transform 1 0 2012 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1712622712
transform 1 0 2012 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1712622712
transform 1 0 1500 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1712622712
transform 1 0 1500 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1712622712
transform 1 0 1428 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1712622712
transform 1 0 1396 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1712622712
transform 1 0 1172 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1712622712
transform 1 0 1132 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1712622712
transform 1 0 852 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1712622712
transform 1 0 836 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1712622712
transform 1 0 628 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1712622712
transform 1 0 268 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1712622712
transform 1 0 268 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1712622712
transform 1 0 268 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1712622712
transform 1 0 260 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1712622712
transform 1 0 244 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1712622712
transform 1 0 236 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1712622712
transform 1 0 212 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1712622712
transform 1 0 212 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1712622712
transform 1 0 204 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1712622712
transform 1 0 204 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1712622712
transform 1 0 188 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1712622712
transform 1 0 188 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1712622712
transform 1 0 188 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1712622712
transform 1 0 2868 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1712622712
transform 1 0 2812 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1712622712
transform 1 0 2812 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1712622712
transform 1 0 2588 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1712622712
transform 1 0 1636 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1712622712
transform 1 0 1524 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1712622712
transform 1 0 1348 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1712622712
transform 1 0 2644 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1712622712
transform 1 0 2644 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1712622712
transform 1 0 2596 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1712622712
transform 1 0 2596 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1712622712
transform 1 0 2580 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1712622712
transform 1 0 2556 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1712622712
transform 1 0 2556 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1712622712
transform 1 0 2556 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1712622712
transform 1 0 2412 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1712622712
transform 1 0 2412 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1712622712
transform 1 0 2372 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1712622712
transform 1 0 2180 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1712622712
transform 1 0 2180 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1712622712
transform 1 0 2124 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1712622712
transform 1 0 2012 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1712622712
transform 1 0 1948 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1712622712
transform 1 0 1884 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1712622712
transform 1 0 1884 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1712622712
transform 1 0 1780 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1712622712
transform 1 0 1676 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1712622712
transform 1 0 1676 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1712622712
transform 1 0 1500 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1712622712
transform 1 0 1492 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1712622712
transform 1 0 1428 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1712622712
transform 1 0 1348 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1712622712
transform 1 0 1332 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1712622712
transform 1 0 1220 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1712622712
transform 1 0 948 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1712622712
transform 1 0 812 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1712622712
transform 1 0 756 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1712622712
transform 1 0 556 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1712622712
transform 1 0 540 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1712622712
transform 1 0 516 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1712622712
transform 1 0 516 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1712622712
transform 1 0 500 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1712622712
transform 1 0 492 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1712622712
transform 1 0 492 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1712622712
transform 1 0 484 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1712622712
transform 1 0 484 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1712622712
transform 1 0 476 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1712622712
transform 1 0 460 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1712622712
transform 1 0 460 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1712622712
transform 1 0 436 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1712622712
transform 1 0 412 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1712622712
transform 1 0 412 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1712622712
transform 1 0 404 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1712622712
transform 1 0 380 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1712622712
transform 1 0 380 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1712622712
transform 1 0 380 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1712622712
transform 1 0 3188 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1712622712
transform 1 0 3140 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1712622712
transform 1 0 3020 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1712622712
transform 1 0 3012 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1712622712
transform 1 0 3308 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1712622712
transform 1 0 3284 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1712622712
transform 1 0 3284 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1712622712
transform 1 0 3236 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1712622712
transform 1 0 3220 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1712622712
transform 1 0 2804 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1712622712
transform 1 0 3076 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1712622712
transform 1 0 3004 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1712622712
transform 1 0 2932 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1712622712
transform 1 0 2884 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1712622712
transform 1 0 2788 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1712622712
transform 1 0 2572 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1712622712
transform 1 0 2452 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1712622712
transform 1 0 2372 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1712622712
transform 1 0 2372 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1712622712
transform 1 0 2372 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1712622712
transform 1 0 2356 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1712622712
transform 1 0 2300 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1712622712
transform 1 0 2244 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1712622712
transform 1 0 2204 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1712622712
transform 1 0 2140 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1712622712
transform 1 0 2124 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1712622712
transform 1 0 2108 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1712622712
transform 1 0 2108 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1712622712
transform 1 0 1996 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1712622712
transform 1 0 1996 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1712622712
transform 1 0 1932 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1712622712
transform 1 0 1932 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1712622712
transform 1 0 1900 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1712622712
transform 1 0 1900 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1712622712
transform 1 0 1900 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1712622712
transform 1 0 1796 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1712622712
transform 1 0 1796 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1712622712
transform 1 0 1772 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1712622712
transform 1 0 1756 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1712622712
transform 1 0 1556 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1712622712
transform 1 0 1524 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1712622712
transform 1 0 1284 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1712622712
transform 1 0 1148 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1712622712
transform 1 0 1132 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1712622712
transform 1 0 1116 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1712622712
transform 1 0 1116 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1712622712
transform 1 0 860 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1712622712
transform 1 0 844 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1712622712
transform 1 0 844 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1712622712
transform 1 0 692 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1712622712
transform 1 0 612 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1712622712
transform 1 0 420 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1712622712
transform 1 0 420 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1712622712
transform 1 0 396 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1712622712
transform 1 0 324 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1712622712
transform 1 0 292 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1712622712
transform 1 0 292 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1712622712
transform 1 0 244 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1712622712
transform 1 0 244 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1712622712
transform 1 0 236 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1712622712
transform 1 0 228 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1712622712
transform 1 0 220 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1712622712
transform 1 0 220 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1712622712
transform 1 0 204 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1712622712
transform 1 0 188 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1712622712
transform 1 0 164 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1712622712
transform 1 0 148 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1712622712
transform 1 0 140 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1712622712
transform 1 0 140 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1712622712
transform 1 0 116 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1712622712
transform 1 0 116 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1712622712
transform 1 0 92 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1712622712
transform 1 0 92 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1712622712
transform 1 0 92 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1712622712
transform 1 0 2764 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1712622712
transform 1 0 2756 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1712622712
transform 1 0 2732 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1712622712
transform 1 0 2716 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1712622712
transform 1 0 2716 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1712622712
transform 1 0 2716 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1712622712
transform 1 0 2716 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1712622712
transform 1 0 2700 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1712622712
transform 1 0 2684 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1712622712
transform 1 0 2684 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1712622712
transform 1 0 2668 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1712622712
transform 1 0 2644 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1712622712
transform 1 0 2628 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1712622712
transform 1 0 2628 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1712622712
transform 1 0 2596 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1712622712
transform 1 0 2572 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1712622712
transform 1 0 2548 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1712622712
transform 1 0 2052 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1712622712
transform 1 0 2052 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1712622712
transform 1 0 2012 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1712622712
transform 1 0 2012 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1712622712
transform 1 0 1892 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1712622712
transform 1 0 1884 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1712622712
transform 1 0 1580 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1712622712
transform 1 0 1580 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1712622712
transform 1 0 1260 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1712622712
transform 1 0 1204 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1712622712
transform 1 0 1196 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1712622712
transform 1 0 1196 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1712622712
transform 1 0 1116 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1712622712
transform 1 0 1116 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1712622712
transform 1 0 2700 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1712622712
transform 1 0 2580 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1712622712
transform 1 0 2540 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1712622712
transform 1 0 2316 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1712622712
transform 1 0 2316 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1712622712
transform 1 0 2148 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1712622712
transform 1 0 2076 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1712622712
transform 1 0 2076 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1712622712
transform 1 0 2036 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1712622712
transform 1 0 2028 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1712622712
transform 1 0 2004 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1712622712
transform 1 0 2004 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1712622712
transform 1 0 1972 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1712622712
transform 1 0 1972 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1712622712
transform 1 0 1908 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1712622712
transform 1 0 1908 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1712622712
transform 1 0 1836 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1712622712
transform 1 0 1836 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1712622712
transform 1 0 1836 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1712622712
transform 1 0 1652 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1712622712
transform 1 0 1564 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1712622712
transform 1 0 1236 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1712622712
transform 1 0 1236 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1712622712
transform 1 0 1180 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1712622712
transform 1 0 1180 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1712622712
transform 1 0 1132 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1712622712
transform 1 0 1132 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1712622712
transform 1 0 1132 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1712622712
transform 1 0 1100 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1712622712
transform 1 0 1100 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1712622712
transform 1 0 1092 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1712622712
transform 1 0 1092 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1712622712
transform 1 0 1060 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1712622712
transform 1 0 1044 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1712622712
transform 1 0 3324 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1712622712
transform 1 0 3268 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1712622712
transform 1 0 3228 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1712622712
transform 1 0 3204 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1712622712
transform 1 0 1724 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1712622712
transform 1 0 1068 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1712622712
transform 1 0 932 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1712622712
transform 1 0 884 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1712622712
transform 1 0 692 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1712622712
transform 1 0 628 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1712622712
transform 1 0 508 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1712622712
transform 1 0 428 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1712622712
transform 1 0 356 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1712622712
transform 1 0 308 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1712622712
transform 1 0 260 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1712622712
transform 1 0 260 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1712622712
transform 1 0 188 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1712622712
transform 1 0 140 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1712622712
transform 1 0 84 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1712622712
transform 1 0 2868 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1712622712
transform 1 0 2676 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1712622712
transform 1 0 2332 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1712622712
transform 1 0 2268 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1712622712
transform 1 0 2236 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1712622712
transform 1 0 2084 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1712622712
transform 1 0 2044 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1712622712
transform 1 0 1884 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1712622712
transform 1 0 1828 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1712622712
transform 1 0 1772 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1712622712
transform 1 0 1764 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1712622712
transform 1 0 1668 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1712622712
transform 1 0 1444 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1712622712
transform 1 0 1372 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1712622712
transform 1 0 1292 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1712622712
transform 1 0 3340 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1712622712
transform 1 0 3332 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1712622712
transform 1 0 3332 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1712622712
transform 1 0 3332 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1712622712
transform 1 0 3284 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1712622712
transform 1 0 3244 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1712622712
transform 1 0 3244 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1712622712
transform 1 0 3220 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1712622712
transform 1 0 3220 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1712622712
transform 1 0 3172 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1712622712
transform 1 0 3124 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1712622712
transform 1 0 3108 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1712622712
transform 1 0 3108 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1712622712
transform 1 0 2996 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1712622712
transform 1 0 2956 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1712622712
transform 1 0 2804 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1712622712
transform 1 0 2780 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1712622712
transform 1 0 2684 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1712622712
transform 1 0 2604 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1712622712
transform 1 0 2452 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1712622712
transform 1 0 2452 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1712622712
transform 1 0 1340 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1712622712
transform 1 0 1780 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1712622712
transform 1 0 1468 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1712622712
transform 1 0 1468 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1712622712
transform 1 0 1252 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1712622712
transform 1 0 1244 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1712622712
transform 1 0 1180 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1712622712
transform 1 0 1100 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1712622712
transform 1 0 1092 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1712622712
transform 1 0 924 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1712622712
transform 1 0 636 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1712622712
transform 1 0 612 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1712622712
transform 1 0 588 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1712622712
transform 1 0 556 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1712622712
transform 1 0 524 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1712622712
transform 1 0 484 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1712622712
transform 1 0 436 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1712622712
transform 1 0 2484 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1712622712
transform 1 0 2444 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1712622712
transform 1 0 2252 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1712622712
transform 1 0 2188 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1712622712
transform 1 0 2116 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1712622712
transform 1 0 1988 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1712622712
transform 1 0 1924 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1712622712
transform 1 0 1668 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1712622712
transform 1 0 1668 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1712622712
transform 1 0 1620 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1712622712
transform 1 0 1444 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1712622712
transform 1 0 1324 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1712622712
transform 1 0 1324 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1712622712
transform 1 0 964 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1712622712
transform 1 0 3340 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1712622712
transform 1 0 3316 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1712622712
transform 1 0 3308 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1712622712
transform 1 0 3292 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1712622712
transform 1 0 3252 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1712622712
transform 1 0 3220 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1712622712
transform 1 0 3204 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1712622712
transform 1 0 3196 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1712622712
transform 1 0 3188 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1712622712
transform 1 0 3188 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1712622712
transform 1 0 3164 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1712622712
transform 1 0 3060 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1712622712
transform 1 0 3052 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1712622712
transform 1 0 3044 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1712622712
transform 1 0 2908 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1712622712
transform 1 0 2620 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1712622712
transform 1 0 2620 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1712622712
transform 1 0 2492 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1712622712
transform 1 0 2492 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1712622712
transform 1 0 1620 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1712622712
transform 1 0 1564 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1712622712
transform 1 0 1564 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1712622712
transform 1 0 1468 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1712622712
transform 1 0 1436 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1712622712
transform 1 0 1396 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1712622712
transform 1 0 2964 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1712622712
transform 1 0 2868 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1712622712
transform 1 0 2820 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1712622712
transform 1 0 2628 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1712622712
transform 1 0 2556 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1712622712
transform 1 0 2428 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1712622712
transform 1 0 2140 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1712622712
transform 1 0 1916 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1712622712
transform 1 0 1916 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1712622712
transform 1 0 1588 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1712622712
transform 1 0 1588 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1712622712
transform 1 0 1540 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1712622712
transform 1 0 1500 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1712622712
transform 1 0 1500 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1712622712
transform 1 0 1460 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1712622712
transform 1 0 1404 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1712622712
transform 1 0 1316 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1712622712
transform 1 0 1244 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1712622712
transform 1 0 1044 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1712622712
transform 1 0 956 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1712622712
transform 1 0 2652 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1712622712
transform 1 0 2572 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1712622712
transform 1 0 2412 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1712622712
transform 1 0 2372 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1712622712
transform 1 0 2364 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1712622712
transform 1 0 2308 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1712622712
transform 1 0 2308 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1712622712
transform 1 0 2196 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1712622712
transform 1 0 2188 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1712622712
transform 1 0 2044 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1712622712
transform 1 0 2044 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1712622712
transform 1 0 1836 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1712622712
transform 1 0 1796 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1712622712
transform 1 0 1756 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1712622712
transform 1 0 1756 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1712622712
transform 1 0 1748 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1712622712
transform 1 0 1628 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1712622712
transform 1 0 1412 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1712622712
transform 1 0 1276 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1712622712
transform 1 0 1140 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1712622712
transform 1 0 1140 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1712622712
transform 1 0 1060 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1712622712
transform 1 0 980 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1712622712
transform 1 0 892 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1712622712
transform 1 0 812 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1712622712
transform 1 0 812 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1712622712
transform 1 0 772 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1712622712
transform 1 0 772 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1712622712
transform 1 0 3108 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1712622712
transform 1 0 3100 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1712622712
transform 1 0 3084 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1712622712
transform 1 0 3084 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1712622712
transform 1 0 3036 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1712622712
transform 1 0 2428 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1712622712
transform 1 0 2172 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1712622712
transform 1 0 2140 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1712622712
transform 1 0 2140 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1712622712
transform 1 0 2124 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1712622712
transform 1 0 2124 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1712622712
transform 1 0 2068 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1712622712
transform 1 0 2068 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1712622712
transform 1 0 2012 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1712622712
transform 1 0 2012 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1712622712
transform 1 0 1980 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1712622712
transform 1 0 1940 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1712622712
transform 1 0 3052 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1712622712
transform 1 0 2988 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1712622712
transform 1 0 2988 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1712622712
transform 1 0 2948 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1712622712
transform 1 0 2820 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1712622712
transform 1 0 2820 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1712622712
transform 1 0 2780 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1712622712
transform 1 0 2764 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1712622712
transform 1 0 2724 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1712622712
transform 1 0 2108 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1712622712
transform 1 0 2100 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1712622712
transform 1 0 1908 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1712622712
transform 1 0 1836 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1712622712
transform 1 0 1836 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1712622712
transform 1 0 1836 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1712622712
transform 1 0 1748 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1712622712
transform 1 0 1748 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1712622712
transform 1 0 1716 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1712622712
transform 1 0 2436 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1712622712
transform 1 0 2388 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1712622712
transform 1 0 2340 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1712622712
transform 1 0 2292 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1712622712
transform 1 0 2292 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1712622712
transform 1 0 2276 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1712622712
transform 1 0 2276 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1712622712
transform 1 0 2276 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1712622712
transform 1 0 2252 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1712622712
transform 1 0 2252 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1712622712
transform 1 0 2244 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1712622712
transform 1 0 2156 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1712622712
transform 1 0 2132 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1712622712
transform 1 0 2188 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1712622712
transform 1 0 2180 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1712622712
transform 1 0 2156 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1712622712
transform 1 0 2108 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1712622712
transform 1 0 2108 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1712622712
transform 1 0 2076 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1712622712
transform 1 0 1876 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1712622712
transform 1 0 1868 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1712622712
transform 1 0 1860 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1712622712
transform 1 0 1796 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1712622712
transform 1 0 1620 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1712622712
transform 1 0 1612 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1712622712
transform 1 0 1604 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1712622712
transform 1 0 1604 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1712622712
transform 1 0 1572 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1712622712
transform 1 0 1572 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1712622712
transform 1 0 2380 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1712622712
transform 1 0 2284 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1712622712
transform 1 0 2284 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1712622712
transform 1 0 1724 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1712622712
transform 1 0 1644 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1712622712
transform 1 0 1636 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1712622712
transform 1 0 1524 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1712622712
transform 1 0 1524 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1712622712
transform 1 0 1388 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1712622712
transform 1 0 1340 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1712622712
transform 1 0 1020 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1712622712
transform 1 0 1020 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1712622712
transform 1 0 812 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1712622712
transform 1 0 732 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1712622712
transform 1 0 732 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1712622712
transform 1 0 668 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1712622712
transform 1 0 660 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1712622712
transform 1 0 660 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1712622712
transform 1 0 1260 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1712622712
transform 1 0 1148 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1712622712
transform 1 0 980 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1712622712
transform 1 0 956 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1712622712
transform 1 0 948 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1712622712
transform 1 0 892 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1712622712
transform 1 0 844 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1712622712
transform 1 0 788 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1712622712
transform 1 0 692 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1712622712
transform 1 0 692 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1712622712
transform 1 0 628 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1712622712
transform 1 0 596 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1712622712
transform 1 0 556 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1712622712
transform 1 0 340 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1712622712
transform 1 0 228 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1712622712
transform 1 0 180 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1712622712
transform 1 0 1628 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1712622712
transform 1 0 1404 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1712622712
transform 1 0 1404 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1712622712
transform 1 0 1252 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1712622712
transform 1 0 1236 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1712622712
transform 1 0 724 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1712622712
transform 1 0 724 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1712622712
transform 1 0 332 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1712622712
transform 1 0 316 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1712622712
transform 1 0 284 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1712622712
transform 1 0 252 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1712622712
transform 1 0 188 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1712622712
transform 1 0 900 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1712622712
transform 1 0 828 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1712622712
transform 1 0 788 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1712622712
transform 1 0 780 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1712622712
transform 1 0 620 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1712622712
transform 1 0 596 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1712622712
transform 1 0 596 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1712622712
transform 1 0 500 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1712622712
transform 1 0 444 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1712622712
transform 1 0 348 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1712622712
transform 1 0 292 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1712622712
transform 1 0 292 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1712622712
transform 1 0 108 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1712622712
transform 1 0 1228 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1712622712
transform 1 0 700 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1712622712
transform 1 0 700 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1712622712
transform 1 0 668 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1712622712
transform 1 0 652 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1712622712
transform 1 0 644 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1712622712
transform 1 0 484 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1712622712
transform 1 0 468 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1712622712
transform 1 0 412 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1712622712
transform 1 0 356 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1712622712
transform 1 0 332 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1712622712
transform 1 0 324 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1712622712
transform 1 0 308 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1712622712
transform 1 0 292 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1712622712
transform 1 0 276 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1712622712
transform 1 0 276 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1712622712
transform 1 0 1292 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1712622712
transform 1 0 1292 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1712622712
transform 1 0 1244 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1712622712
transform 1 0 1212 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1712622712
transform 1 0 1148 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1712622712
transform 1 0 1148 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1712622712
transform 1 0 1044 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1712622712
transform 1 0 1028 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1712622712
transform 1 0 1028 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1712622712
transform 1 0 980 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1712622712
transform 1 0 956 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1712622712
transform 1 0 948 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1712622712
transform 1 0 948 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1712622712
transform 1 0 892 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1712622712
transform 1 0 820 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1712622712
transform 1 0 764 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1712622712
transform 1 0 660 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1712622712
transform 1 0 628 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1712622712
transform 1 0 3436 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1712622712
transform 1 0 3436 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1712622712
transform 1 0 3436 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1712622712
transform 1 0 3420 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1712622712
transform 1 0 3380 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1712622712
transform 1 0 3380 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1712622712
transform 1 0 3372 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1712622712
transform 1 0 3276 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1712622712
transform 1 0 3276 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1712622712
transform 1 0 3276 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1712622712
transform 1 0 3260 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1712622712
transform 1 0 3260 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1712622712
transform 1 0 3260 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1712622712
transform 1 0 3244 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1712622712
transform 1 0 3236 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1712622712
transform 1 0 3172 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1712622712
transform 1 0 3036 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1712622712
transform 1 0 3396 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1712622712
transform 1 0 3204 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1712622712
transform 1 0 3148 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1712622712
transform 1 0 3140 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1712622712
transform 1 0 3076 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1712622712
transform 1 0 3356 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1712622712
transform 1 0 2916 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1712622712
transform 1 0 2700 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1712622712
transform 1 0 2692 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1712622712
transform 1 0 1748 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1712622712
transform 1 0 3284 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1712622712
transform 1 0 3140 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1712622712
transform 1 0 2692 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1712622712
transform 1 0 2676 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1712622712
transform 1 0 2660 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1712622712
transform 1 0 2628 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1712622712
transform 1 0 2620 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1712622712
transform 1 0 1684 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1712622712
transform 1 0 1620 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1712622712
transform 1 0 1620 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1712622712
transform 1 0 1572 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1712622712
transform 1 0 1444 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1712622712
transform 1 0 1444 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1712622712
transform 1 0 1068 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1712622712
transform 1 0 1404 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1712622712
transform 1 0 1348 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1712622712
transform 1 0 1260 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1712622712
transform 1 0 1188 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1712622712
transform 1 0 3004 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1712622712
transform 1 0 2980 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1712622712
transform 1 0 2980 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1712622712
transform 1 0 2916 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1712622712
transform 1 0 2852 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1712622712
transform 1 0 2844 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1712622712
transform 1 0 2828 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1712622712
transform 1 0 2716 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1712622712
transform 1 0 2348 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1712622712
transform 1 0 1604 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1712622712
transform 1 0 1604 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1712622712
transform 1 0 1580 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1712622712
transform 1 0 1460 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1712622712
transform 1 0 1332 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1712622712
transform 1 0 1332 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1712622712
transform 1 0 3276 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1712622712
transform 1 0 3212 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1712622712
transform 1 0 3212 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1712622712
transform 1 0 3172 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1712622712
transform 1 0 3236 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1712622712
transform 1 0 2796 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1712622712
transform 1 0 2292 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1712622712
transform 1 0 2292 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1712622712
transform 1 0 1620 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1712622712
transform 1 0 3332 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1712622712
transform 1 0 3228 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1712622712
transform 1 0 3180 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1712622712
transform 1 0 3196 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1712622712
transform 1 0 2372 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1712622712
transform 1 0 3396 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1712622712
transform 1 0 3324 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1712622712
transform 1 0 1444 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1712622712
transform 1 0 1316 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1712622712
transform 1 0 1316 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1712622712
transform 1 0 1276 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1712622712
transform 1 0 1188 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1712622712
transform 1 0 1148 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1712622712
transform 1 0 1428 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1712622712
transform 1 0 1308 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1712622712
transform 1 0 836 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1712622712
transform 1 0 700 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1712622712
transform 1 0 676 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1712622712
transform 1 0 1388 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1712622712
transform 1 0 1308 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1712622712
transform 1 0 1308 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1712622712
transform 1 0 1236 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1712622712
transform 1 0 1236 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1712622712
transform 1 0 1068 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1712622712
transform 1 0 1068 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1712622712
transform 1 0 964 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1712622712
transform 1 0 964 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1712622712
transform 1 0 836 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1712622712
transform 1 0 2260 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1712622712
transform 1 0 2044 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1712622712
transform 1 0 2036 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1712622712
transform 1 0 1964 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1712622712
transform 1 0 1948 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1712622712
transform 1 0 1604 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1712622712
transform 1 0 1564 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1712622712
transform 1 0 1564 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1712622712
transform 1 0 1444 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1712622712
transform 1 0 1340 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1712622712
transform 1 0 908 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1712622712
transform 1 0 740 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1712622712
transform 1 0 1084 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1712622712
transform 1 0 700 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1712622712
transform 1 0 540 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1712622712
transform 1 0 524 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1712622712
transform 1 0 476 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1712622712
transform 1 0 476 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1712622712
transform 1 0 476 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1712622712
transform 1 0 388 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1712622712
transform 1 0 388 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1712622712
transform 1 0 388 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1712622712
transform 1 0 236 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1712622712
transform 1 0 212 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1712622712
transform 1 0 212 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1712622712
transform 1 0 3084 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1712622712
transform 1 0 3044 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1712622712
transform 1 0 2908 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1712622712
transform 1 0 2900 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1712622712
transform 1 0 2740 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1712622712
transform 1 0 2740 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1712622712
transform 1 0 2684 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1712622712
transform 1 0 2532 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1712622712
transform 1 0 2532 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1712622712
transform 1 0 2172 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1712622712
transform 1 0 2084 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1712622712
transform 1 0 1108 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1712622712
transform 1 0 900 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1712622712
transform 1 0 900 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1712622712
transform 1 0 596 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1712622712
transform 1 0 548 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1712622712
transform 1 0 540 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1712622712
transform 1 0 316 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1712622712
transform 1 0 268 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1712622712
transform 1 0 268 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1712622712
transform 1 0 220 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1712622712
transform 1 0 212 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1712622712
transform 1 0 2652 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1712622712
transform 1 0 2564 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1712622712
transform 1 0 2540 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1712622712
transform 1 0 2500 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1712622712
transform 1 0 2492 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1712622712
transform 1 0 2476 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1712622712
transform 1 0 2476 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1712622712
transform 1 0 2460 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1712622712
transform 1 0 2460 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1712622712
transform 1 0 2348 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1712622712
transform 1 0 2348 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1712622712
transform 1 0 2340 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1712622712
transform 1 0 2316 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1712622712
transform 1 0 2148 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1712622712
transform 1 0 2148 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1712622712
transform 1 0 2060 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1712622712
transform 1 0 2060 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1712622712
transform 1 0 2052 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1712622712
transform 1 0 1868 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1712622712
transform 1 0 1852 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1712622712
transform 1 0 1844 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1712622712
transform 1 0 1828 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1712622712
transform 1 0 1828 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1712622712
transform 1 0 1748 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1712622712
transform 1 0 1748 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1712622712
transform 1 0 1636 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1712622712
transform 1 0 1596 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1712622712
transform 1 0 1580 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1712622712
transform 1 0 1580 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1712622712
transform 1 0 1580 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1712622712
transform 1 0 1524 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1712622712
transform 1 0 1524 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1712622712
transform 1 0 1444 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1712622712
transform 1 0 1436 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1712622712
transform 1 0 1420 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1712622712
transform 1 0 1420 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1712622712
transform 1 0 1356 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1712622712
transform 1 0 1348 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1712622712
transform 1 0 1292 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1712622712
transform 1 0 1164 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1712622712
transform 1 0 1164 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1712622712
transform 1 0 892 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1712622712
transform 1 0 724 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1712622712
transform 1 0 684 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1712622712
transform 1 0 516 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1712622712
transform 1 0 500 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1712622712
transform 1 0 500 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1712622712
transform 1 0 500 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1712622712
transform 1 0 500 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1712622712
transform 1 0 484 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1712622712
transform 1 0 484 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1712622712
transform 1 0 468 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1712622712
transform 1 0 436 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1712622712
transform 1 0 436 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1712622712
transform 1 0 428 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1712622712
transform 1 0 420 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1712622712
transform 1 0 412 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1712622712
transform 1 0 380 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1712622712
transform 1 0 372 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1712622712
transform 1 0 2716 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1712622712
transform 1 0 2676 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1712622712
transform 1 0 2580 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1712622712
transform 1 0 2204 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1712622712
transform 1 0 2204 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1712622712
transform 1 0 2188 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1712622712
transform 1 0 3420 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1712622712
transform 1 0 3364 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1712622712
transform 1 0 3364 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1712622712
transform 1 0 3260 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1712622712
transform 1 0 3188 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1712622712
transform 1 0 3076 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1712622712
transform 1 0 3068 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1712622712
transform 1 0 2972 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1712622712
transform 1 0 3340 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1712622712
transform 1 0 3284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1712622712
transform 1 0 3436 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1712622712
transform 1 0 3388 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1712622712
transform 1 0 3412 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1712622712
transform 1 0 3412 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1712622712
transform 1 0 3388 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1712622712
transform 1 0 3356 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1712622712
transform 1 0 3348 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1712622712
transform 1 0 3324 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1712622712
transform 1 0 2980 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1712622712
transform 1 0 2908 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1712622712
transform 1 0 2812 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1712622712
transform 1 0 2748 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1712622712
transform 1 0 3356 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1712622712
transform 1 0 3300 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1712622712
transform 1 0 2732 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1712622712
transform 1 0 2652 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1712622712
transform 1 0 2548 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1712622712
transform 1 0 3220 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1712622712
transform 1 0 2748 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1712622712
transform 1 0 2628 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1712622712
transform 1 0 3220 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1712622712
transform 1 0 3124 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1712622712
transform 1 0 2700 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1712622712
transform 1 0 2660 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1712622712
transform 1 0 2620 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1712622712
transform 1 0 2612 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1712622712
transform 1 0 2924 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1712622712
transform 1 0 2724 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1712622712
transform 1 0 2724 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1712622712
transform 1 0 2668 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1712622712
transform 1 0 2780 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1712622712
transform 1 0 2772 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1712622712
transform 1 0 2716 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1712622712
transform 1 0 2692 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1712622712
transform 1 0 2692 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1712622712
transform 1 0 3260 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1712622712
transform 1 0 3132 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1712622712
transform 1 0 3220 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1712622712
transform 1 0 3164 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1712622712
transform 1 0 3396 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1712622712
transform 1 0 3300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1712622712
transform 1 0 3260 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1712622712
transform 1 0 3172 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1712622712
transform 1 0 2860 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1712622712
transform 1 0 2820 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1712622712
transform 1 0 2260 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1712622712
transform 1 0 2228 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1712622712
transform 1 0 2068 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1712622712
transform 1 0 2028 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1712622712
transform 1 0 1876 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1712622712
transform 1 0 1828 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1712622712
transform 1 0 1812 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1712622712
transform 1 0 1692 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1712622712
transform 1 0 1684 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1712622712
transform 1 0 1580 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1712622712
transform 1 0 292 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1712622712
transform 1 0 244 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1712622712
transform 1 0 340 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1712622712
transform 1 0 244 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1712622712
transform 1 0 412 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1712622712
transform 1 0 364 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1712622712
transform 1 0 1364 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1712622712
transform 1 0 1212 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1712622712
transform 1 0 2092 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1712622712
transform 1 0 1732 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1712622712
transform 1 0 3420 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1712622712
transform 1 0 3380 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1712622712
transform 1 0 3228 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1712622712
transform 1 0 3044 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1712622712
transform 1 0 2924 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1712622712
transform 1 0 2868 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1712622712
transform 1 0 3244 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1712622712
transform 1 0 3212 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1712622712
transform 1 0 2772 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1712622712
transform 1 0 2724 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1712622712
transform 1 0 2612 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1712622712
transform 1 0 3364 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2584
timestamp 1712622712
transform 1 0 3340 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1712622712
transform 1 0 3404 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1712622712
transform 1 0 3308 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1712622712
transform 1 0 2940 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1712622712
transform 1 0 1756 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1712622712
transform 1 0 1756 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1712622712
transform 1 0 1756 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1712622712
transform 1 0 1700 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1712622712
transform 1 0 1700 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1712622712
transform 1 0 1660 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1712622712
transform 1 0 1660 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1712622712
transform 1 0 1724 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1712622712
transform 1 0 1668 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1712622712
transform 1 0 1740 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1712622712
transform 1 0 1580 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2599
timestamp 1712622712
transform 1 0 1556 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1712622712
transform 1 0 1532 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1712622712
transform 1 0 1524 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1712622712
transform 1 0 1468 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1712622712
transform 1 0 1500 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1712622712
transform 1 0 1484 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1712622712
transform 1 0 1532 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1712622712
transform 1 0 1476 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1712622712
transform 1 0 1492 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1712622712
transform 1 0 1484 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1712622712
transform 1 0 1476 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1712622712
transform 1 0 1452 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1712622712
transform 1 0 1452 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1712622712
transform 1 0 1452 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1712622712
transform 1 0 2068 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1712622712
transform 1 0 1452 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1712622712
transform 1 0 1460 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1712622712
transform 1 0 980 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1712622712
transform 1 0 924 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1712622712
transform 1 0 284 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1712622712
transform 1 0 1100 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1712622712
transform 1 0 964 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1712622712
transform 1 0 972 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1712622712
transform 1 0 684 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1712622712
transform 1 0 1004 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1712622712
transform 1 0 964 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1712622712
transform 1 0 1684 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1712622712
transform 1 0 996 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1712622712
transform 1 0 780 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1712622712
transform 1 0 1068 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1712622712
transform 1 0 1020 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1712622712
transform 1 0 1540 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1712622712
transform 1 0 1436 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1712622712
transform 1 0 1436 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1712622712
transform 1 0 1372 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1712622712
transform 1 0 1060 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1712622712
transform 1 0 1244 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1712622712
transform 1 0 1172 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1712622712
transform 1 0 1084 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1712622712
transform 1 0 652 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1712622712
transform 1 0 548 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1712622712
transform 1 0 548 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1712622712
transform 1 0 388 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1712622712
transform 1 0 692 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1712622712
transform 1 0 644 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1712622712
transform 1 0 1148 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1712622712
transform 1 0 1084 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1712622712
transform 1 0 1044 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1712622712
transform 1 0 900 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1712622712
transform 1 0 836 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1712622712
transform 1 0 1364 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1712622712
transform 1 0 1172 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1712622712
transform 1 0 1164 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1712622712
transform 1 0 1132 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1712622712
transform 1 0 236 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1712622712
transform 1 0 212 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1712622712
transform 1 0 268 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1712622712
transform 1 0 196 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1712622712
transform 1 0 220 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1712622712
transform 1 0 172 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1712622712
transform 1 0 308 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1712622712
transform 1 0 252 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1712622712
transform 1 0 204 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1712622712
transform 1 0 532 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1712622712
transform 1 0 308 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1712622712
transform 1 0 308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1712622712
transform 1 0 260 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1712622712
transform 1 0 260 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1712622712
transform 1 0 252 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1712622712
transform 1 0 316 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1712622712
transform 1 0 276 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1712622712
transform 1 0 212 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1712622712
transform 1 0 508 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1712622712
transform 1 0 172 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1712622712
transform 1 0 2212 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1712622712
transform 1 0 2132 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1712622712
transform 1 0 2252 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1712622712
transform 1 0 2212 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1712622712
transform 1 0 2204 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1712622712
transform 1 0 1788 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1712622712
transform 1 0 2308 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1712622712
transform 1 0 2292 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1712622712
transform 1 0 2324 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1712622712
transform 1 0 2212 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1712622712
transform 1 0 2372 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1712622712
transform 1 0 2132 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1712622712
transform 1 0 2100 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1712622712
transform 1 0 1956 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1712622712
transform 1 0 1444 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1712622712
transform 1 0 1076 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1712622712
transform 1 0 1036 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1712622712
transform 1 0 964 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1712622712
transform 1 0 1052 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1712622712
transform 1 0 956 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1712622712
transform 1 0 972 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1712622712
transform 1 0 876 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1712622712
transform 1 0 428 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1712622712
transform 1 0 332 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1712622712
transform 1 0 1572 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1712622712
transform 1 0 1492 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1712622712
transform 1 0 2244 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1712622712
transform 1 0 1516 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1712622712
transform 1 0 2428 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1712622712
transform 1 0 2308 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1712622712
transform 1 0 2308 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1712622712
transform 1 0 2204 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1712622712
transform 1 0 2252 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1712622712
transform 1 0 2148 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1712622712
transform 1 0 1700 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1712622712
transform 1 0 1596 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1712622712
transform 1 0 1580 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1712622712
transform 1 0 1444 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1712622712
transform 1 0 1444 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1712622712
transform 1 0 1284 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1712622712
transform 1 0 1908 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1712622712
transform 1 0 1700 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1712622712
transform 1 0 1692 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1712622712
transform 1 0 1508 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1712622712
transform 1 0 1692 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2718
timestamp 1712622712
transform 1 0 1524 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1712622712
transform 1 0 1524 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1712622712
transform 1 0 396 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1712622712
transform 1 0 532 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1712622712
transform 1 0 532 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1712622712
transform 1 0 476 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1712622712
transform 1 0 396 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1712622712
transform 1 0 444 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1712622712
transform 1 0 420 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1712622712
transform 1 0 780 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1712622712
transform 1 0 412 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1712622712
transform 1 0 868 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1712622712
transform 1 0 804 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1712622712
transform 1 0 924 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1712622712
transform 1 0 812 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1712622712
transform 1 0 892 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1712622712
transform 1 0 748 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1712622712
transform 1 0 2988 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1712622712
transform 1 0 2940 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1712622712
transform 1 0 2940 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1712622712
transform 1 0 2868 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1712622712
transform 1 0 2588 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1712622712
transform 1 0 2508 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1712622712
transform 1 0 2508 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1712622712
transform 1 0 2500 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2743
timestamp 1712622712
transform 1 0 1652 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1712622712
transform 1 0 1644 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1712622712
transform 1 0 1620 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1712622712
transform 1 0 2652 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1712622712
transform 1 0 2604 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1712622712
transform 1 0 1748 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1712622712
transform 1 0 1748 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1712622712
transform 1 0 1652 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1712622712
transform 1 0 492 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1712622712
transform 1 0 444 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1712622712
transform 1 0 420 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1712622712
transform 1 0 436 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1712622712
transform 1 0 380 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1712622712
transform 1 0 484 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2757
timestamp 1712622712
transform 1 0 412 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1712622712
transform 1 0 980 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1712622712
transform 1 0 412 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1712622712
transform 1 0 500 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1712622712
transform 1 0 420 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1712622712
transform 1 0 1188 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2763
timestamp 1712622712
transform 1 0 1004 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1712622712
transform 1 0 956 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1712622712
transform 1 0 988 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1712622712
transform 1 0 948 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2767
timestamp 1712622712
transform 1 0 884 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1712622712
transform 1 0 540 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1712622712
transform 1 0 476 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1712622712
transform 1 0 492 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1712622712
transform 1 0 460 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1712622712
transform 1 0 388 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1712622712
transform 1 0 1772 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1712622712
transform 1 0 1684 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1712622712
transform 1 0 1772 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1712622712
transform 1 0 1740 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1712622712
transform 1 0 1628 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1712622712
transform 1 0 1652 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1712622712
transform 1 0 1572 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1712622712
transform 1 0 1524 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1712622712
transform 1 0 1124 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1712622712
transform 1 0 1116 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1712622712
transform 1 0 956 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1712622712
transform 1 0 812 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1712622712
transform 1 0 812 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1712622712
transform 1 0 796 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1712622712
transform 1 0 796 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1712622712
transform 1 0 660 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1712622712
transform 1 0 1532 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1712622712
transform 1 0 1308 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1712622712
transform 1 0 1588 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1712622712
transform 1 0 1492 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1712622712
transform 1 0 940 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1712622712
transform 1 0 628 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1712622712
transform 1 0 196 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1712622712
transform 1 0 196 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1712622712
transform 1 0 196 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1712622712
transform 1 0 148 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1712622712
transform 1 0 140 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1712622712
transform 1 0 140 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1712622712
transform 1 0 92 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1712622712
transform 1 0 1764 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1712622712
transform 1 0 1740 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1712622712
transform 1 0 2244 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1712622712
transform 1 0 1836 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1712622712
transform 1 0 2492 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2807
timestamp 1712622712
transform 1 0 2372 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1712622712
transform 1 0 2268 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1712622712
transform 1 0 2188 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1712622712
transform 1 0 2364 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1712622712
transform 1 0 2236 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1712622712
transform 1 0 2500 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1712622712
transform 1 0 2276 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1712622712
transform 1 0 2236 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1712622712
transform 1 0 2260 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2816
timestamp 1712622712
transform 1 0 2180 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1712622712
transform 1 0 2444 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1712622712
transform 1 0 2284 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1712622712
transform 1 0 2284 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1712622712
transform 1 0 2228 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1712622712
transform 1 0 1868 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1712622712
transform 1 0 1804 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1712622712
transform 1 0 1724 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1712622712
transform 1 0 1940 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1712622712
transform 1 0 1732 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1712622712
transform 1 0 1652 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2827
timestamp 1712622712
transform 1 0 1388 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2828
timestamp 1712622712
transform 1 0 2588 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1712622712
transform 1 0 1900 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1712622712
transform 1 0 1844 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1712622712
transform 1 0 1292 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1712622712
transform 1 0 1268 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1712622712
transform 1 0 2204 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1712622712
transform 1 0 2156 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1712622712
transform 1 0 1868 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2836
timestamp 1712622712
transform 1 0 1844 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1712622712
transform 1 0 1828 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1712622712
transform 1 0 1796 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1712622712
transform 1 0 1748 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2840
timestamp 1712622712
transform 1 0 1540 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1712622712
transform 1 0 2116 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1712622712
transform 1 0 1932 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1712622712
transform 1 0 1948 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1712622712
transform 1 0 1876 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1712622712
transform 1 0 1764 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2846
timestamp 1712622712
transform 1 0 2628 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1712622712
transform 1 0 2596 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1712622712
transform 1 0 2764 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1712622712
transform 1 0 2764 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1712622712
transform 1 0 2660 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1712622712
transform 1 0 2572 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1712622712
transform 1 0 2588 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1712622712
transform 1 0 2524 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1712622712
transform 1 0 2492 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1712622712
transform 1 0 2652 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1712622712
transform 1 0 2452 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1712622712
transform 1 0 1628 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1712622712
transform 1 0 1404 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1712622712
transform 1 0 1412 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1712622712
transform 1 0 884 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1712622712
transform 1 0 836 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1712622712
transform 1 0 588 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1712622712
transform 1 0 964 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1712622712
transform 1 0 964 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1712622712
transform 1 0 884 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1712622712
transform 1 0 868 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1712622712
transform 1 0 844 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1712622712
transform 1 0 652 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1712622712
transform 1 0 1668 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1712622712
transform 1 0 892 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2871
timestamp 1712622712
transform 1 0 1660 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1712622712
transform 1 0 1068 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2873
timestamp 1712622712
transform 1 0 1140 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1712622712
transform 1 0 1044 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1712622712
transform 1 0 1044 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2876
timestamp 1712622712
transform 1 0 924 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1712622712
transform 1 0 1204 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1712622712
transform 1 0 1084 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1712622712
transform 1 0 988 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1712622712
transform 1 0 2596 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1712622712
transform 1 0 2596 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1712622712
transform 1 0 2572 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1712622712
transform 1 0 1684 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1712622712
transform 1 0 596 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1712622712
transform 1 0 508 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1712622712
transform 1 0 652 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1712622712
transform 1 0 540 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1712622712
transform 1 0 644 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1712622712
transform 1 0 516 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1712622712
transform 1 0 620 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1712622712
transform 1 0 556 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1712622712
transform 1 0 668 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1712622712
transform 1 0 572 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1712622712
transform 1 0 524 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1712622712
transform 1 0 492 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1712622712
transform 1 0 724 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1712622712
transform 1 0 652 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1712622712
transform 1 0 556 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1712622712
transform 1 0 1044 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1712622712
transform 1 0 852 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1712622712
transform 1 0 852 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1712622712
transform 1 0 756 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1712622712
transform 1 0 756 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1712622712
transform 1 0 684 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1712622712
transform 1 0 996 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1712622712
transform 1 0 964 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1712622712
transform 1 0 2100 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1712622712
transform 1 0 2084 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1712622712
transform 1 0 2052 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1712622712
transform 1 0 2044 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1712622712
transform 1 0 1828 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1712622712
transform 1 0 1316 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1712622712
transform 1 0 1292 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1712622712
transform 1 0 1228 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1712622712
transform 1 0 1172 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1712622712
transform 1 0 652 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1712622712
transform 1 0 516 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1712622712
transform 1 0 668 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1712622712
transform 1 0 564 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1712622712
transform 1 0 2308 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1712622712
transform 1 0 1636 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1712622712
transform 1 0 1756 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1712622712
transform 1 0 1644 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1712622712
transform 1 0 2308 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1712622712
transform 1 0 1780 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1712622712
transform 1 0 1836 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1712622712
transform 1 0 1804 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1712622712
transform 1 0 1884 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1712622712
transform 1 0 1860 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1712622712
transform 1 0 1892 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1712622712
transform 1 0 1788 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1712622712
transform 1 0 2292 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1712622712
transform 1 0 2292 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1712622712
transform 1 0 2244 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1712622712
transform 1 0 2244 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1712622712
transform 1 0 2220 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1712622712
transform 1 0 2212 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1712622712
transform 1 0 2204 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1712622712
transform 1 0 2204 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1712622712
transform 1 0 2140 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1712622712
transform 1 0 2076 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1712622712
transform 1 0 2028 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1712622712
transform 1 0 2004 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1712622712
transform 1 0 1580 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1712622712
transform 1 0 1556 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1712622712
transform 1 0 1460 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1712622712
transform 1 0 2404 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1712622712
transform 1 0 2332 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1712622712
transform 1 0 2388 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1712622712
transform 1 0 2348 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1712622712
transform 1 0 2436 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1712622712
transform 1 0 2372 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1712622712
transform 1 0 2100 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1712622712
transform 1 0 2404 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1712622712
transform 1 0 2188 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2956
timestamp 1712622712
transform 1 0 2420 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1712622712
transform 1 0 2348 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1712622712
transform 1 0 2220 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1712622712
transform 1 0 2420 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1712622712
transform 1 0 2316 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2961
timestamp 1712622712
transform 1 0 2156 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1712622712
transform 1 0 2396 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2963
timestamp 1712622712
transform 1 0 2276 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1712622712
transform 1 0 2284 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1712622712
transform 1 0 2260 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1712622712
transform 1 0 2244 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1712622712
transform 1 0 2204 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1712622712
transform 1 0 2020 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1712622712
transform 1 0 2420 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1712622712
transform 1 0 2420 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1712622712
transform 1 0 2348 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1712622712
transform 1 0 2348 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2973
timestamp 1712622712
transform 1 0 2308 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1712622712
transform 1 0 2292 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1712622712
transform 1 0 2516 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1712622712
transform 1 0 2436 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1712622712
transform 1 0 2380 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1712622712
transform 1 0 1556 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1712622712
transform 1 0 1236 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1712622712
transform 1 0 1772 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1712622712
transform 1 0 1772 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1712622712
transform 1 0 1748 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1712622712
transform 1 0 1708 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1712622712
transform 1 0 1572 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1712622712
transform 1 0 1612 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1712622712
transform 1 0 1476 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1712622712
transform 1 0 1340 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1712622712
transform 1 0 1228 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1712622712
transform 1 0 1140 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1712622712
transform 1 0 1260 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1712622712
transform 1 0 1228 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1712622712
transform 1 0 1188 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1712622712
transform 1 0 1428 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1712622712
transform 1 0 1380 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2995
timestamp 1712622712
transform 1 0 1364 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2996
timestamp 1712622712
transform 1 0 1300 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2997
timestamp 1712622712
transform 1 0 1300 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1712622712
transform 1 0 468 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1712622712
transform 1 0 444 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1712622712
transform 1 0 196 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1712622712
transform 1 0 196 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1712622712
transform 1 0 100 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1712622712
transform 1 0 2052 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1712622712
transform 1 0 1940 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1712622712
transform 1 0 1940 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1712622712
transform 1 0 1532 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1712622712
transform 1 0 1540 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1712622712
transform 1 0 820 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3009
timestamp 1712622712
transform 1 0 732 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1712622712
transform 1 0 532 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1712622712
transform 1 0 932 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1712622712
transform 1 0 820 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3013
timestamp 1712622712
transform 1 0 1348 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1712622712
transform 1 0 1292 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1712622712
transform 1 0 1284 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1712622712
transform 1 0 996 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1712622712
transform 1 0 940 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1712622712
transform 1 0 940 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3019
timestamp 1712622712
transform 1 0 916 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1712622712
transform 1 0 884 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1712622712
transform 1 0 332 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1712622712
transform 1 0 332 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1712622712
transform 1 0 308 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3024
timestamp 1712622712
transform 1 0 1036 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1712622712
transform 1 0 940 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1712622712
transform 1 0 916 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1712622712
transform 1 0 916 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1712622712
transform 1 0 836 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1712622712
transform 1 0 996 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1712622712
transform 1 0 956 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3031
timestamp 1712622712
transform 1 0 932 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1712622712
transform 1 0 940 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1712622712
transform 1 0 788 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1712622712
transform 1 0 804 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1712622712
transform 1 0 732 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1712622712
transform 1 0 1052 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1712622712
transform 1 0 980 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1712622712
transform 1 0 916 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1712622712
transform 1 0 916 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3040
timestamp 1712622712
transform 1 0 684 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1712622712
transform 1 0 588 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1712622712
transform 1 0 756 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1712622712
transform 1 0 740 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1712622712
transform 1 0 692 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1712622712
transform 1 0 684 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1712622712
transform 1 0 1076 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1712622712
transform 1 0 892 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1712622712
transform 1 0 1388 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3049
timestamp 1712622712
transform 1 0 1212 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1712622712
transform 1 0 1140 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3051
timestamp 1712622712
transform 1 0 1140 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1712622712
transform 1 0 1020 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1712622712
transform 1 0 956 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1712622712
transform 1 0 812 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1712622712
transform 1 0 732 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1712622712
transform 1 0 684 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1712622712
transform 1 0 620 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1712622712
transform 1 0 860 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1712622712
transform 1 0 804 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1712622712
transform 1 0 756 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1712622712
transform 1 0 756 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1712622712
transform 1 0 636 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1712622712
transform 1 0 580 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1712622712
transform 1 0 988 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1712622712
transform 1 0 892 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1712622712
transform 1 0 788 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1712622712
transform 1 0 684 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1712622712
transform 1 0 636 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1712622712
transform 1 0 636 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1712622712
transform 1 0 2484 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1712622712
transform 1 0 2444 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1712622712
transform 1 0 2188 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1712622712
transform 1 0 2188 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1712622712
transform 1 0 1484 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1712622712
transform 1 0 1140 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1712622712
transform 1 0 1092 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1712622712
transform 1 0 1044 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1712622712
transform 1 0 996 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1712622712
transform 1 0 812 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1712622712
transform 1 0 612 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1712622712
transform 1 0 1004 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1712622712
transform 1 0 852 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1712622712
transform 1 0 668 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1712622712
transform 1 0 588 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1712622712
transform 1 0 588 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1712622712
transform 1 0 500 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1712622712
transform 1 0 572 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1712622712
transform 1 0 508 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1712622712
transform 1 0 812 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1712622712
transform 1 0 724 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1712622712
transform 1 0 724 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1712622712
transform 1 0 580 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1712622712
transform 1 0 548 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1712622712
transform 1 0 796 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1712622712
transform 1 0 708 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1712622712
transform 1 0 668 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1712622712
transform 1 0 644 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1712622712
transform 1 0 588 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1712622712
transform 1 0 588 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1712622712
transform 1 0 2060 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1712622712
transform 1 0 2036 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1712622712
transform 1 0 2532 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1712622712
transform 1 0 2028 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1712622712
transform 1 0 2036 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1712622712
transform 1 0 1444 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1712622712
transform 1 0 2316 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1712622712
transform 1 0 2292 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1712622712
transform 1 0 2260 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1712622712
transform 1 0 2196 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1712622712
transform 1 0 1812 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1712622712
transform 1 0 1724 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1712622712
transform 1 0 1724 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1712622712
transform 1 0 1668 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1712622712
transform 1 0 1588 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1712622712
transform 1 0 1412 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1712622712
transform 1 0 1460 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1712622712
transform 1 0 1412 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1712622712
transform 1 0 1492 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1712622712
transform 1 0 1484 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1712622712
transform 1 0 1404 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1712622712
transform 1 0 1404 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1712622712
transform 1 0 1364 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1712622712
transform 1 0 1340 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1712622712
transform 1 0 1236 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1712622712
transform 1 0 1476 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1712622712
transform 1 0 1420 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1712622712
transform 1 0 1420 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1712622712
transform 1 0 1172 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1712622712
transform 1 0 2060 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1712622712
transform 1 0 1988 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1712622712
transform 1 0 2252 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1712622712
transform 1 0 2092 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1712622712
transform 1 0 2516 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1712622712
transform 1 0 2196 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1712622712
transform 1 0 2196 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1712622712
transform 1 0 2012 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1712622712
transform 1 0 1612 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1712622712
transform 1 0 1612 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1712622712
transform 1 0 1564 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3140
timestamp 1712622712
transform 1 0 2252 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1712622712
transform 1 0 1892 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1712622712
transform 1 0 1820 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1712622712
transform 1 0 1940 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1712622712
transform 1 0 1924 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1712622712
transform 1 0 1916 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1712622712
transform 1 0 1876 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1712622712
transform 1 0 1852 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1712622712
transform 1 0 2004 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1712622712
transform 1 0 1820 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1712622712
transform 1 0 1820 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1712622712
transform 1 0 1724 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1712622712
transform 1 0 1724 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1712622712
transform 1 0 1628 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1712622712
transform 1 0 2612 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1712622712
transform 1 0 2516 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1712622712
transform 1 0 2460 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1712622712
transform 1 0 2436 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1712622712
transform 1 0 2428 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1712622712
transform 1 0 2428 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1712622712
transform 1 0 2388 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1712622712
transform 1 0 2388 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1712622712
transform 1 0 2348 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1712622712
transform 1 0 2340 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1712622712
transform 1 0 2652 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1712622712
transform 1 0 2548 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3166
timestamp 1712622712
transform 1 0 2548 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1712622712
transform 1 0 2524 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1712622712
transform 1 0 2524 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1712622712
transform 1 0 2516 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1712622712
transform 1 0 2476 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1712622712
transform 1 0 2132 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1712622712
transform 1 0 2100 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3173
timestamp 1712622712
transform 1 0 3108 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1712622712
transform 1 0 3108 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1712622712
transform 1 0 3028 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1712622712
transform 1 0 2972 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1712622712
transform 1 0 2908 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1712622712
transform 1 0 2548 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1712622712
transform 1 0 2548 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3180
timestamp 1712622712
transform 1 0 2500 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1712622712
transform 1 0 2276 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1712622712
transform 1 0 2260 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1712622712
transform 1 0 2260 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1712622712
transform 1 0 2244 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1712622712
transform 1 0 2156 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3186
timestamp 1712622712
transform 1 0 2140 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1712622712
transform 1 0 2052 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1712622712
transform 1 0 2028 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1712622712
transform 1 0 2060 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1712622712
transform 1 0 2028 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1712622712
transform 1 0 2020 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1712622712
transform 1 0 2004 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1712622712
transform 1 0 1908 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3194
timestamp 1712622712
transform 1 0 1868 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1712622712
transform 1 0 1788 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1712622712
transform 1 0 1732 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3197
timestamp 1712622712
transform 1 0 2260 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1712622712
transform 1 0 2132 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1712622712
transform 1 0 2124 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1712622712
transform 1 0 2116 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1712622712
transform 1 0 2108 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1712622712
transform 1 0 2084 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1712622712
transform 1 0 2076 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1712622712
transform 1 0 1988 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1712622712
transform 1 0 1668 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3206
timestamp 1712622712
transform 1 0 1628 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1712622712
transform 1 0 3300 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1712622712
transform 1 0 1940 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1712622712
transform 1 0 1628 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1712622712
transform 1 0 1564 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1712622712
transform 1 0 1348 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1712622712
transform 1 0 1548 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1712622712
transform 1 0 1532 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1712622712
transform 1 0 1884 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1712622712
transform 1 0 1620 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1712622712
transform 1 0 1612 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1712622712
transform 1 0 1524 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1712622712
transform 1 0 1508 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3219
timestamp 1712622712
transform 1 0 372 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3220
timestamp 1712622712
transform 1 0 1572 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3221
timestamp 1712622712
transform 1 0 1524 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1712622712
transform 1 0 1540 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3223
timestamp 1712622712
transform 1 0 1524 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1712622712
transform 1 0 1540 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1712622712
transform 1 0 804 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1712622712
transform 1 0 764 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1712622712
transform 1 0 724 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3228
timestamp 1712622712
transform 1 0 572 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1712622712
transform 1 0 516 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1712622712
transform 1 0 524 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1712622712
transform 1 0 476 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1712622712
transform 1 0 524 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1712622712
transform 1 0 380 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3234
timestamp 1712622712
transform 1 0 1524 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3235
timestamp 1712622712
transform 1 0 1332 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1712622712
transform 1 0 1300 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1712622712
transform 1 0 2068 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3238
timestamp 1712622712
transform 1 0 2044 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1712622712
transform 1 0 1900 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3240
timestamp 1712622712
transform 1 0 1884 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3241
timestamp 1712622712
transform 1 0 1812 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1712622712
transform 1 0 1812 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1712622712
transform 1 0 1580 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3244
timestamp 1712622712
transform 1 0 356 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1712622712
transform 1 0 340 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1712622712
transform 1 0 388 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3247
timestamp 1712622712
transform 1 0 356 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3248
timestamp 1712622712
transform 1 0 428 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1712622712
transform 1 0 356 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1712622712
transform 1 0 388 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1712622712
transform 1 0 372 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1712622712
transform 1 0 428 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1712622712
transform 1 0 340 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1712622712
transform 1 0 412 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1712622712
transform 1 0 332 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1712622712
transform 1 0 476 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1712622712
transform 1 0 412 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1712622712
transform 1 0 412 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1712622712
transform 1 0 364 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1712622712
transform 1 0 452 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1712622712
transform 1 0 420 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1712622712
transform 1 0 340 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1712622712
transform 1 0 372 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1712622712
transform 1 0 332 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3265
timestamp 1712622712
transform 1 0 1916 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1712622712
transform 1 0 1852 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1712622712
transform 1 0 2756 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1712622712
transform 1 0 2756 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1712622712
transform 1 0 2724 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1712622712
transform 1 0 1868 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1712622712
transform 1 0 2828 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1712622712
transform 1 0 2796 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1712622712
transform 1 0 2788 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1712622712
transform 1 0 2692 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1712622712
transform 1 0 2716 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1712622712
transform 1 0 2652 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1712622712
transform 1 0 2612 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1712622712
transform 1 0 2540 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1712622712
transform 1 0 2236 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1712622712
transform 1 0 2668 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1712622712
transform 1 0 2468 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1712622712
transform 1 0 2332 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1712622712
transform 1 0 2724 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1712622712
transform 1 0 2548 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1712622712
transform 1 0 2548 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1712622712
transform 1 0 2492 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1712622712
transform 1 0 1900 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1712622712
transform 1 0 1876 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1712622712
transform 1 0 2196 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3290
timestamp 1712622712
transform 1 0 1956 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1712622712
transform 1 0 2412 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3292
timestamp 1712622712
transform 1 0 2316 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1712622712
transform 1 0 2180 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1712622712
transform 1 0 2212 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1712622712
transform 1 0 2156 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1712622712
transform 1 0 1988 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1712622712
transform 1 0 1924 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1712622712
transform 1 0 1860 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1712622712
transform 1 0 1908 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1712622712
transform 1 0 1836 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1712622712
transform 1 0 1748 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3302
timestamp 1712622712
transform 1 0 1996 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1712622712
transform 1 0 1540 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1712622712
transform 1 0 1556 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3305
timestamp 1712622712
transform 1 0 1284 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3306
timestamp 1712622712
transform 1 0 1260 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1712622712
transform 1 0 1220 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1712622712
transform 1 0 1372 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3309
timestamp 1712622712
transform 1 0 1284 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1712622712
transform 1 0 1268 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1712622712
transform 1 0 1268 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1712622712
transform 1 0 1196 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3313
timestamp 1712622712
transform 1 0 1244 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3314
timestamp 1712622712
transform 1 0 1172 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3315
timestamp 1712622712
transform 1 0 1124 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3316
timestamp 1712622712
transform 1 0 932 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1712622712
transform 1 0 2460 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3318
timestamp 1712622712
transform 1 0 2036 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1712622712
transform 1 0 2476 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3320
timestamp 1712622712
transform 1 0 2180 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3321
timestamp 1712622712
transform 1 0 2092 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3322
timestamp 1712622712
transform 1 0 1852 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3323
timestamp 1712622712
transform 1 0 1660 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3324
timestamp 1712622712
transform 1 0 1332 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1712622712
transform 1 0 1332 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1712622712
transform 1 0 1300 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3327
timestamp 1712622712
transform 1 0 188 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1712622712
transform 1 0 1308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1712622712
transform 1 0 1124 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3330
timestamp 1712622712
transform 1 0 1124 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3331
timestamp 1712622712
transform 1 0 1004 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3332
timestamp 1712622712
transform 1 0 1004 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3333
timestamp 1712622712
transform 1 0 908 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3334
timestamp 1712622712
transform 1 0 908 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1712622712
transform 1 0 772 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3336
timestamp 1712622712
transform 1 0 772 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3337
timestamp 1712622712
transform 1 0 660 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3338
timestamp 1712622712
transform 1 0 1684 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3339
timestamp 1712622712
transform 1 0 1324 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1712622712
transform 1 0 2012 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3341
timestamp 1712622712
transform 1 0 1708 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1712622712
transform 1 0 2164 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3343
timestamp 1712622712
transform 1 0 1700 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1712622712
transform 1 0 1684 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3345
timestamp 1712622712
transform 1 0 1652 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3346
timestamp 1712622712
transform 1 0 1708 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1712622712
transform 1 0 1636 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1712622712
transform 1 0 1604 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1712622712
transform 1 0 1620 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1712622712
transform 1 0 1516 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3351
timestamp 1712622712
transform 1 0 1412 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3352
timestamp 1712622712
transform 1 0 1212 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1712622712
transform 1 0 1084 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3354
timestamp 1712622712
transform 1 0 1084 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3355
timestamp 1712622712
transform 1 0 1052 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1712622712
transform 1 0 2212 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1712622712
transform 1 0 2188 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1712622712
transform 1 0 2220 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1712622712
transform 1 0 2188 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3360
timestamp 1712622712
transform 1 0 2244 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1712622712
transform 1 0 2188 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1712622712
transform 1 0 2052 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3363
timestamp 1712622712
transform 1 0 1988 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1712622712
transform 1 0 2220 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1712622712
transform 1 0 1988 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3366
timestamp 1712622712
transform 1 0 2124 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1712622712
transform 1 0 1980 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3368
timestamp 1712622712
transform 1 0 2108 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3369
timestamp 1712622712
transform 1 0 2076 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1712622712
transform 1 0 2060 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3371
timestamp 1712622712
transform 1 0 2012 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1712622712
transform 1 0 1956 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1712622712
transform 1 0 1988 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1712622712
transform 1 0 1852 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3375
timestamp 1712622712
transform 1 0 2396 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1712622712
transform 1 0 2204 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3377
timestamp 1712622712
transform 1 0 2180 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3378
timestamp 1712622712
transform 1 0 2068 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3379
timestamp 1712622712
transform 1 0 2332 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3380
timestamp 1712622712
transform 1 0 2236 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3381
timestamp 1712622712
transform 1 0 2172 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3382
timestamp 1712622712
transform 1 0 2124 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3383
timestamp 1712622712
transform 1 0 2028 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3384
timestamp 1712622712
transform 1 0 2052 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3385
timestamp 1712622712
transform 1 0 1908 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3386
timestamp 1712622712
transform 1 0 1868 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3387
timestamp 1712622712
transform 1 0 636 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1712622712
transform 1 0 300 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3389
timestamp 1712622712
transform 1 0 260 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1712622712
transform 1 0 108 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3391
timestamp 1712622712
transform 1 0 268 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1712622712
transform 1 0 220 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1712622712
transform 1 0 820 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3394
timestamp 1712622712
transform 1 0 788 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3395
timestamp 1712622712
transform 1 0 684 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3396
timestamp 1712622712
transform 1 0 700 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3397
timestamp 1712622712
transform 1 0 556 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3398
timestamp 1712622712
transform 1 0 460 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3399
timestamp 1712622712
transform 1 0 172 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3400
timestamp 1712622712
transform 1 0 300 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3401
timestamp 1712622712
transform 1 0 172 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3402
timestamp 1712622712
transform 1 0 1236 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1712622712
transform 1 0 212 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3404
timestamp 1712622712
transform 1 0 204 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3405
timestamp 1712622712
transform 1 0 124 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3406
timestamp 1712622712
transform 1 0 596 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3407
timestamp 1712622712
transform 1 0 492 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3408
timestamp 1712622712
transform 1 0 340 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3409
timestamp 1712622712
transform 1 0 172 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3410
timestamp 1712622712
transform 1 0 148 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3411
timestamp 1712622712
transform 1 0 1796 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3412
timestamp 1712622712
transform 1 0 1620 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3413
timestamp 1712622712
transform 1 0 1604 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1712622712
transform 1 0 1452 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3415
timestamp 1712622712
transform 1 0 3204 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3416
timestamp 1712622712
transform 1 0 1692 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1712622712
transform 1 0 1684 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3418
timestamp 1712622712
transform 1 0 1636 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3419
timestamp 1712622712
transform 1 0 1588 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3420
timestamp 1712622712
transform 1 0 1508 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3421
timestamp 1712622712
transform 1 0 1420 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1712622712
transform 1 0 1420 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1712622712
transform 1 0 1396 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3424
timestamp 1712622712
transform 1 0 1396 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3425
timestamp 1712622712
transform 1 0 1380 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3426
timestamp 1712622712
transform 1 0 1380 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3427
timestamp 1712622712
transform 1 0 900 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3428
timestamp 1712622712
transform 1 0 1428 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3429
timestamp 1712622712
transform 1 0 380 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1712622712
transform 1 0 356 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3431
timestamp 1712622712
transform 1 0 300 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3432
timestamp 1712622712
transform 1 0 372 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3433
timestamp 1712622712
transform 1 0 356 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1712622712
transform 1 0 1012 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3435
timestamp 1712622712
transform 1 0 492 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1712622712
transform 1 0 492 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3437
timestamp 1712622712
transform 1 0 252 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3438
timestamp 1712622712
transform 1 0 396 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1712622712
transform 1 0 340 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1712622712
transform 1 0 332 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3441
timestamp 1712622712
transform 1 0 292 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1712622712
transform 1 0 412 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3443
timestamp 1712622712
transform 1 0 356 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1712622712
transform 1 0 356 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3445
timestamp 1712622712
transform 1 0 268 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3446
timestamp 1712622712
transform 1 0 1644 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1712622712
transform 1 0 1500 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3448
timestamp 1712622712
transform 1 0 1500 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1712622712
transform 1 0 1324 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3450
timestamp 1712622712
transform 1 0 892 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3451
timestamp 1712622712
transform 1 0 548 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1712622712
transform 1 0 1972 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3453
timestamp 1712622712
transform 1 0 1732 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1712622712
transform 1 0 1732 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1712622712
transform 1 0 1660 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1712622712
transform 1 0 1660 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3457
timestamp 1712622712
transform 1 0 540 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3458
timestamp 1712622712
transform 1 0 324 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1712622712
transform 1 0 292 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1712622712
transform 1 0 348 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1712622712
transform 1 0 292 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3462
timestamp 1712622712
transform 1 0 324 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1712622712
transform 1 0 292 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1712622712
transform 1 0 356 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3465
timestamp 1712622712
transform 1 0 252 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1712622712
transform 1 0 2172 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1712622712
transform 1 0 2092 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1712622712
transform 1 0 2084 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3469
timestamp 1712622712
transform 1 0 668 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1712622712
transform 1 0 2140 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3471
timestamp 1712622712
transform 1 0 2028 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3472
timestamp 1712622712
transform 1 0 1956 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1712622712
transform 1 0 1940 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3474
timestamp 1712622712
transform 1 0 1612 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1712622712
transform 1 0 1612 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3476
timestamp 1712622712
transform 1 0 868 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3477
timestamp 1712622712
transform 1 0 828 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1712622712
transform 1 0 772 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3479
timestamp 1712622712
transform 1 0 380 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3480
timestamp 1712622712
transform 1 0 308 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3481
timestamp 1712622712
transform 1 0 284 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3482
timestamp 1712622712
transform 1 0 372 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3483
timestamp 1712622712
transform 1 0 308 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1712622712
transform 1 0 308 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3485
timestamp 1712622712
transform 1 0 228 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1712622712
transform 1 0 2148 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3487
timestamp 1712622712
transform 1 0 564 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3488
timestamp 1712622712
transform 1 0 988 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3489
timestamp 1712622712
transform 1 0 828 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1712622712
transform 1 0 580 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3491
timestamp 1712622712
transform 1 0 540 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3492
timestamp 1712622712
transform 1 0 452 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3493
timestamp 1712622712
transform 1 0 460 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3494
timestamp 1712622712
transform 1 0 300 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3495
timestamp 1712622712
transform 1 0 276 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3496
timestamp 1712622712
transform 1 0 988 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3497
timestamp 1712622712
transform 1 0 972 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3498
timestamp 1712622712
transform 1 0 956 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1712622712
transform 1 0 956 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1712622712
transform 1 0 820 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3501
timestamp 1712622712
transform 1 0 492 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3502
timestamp 1712622712
transform 1 0 708 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3503
timestamp 1712622712
transform 1 0 708 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3504
timestamp 1712622712
transform 1 0 628 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3505
timestamp 1712622712
transform 1 0 620 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3506
timestamp 1712622712
transform 1 0 612 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3507
timestamp 1712622712
transform 1 0 612 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3508
timestamp 1712622712
transform 1 0 580 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1712622712
transform 1 0 580 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3510
timestamp 1712622712
transform 1 0 572 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3511
timestamp 1712622712
transform 1 0 516 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3512
timestamp 1712622712
transform 1 0 516 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1712622712
transform 1 0 492 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1712622712
transform 1 0 724 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3515
timestamp 1712622712
transform 1 0 724 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3516
timestamp 1712622712
transform 1 0 700 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1712622712
transform 1 0 676 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3518
timestamp 1712622712
transform 1 0 676 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3519
timestamp 1712622712
transform 1 0 564 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3520
timestamp 1712622712
transform 1 0 564 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3521
timestamp 1712622712
transform 1 0 548 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3522
timestamp 1712622712
transform 1 0 500 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3523
timestamp 1712622712
transform 1 0 1940 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3524
timestamp 1712622712
transform 1 0 1724 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3525
timestamp 1712622712
transform 1 0 1508 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1712622712
transform 1 0 1508 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3527
timestamp 1712622712
transform 1 0 1468 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3528
timestamp 1712622712
transform 1 0 1508 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1712622712
transform 1 0 1468 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3530
timestamp 1712622712
transform 1 0 1420 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1712622712
transform 1 0 1372 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3532
timestamp 1712622712
transform 1 0 1028 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3533
timestamp 1712622712
transform 1 0 844 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3534
timestamp 1712622712
transform 1 0 836 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3535
timestamp 1712622712
transform 1 0 620 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3536
timestamp 1712622712
transform 1 0 612 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3537
timestamp 1712622712
transform 1 0 412 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3538
timestamp 1712622712
transform 1 0 412 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3539
timestamp 1712622712
transform 1 0 140 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3540
timestamp 1712622712
transform 1 0 1628 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3541
timestamp 1712622712
transform 1 0 1468 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1712622712
transform 1 0 1516 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3543
timestamp 1712622712
transform 1 0 1452 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3544
timestamp 1712622712
transform 1 0 1380 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1712622712
transform 1 0 2404 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1712622712
transform 1 0 1804 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3547
timestamp 1712622712
transform 1 0 1868 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3548
timestamp 1712622712
transform 1 0 1868 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3549
timestamp 1712622712
transform 1 0 1852 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3550
timestamp 1712622712
transform 1 0 1820 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3551
timestamp 1712622712
transform 1 0 1940 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3552
timestamp 1712622712
transform 1 0 1812 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1712622712
transform 1 0 1844 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3554
timestamp 1712622712
transform 1 0 1348 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3555
timestamp 1712622712
transform 1 0 1484 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3556
timestamp 1712622712
transform 1 0 1428 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1712622712
transform 1 0 1260 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3558
timestamp 1712622712
transform 1 0 1332 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3559
timestamp 1712622712
transform 1 0 1164 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3560
timestamp 1712622712
transform 1 0 1836 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1712622712
transform 1 0 1820 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1712622712
transform 1 0 1724 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3563
timestamp 1712622712
transform 1 0 1724 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3564
timestamp 1712622712
transform 1 0 1716 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3565
timestamp 1712622712
transform 1 0 1668 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3566
timestamp 1712622712
transform 1 0 1660 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1712622712
transform 1 0 1572 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1712622712
transform 1 0 1308 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3569
timestamp 1712622712
transform 1 0 1180 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1712622712
transform 1 0 996 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1712622712
transform 1 0 2380 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3572
timestamp 1712622712
transform 1 0 1964 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3573
timestamp 1712622712
transform 1 0 2476 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3574
timestamp 1712622712
transform 1 0 2348 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3575
timestamp 1712622712
transform 1 0 2388 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3576
timestamp 1712622712
transform 1 0 2308 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3577
timestamp 1712622712
transform 1 0 2956 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1712622712
transform 1 0 2940 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3579
timestamp 1712622712
transform 1 0 2476 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3580
timestamp 1712622712
transform 1 0 2412 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3581
timestamp 1712622712
transform 1 0 2324 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3582
timestamp 1712622712
transform 1 0 2284 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3583
timestamp 1712622712
transform 1 0 1932 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3584
timestamp 1712622712
transform 1 0 2628 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3585
timestamp 1712622712
transform 1 0 2620 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3586
timestamp 1712622712
transform 1 0 2564 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3587
timestamp 1712622712
transform 1 0 2548 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3588
timestamp 1712622712
transform 1 0 2548 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3589
timestamp 1712622712
transform 1 0 2532 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1712622712
transform 1 0 2404 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3591
timestamp 1712622712
transform 1 0 1836 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3592
timestamp 1712622712
transform 1 0 1764 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3593
timestamp 1712622712
transform 1 0 2244 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1712622712
transform 1 0 2084 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3595
timestamp 1712622712
transform 1 0 2084 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3596
timestamp 1712622712
transform 1 0 1764 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3597
timestamp 1712622712
transform 1 0 1828 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3598
timestamp 1712622712
transform 1 0 1772 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3599
timestamp 1712622712
transform 1 0 1860 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1712622712
transform 1 0 1820 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1712622712
transform 1 0 2044 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3602
timestamp 1712622712
transform 1 0 1940 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3603
timestamp 1712622712
transform 1 0 1876 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3604
timestamp 1712622712
transform 1 0 1868 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3605
timestamp 1712622712
transform 1 0 2908 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3606
timestamp 1712622712
transform 1 0 2852 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3607
timestamp 1712622712
transform 1 0 2636 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1712622712
transform 1 0 2628 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1712622712
transform 1 0 2596 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1712622712
transform 1 0 2556 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3611
timestamp 1712622712
transform 1 0 2436 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1712622712
transform 1 0 2044 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1712622712
transform 1 0 2036 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1712622712
transform 1 0 2004 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3615
timestamp 1712622712
transform 1 0 1908 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1712622712
transform 1 0 3044 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3617
timestamp 1712622712
transform 1 0 2900 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1712622712
transform 1 0 2484 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1712622712
transform 1 0 2740 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1712622712
transform 1 0 2076 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1712622712
transform 1 0 2076 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3622
timestamp 1712622712
transform 1 0 1876 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1712622712
transform 1 0 2276 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1712622712
transform 1 0 2236 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3625
timestamp 1712622712
transform 1 0 2468 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1712622712
transform 1 0 2356 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3627
timestamp 1712622712
transform 1 0 2356 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3628
timestamp 1712622712
transform 1 0 2340 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3629
timestamp 1712622712
transform 1 0 2340 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3630
timestamp 1712622712
transform 1 0 2260 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3631
timestamp 1712622712
transform 1 0 3100 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1712622712
transform 1 0 3084 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1712622712
transform 1 0 2748 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1712622712
transform 1 0 2740 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1712622712
transform 1 0 2644 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1712622712
transform 1 0 2644 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3637
timestamp 1712622712
transform 1 0 2620 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3638
timestamp 1712622712
transform 1 0 2492 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3639
timestamp 1712622712
transform 1 0 2404 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3640
timestamp 1712622712
transform 1 0 2388 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1712622712
transform 1 0 2324 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3642
timestamp 1712622712
transform 1 0 2300 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1712622712
transform 1 0 2268 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1712622712
transform 1 0 2428 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1712622712
transform 1 0 2252 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3646
timestamp 1712622712
transform 1 0 2196 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3647
timestamp 1712622712
transform 1 0 2708 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3648
timestamp 1712622712
transform 1 0 2652 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1712622712
transform 1 0 3156 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3650
timestamp 1712622712
transform 1 0 3044 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1712622712
transform 1 0 3036 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3652
timestamp 1712622712
transform 1 0 3028 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1712622712
transform 1 0 2996 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1712622712
transform 1 0 2988 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1712622712
transform 1 0 1788 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1712622712
transform 1 0 1636 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1712622712
transform 1 0 1628 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3658
timestamp 1712622712
transform 1 0 132 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3659
timestamp 1712622712
transform 1 0 148 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3660
timestamp 1712622712
transform 1 0 124 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1712622712
transform 1 0 116 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1712622712
transform 1 0 84 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_3663
timestamp 1712622712
transform 1 0 132 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1712622712
transform 1 0 84 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3665
timestamp 1712622712
transform 1 0 124 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1712622712
transform 1 0 124 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3667
timestamp 1712622712
transform 1 0 700 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1712622712
transform 1 0 132 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3669
timestamp 1712622712
transform 1 0 2140 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3670
timestamp 1712622712
transform 1 0 1676 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_3671
timestamp 1712622712
transform 1 0 1676 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3672
timestamp 1712622712
transform 1 0 1276 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3673
timestamp 1712622712
transform 1 0 1276 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_3674
timestamp 1712622712
transform 1 0 1212 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1712622712
transform 1 0 1212 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1712622712
transform 1 0 740 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3677
timestamp 1712622712
transform 1 0 580 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3678
timestamp 1712622712
transform 1 0 572 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3679
timestamp 1712622712
transform 1 0 372 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3680
timestamp 1712622712
transform 1 0 332 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3681
timestamp 1712622712
transform 1 0 108 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3682
timestamp 1712622712
transform 1 0 140 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1712622712
transform 1 0 108 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3684
timestamp 1712622712
transform 1 0 1004 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3685
timestamp 1712622712
transform 1 0 748 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1712622712
transform 1 0 148 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3687
timestamp 1712622712
transform 1 0 84 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1712622712
transform 1 0 156 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3689
timestamp 1712622712
transform 1 0 84 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3690
timestamp 1712622712
transform 1 0 140 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3691
timestamp 1712622712
transform 1 0 140 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1712622712
transform 1 0 84 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1712622712
transform 1 0 84 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3694
timestamp 1712622712
transform 1 0 196 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3695
timestamp 1712622712
transform 1 0 108 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3696
timestamp 1712622712
transform 1 0 236 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1712622712
transform 1 0 124 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1712622712
transform 1 0 540 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3699
timestamp 1712622712
transform 1 0 228 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3700
timestamp 1712622712
transform 1 0 252 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3701
timestamp 1712622712
transform 1 0 204 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3702
timestamp 1712622712
transform 1 0 100 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3703
timestamp 1712622712
transform 1 0 1164 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3704
timestamp 1712622712
transform 1 0 1140 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3705
timestamp 1712622712
transform 1 0 1268 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3706
timestamp 1712622712
transform 1 0 1220 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1712622712
transform 1 0 1460 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3708
timestamp 1712622712
transform 1 0 1364 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1712622712
transform 1 0 1364 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1712622712
transform 1 0 1244 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3711
timestamp 1712622712
transform 1 0 1196 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3712
timestamp 1712622712
transform 1 0 1348 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3713
timestamp 1712622712
transform 1 0 1308 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1712622712
transform 1 0 1244 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1712622712
transform 1 0 1436 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3716
timestamp 1712622712
transform 1 0 1348 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3717
timestamp 1712622712
transform 1 0 1164 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3718
timestamp 1712622712
transform 1 0 1156 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3719
timestamp 1712622712
transform 1 0 1132 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3720
timestamp 1712622712
transform 1 0 1620 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3721
timestamp 1712622712
transform 1 0 1508 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3722
timestamp 1712622712
transform 1 0 1340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3723
timestamp 1712622712
transform 1 0 1292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1712622712
transform 1 0 1292 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1712622712
transform 1 0 1156 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3726
timestamp 1712622712
transform 1 0 1924 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1712622712
transform 1 0 1756 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3728
timestamp 1712622712
transform 1 0 1908 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3729
timestamp 1712622712
transform 1 0 1748 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1712622712
transform 1 0 2068 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3731
timestamp 1712622712
transform 1 0 1932 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1712622712
transform 1 0 1932 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1712622712
transform 1 0 1532 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1712622712
transform 1 0 1364 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3735
timestamp 1712622712
transform 1 0 2508 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3736
timestamp 1712622712
transform 1 0 2508 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3737
timestamp 1712622712
transform 1 0 2444 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1712622712
transform 1 0 2428 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3739
timestamp 1712622712
transform 1 0 2404 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3740
timestamp 1712622712
transform 1 0 2108 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1712622712
transform 1 0 1996 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3742
timestamp 1712622712
transform 1 0 1996 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3743
timestamp 1712622712
transform 1 0 1996 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1712622712
transform 1 0 1980 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3745
timestamp 1712622712
transform 1 0 1980 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3746
timestamp 1712622712
transform 1 0 1956 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1712622712
transform 1 0 1948 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3748
timestamp 1712622712
transform 1 0 1948 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3749
timestamp 1712622712
transform 1 0 1924 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3750
timestamp 1712622712
transform 1 0 1916 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3751
timestamp 1712622712
transform 1 0 1916 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3752
timestamp 1712622712
transform 1 0 1844 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3753
timestamp 1712622712
transform 1 0 1796 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1712622712
transform 1 0 2108 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3755
timestamp 1712622712
transform 1 0 1996 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3756
timestamp 1712622712
transform 1 0 1972 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1712622712
transform 1 0 1724 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3758
timestamp 1712622712
transform 1 0 2964 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3759
timestamp 1712622712
transform 1 0 2604 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3760
timestamp 1712622712
transform 1 0 2556 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3761
timestamp 1712622712
transform 1 0 2532 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3762
timestamp 1712622712
transform 1 0 2532 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3763
timestamp 1712622712
transform 1 0 2444 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3764
timestamp 1712622712
transform 1 0 2444 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3765
timestamp 1712622712
transform 1 0 2324 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3766
timestamp 1712622712
transform 1 0 2276 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3767
timestamp 1712622712
transform 1 0 2196 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3768
timestamp 1712622712
transform 1 0 2172 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3769
timestamp 1712622712
transform 1 0 2172 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3770
timestamp 1712622712
transform 1 0 2172 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3771
timestamp 1712622712
transform 1 0 2068 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3772
timestamp 1712622712
transform 1 0 2052 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3773
timestamp 1712622712
transform 1 0 2052 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3774
timestamp 1712622712
transform 1 0 2044 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3775
timestamp 1712622712
transform 1 0 2028 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3776
timestamp 1712622712
transform 1 0 2180 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3777
timestamp 1712622712
transform 1 0 2092 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3778
timestamp 1712622712
transform 1 0 2156 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3779
timestamp 1712622712
transform 1 0 2052 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1712622712
transform 1 0 1724 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3781
timestamp 1712622712
transform 1 0 1604 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3782
timestamp 1712622712
transform 1 0 2244 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3783
timestamp 1712622712
transform 1 0 1740 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1712622712
transform 1 0 2220 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3785
timestamp 1712622712
transform 1 0 2148 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3786
timestamp 1712622712
transform 1 0 1956 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3787
timestamp 1712622712
transform 1 0 1820 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3788
timestamp 1712622712
transform 1 0 1820 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3789
timestamp 1712622712
transform 1 0 1740 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3790
timestamp 1712622712
transform 1 0 1740 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3791
timestamp 1712622712
transform 1 0 1588 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3792
timestamp 1712622712
transform 1 0 1612 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3793
timestamp 1712622712
transform 1 0 1148 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1712622712
transform 1 0 1148 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3795
timestamp 1712622712
transform 1 0 1052 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3796
timestamp 1712622712
transform 1 0 1052 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1712622712
transform 1 0 1036 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1712622712
transform 1 0 804 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3799
timestamp 1712622712
transform 1 0 804 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1712622712
transform 1 0 676 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1712622712
transform 1 0 652 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3802
timestamp 1712622712
transform 1 0 2108 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3803
timestamp 1712622712
transform 1 0 1940 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3804
timestamp 1712622712
transform 1 0 1948 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3805
timestamp 1712622712
transform 1 0 1908 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3806
timestamp 1712622712
transform 1 0 1932 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3807
timestamp 1712622712
transform 1 0 1804 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3808
timestamp 1712622712
transform 1 0 1964 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3809
timestamp 1712622712
transform 1 0 1884 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3810
timestamp 1712622712
transform 1 0 1532 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_3811
timestamp 1712622712
transform 1 0 1404 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_3812
timestamp 1712622712
transform 1 0 1596 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1712622712
transform 1 0 1500 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1712622712
transform 1 0 1492 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1712622712
transform 1 0 1444 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3816
timestamp 1712622712
transform 1 0 1276 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3817
timestamp 1712622712
transform 1 0 1164 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3818
timestamp 1712622712
transform 1 0 1084 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3819
timestamp 1712622712
transform 1 0 1084 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3820
timestamp 1712622712
transform 1 0 972 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3821
timestamp 1712622712
transform 1 0 940 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1712622712
transform 1 0 908 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1712622712
transform 1 0 892 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3824
timestamp 1712622712
transform 1 0 804 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1712622712
transform 1 0 524 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1712622712
transform 1 0 3212 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1712622712
transform 1 0 2716 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1712622712
transform 1 0 2700 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1712622712
transform 1 0 1572 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1712622712
transform 1 0 1564 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_3831
timestamp 1712622712
transform 1 0 1404 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1712622712
transform 1 0 1732 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3833
timestamp 1712622712
transform 1 0 1636 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1712622712
transform 1 0 1300 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3835
timestamp 1712622712
transform 1 0 1236 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3836
timestamp 1712622712
transform 1 0 1212 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1712622712
transform 1 0 1180 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1712622712
transform 1 0 1148 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1712622712
transform 1 0 1148 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1712622712
transform 1 0 1124 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3841
timestamp 1712622712
transform 1 0 1268 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3842
timestamp 1712622712
transform 1 0 1260 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1712622712
transform 1 0 1236 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3844
timestamp 1712622712
transform 1 0 1172 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3845
timestamp 1712622712
transform 1 0 868 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3846
timestamp 1712622712
transform 1 0 1372 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1712622712
transform 1 0 1340 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1712622712
transform 1 0 1332 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3849
timestamp 1712622712
transform 1 0 1308 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1712622712
transform 1 0 1356 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1712622712
transform 1 0 1220 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3852
timestamp 1712622712
transform 1 0 1212 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3853
timestamp 1712622712
transform 1 0 1196 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3854
timestamp 1712622712
transform 1 0 1028 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3855
timestamp 1712622712
transform 1 0 1028 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1712622712
transform 1 0 716 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3857
timestamp 1712622712
transform 1 0 716 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3858
timestamp 1712622712
transform 1 0 524 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3859
timestamp 1712622712
transform 1 0 1292 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3860
timestamp 1712622712
transform 1 0 956 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3861
timestamp 1712622712
transform 1 0 1364 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3862
timestamp 1712622712
transform 1 0 1260 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3863
timestamp 1712622712
transform 1 0 1100 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3864
timestamp 1712622712
transform 1 0 812 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3865
timestamp 1712622712
transform 1 0 812 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3866
timestamp 1712622712
transform 1 0 540 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3867
timestamp 1712622712
transform 1 0 532 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3868
timestamp 1712622712
transform 1 0 412 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3869
timestamp 1712622712
transform 1 0 332 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3870
timestamp 1712622712
transform 1 0 1164 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3871
timestamp 1712622712
transform 1 0 1116 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3872
timestamp 1712622712
transform 1 0 1068 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3873
timestamp 1712622712
transform 1 0 1428 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3874
timestamp 1712622712
transform 1 0 1380 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3875
timestamp 1712622712
transform 1 0 1004 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3876
timestamp 1712622712
transform 1 0 980 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3877
timestamp 1712622712
transform 1 0 908 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3878
timestamp 1712622712
transform 1 0 876 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3879
timestamp 1712622712
transform 1 0 876 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3880
timestamp 1712622712
transform 1 0 860 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3881
timestamp 1712622712
transform 1 0 788 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3882
timestamp 1712622712
transform 1 0 788 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3883
timestamp 1712622712
transform 1 0 1108 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_3884
timestamp 1712622712
transform 1 0 780 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1712622712
transform 1 0 1412 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3886
timestamp 1712622712
transform 1 0 1084 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3887
timestamp 1712622712
transform 1 0 1164 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1712622712
transform 1 0 1092 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1712622712
transform 1 0 1116 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1712622712
transform 1 0 1020 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3891
timestamp 1712622712
transform 1 0 1020 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3892
timestamp 1712622712
transform 1 0 868 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3893
timestamp 1712622712
transform 1 0 868 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3894
timestamp 1712622712
transform 1 0 812 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3895
timestamp 1712622712
transform 1 0 396 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3896
timestamp 1712622712
transform 1 0 396 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3897
timestamp 1712622712
transform 1 0 372 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3898
timestamp 1712622712
transform 1 0 308 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1712622712
transform 1 0 300 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3900
timestamp 1712622712
transform 1 0 300 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3901
timestamp 1712622712
transform 1 0 284 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1712622712
transform 1 0 1180 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3903
timestamp 1712622712
transform 1 0 1108 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3904
timestamp 1712622712
transform 1 0 1068 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3905
timestamp 1712622712
transform 1 0 3260 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3906
timestamp 1712622712
transform 1 0 3140 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3907
timestamp 1712622712
transform 1 0 3068 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3908
timestamp 1712622712
transform 1 0 3004 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1712622712
transform 1 0 868 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3910
timestamp 1712622712
transform 1 0 716 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3911
timestamp 1712622712
transform 1 0 1372 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3912
timestamp 1712622712
transform 1 0 1188 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3913
timestamp 1712622712
transform 1 0 1188 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3914
timestamp 1712622712
transform 1 0 844 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3915
timestamp 1712622712
transform 1 0 1004 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3916
timestamp 1712622712
transform 1 0 932 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3917
timestamp 1712622712
transform 1 0 932 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1712622712
transform 1 0 852 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1712622712
transform 1 0 1268 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3920
timestamp 1712622712
transform 1 0 1164 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3921
timestamp 1712622712
transform 1 0 1164 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3922
timestamp 1712622712
transform 1 0 1156 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3923
timestamp 1712622712
transform 1 0 1132 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1712622712
transform 1 0 964 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3925
timestamp 1712622712
transform 1 0 932 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3926
timestamp 1712622712
transform 1 0 932 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1712622712
transform 1 0 924 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1712622712
transform 1 0 860 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1712622712
transform 1 0 1236 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3930
timestamp 1712622712
transform 1 0 1188 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3931
timestamp 1712622712
transform 1 0 2852 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1712622712
transform 1 0 2316 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1712622712
transform 1 0 1740 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3934
timestamp 1712622712
transform 1 0 1740 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3935
timestamp 1712622712
transform 1 0 1468 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3936
timestamp 1712622712
transform 1 0 1340 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3937
timestamp 1712622712
transform 1 0 1252 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1712622712
transform 1 0 1252 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1712622712
transform 1 0 1212 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1712622712
transform 1 0 3004 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3941
timestamp 1712622712
transform 1 0 3004 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1712622712
transform 1 0 2900 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1712622712
transform 1 0 1660 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1712622712
transform 1 0 1444 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1712622712
transform 1 0 1444 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1712622712
transform 1 0 1348 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1712622712
transform 1 0 1324 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3948
timestamp 1712622712
transform 1 0 1260 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3949
timestamp 1712622712
transform 1 0 1228 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1712622712
transform 1 0 1220 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1712622712
transform 1 0 1348 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1712622712
transform 1 0 1324 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3953
timestamp 1712622712
transform 1 0 1420 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1712622712
transform 1 0 1348 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3955
timestamp 1712622712
transform 1 0 1124 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3956
timestamp 1712622712
transform 1 0 1084 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3957
timestamp 1712622712
transform 1 0 1084 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1712622712
transform 1 0 1084 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3959
timestamp 1712622712
transform 1 0 1068 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3960
timestamp 1712622712
transform 1 0 1004 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1712622712
transform 1 0 908 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3962
timestamp 1712622712
transform 1 0 1540 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1712622712
transform 1 0 1436 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1712622712
transform 1 0 604 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3965
timestamp 1712622712
transform 1 0 516 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3966
timestamp 1712622712
transform 1 0 812 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3967
timestamp 1712622712
transform 1 0 596 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3968
timestamp 1712622712
transform 1 0 924 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3969
timestamp 1712622712
transform 1 0 788 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3970
timestamp 1712622712
transform 1 0 1132 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3971
timestamp 1712622712
transform 1 0 1100 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3972
timestamp 1712622712
transform 1 0 980 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3973
timestamp 1712622712
transform 1 0 940 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3974
timestamp 1712622712
transform 1 0 748 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3975
timestamp 1712622712
transform 1 0 740 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3976
timestamp 1712622712
transform 1 0 732 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3977
timestamp 1712622712
transform 1 0 308 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3978
timestamp 1712622712
transform 1 0 300 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3979
timestamp 1712622712
transform 1 0 236 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3980
timestamp 1712622712
transform 1 0 884 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3981
timestamp 1712622712
transform 1 0 764 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3982
timestamp 1712622712
transform 1 0 1244 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3983
timestamp 1712622712
transform 1 0 1116 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3984
timestamp 1712622712
transform 1 0 1156 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3985
timestamp 1712622712
transform 1 0 1132 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3986
timestamp 1712622712
transform 1 0 1572 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3987
timestamp 1712622712
transform 1 0 1556 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3988
timestamp 1712622712
transform 1 0 1268 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3989
timestamp 1712622712
transform 1 0 1196 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3990
timestamp 1712622712
transform 1 0 940 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3991
timestamp 1712622712
transform 1 0 1228 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1712622712
transform 1 0 1188 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3993
timestamp 1712622712
transform 1 0 2820 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1712622712
transform 1 0 2788 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3995
timestamp 1712622712
transform 1 0 2708 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3996
timestamp 1712622712
transform 1 0 1788 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3997
timestamp 1712622712
transform 1 0 1788 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3998
timestamp 1712622712
transform 1 0 1684 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3999
timestamp 1712622712
transform 1 0 1636 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4000
timestamp 1712622712
transform 1 0 1628 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4001
timestamp 1712622712
transform 1 0 1388 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4002
timestamp 1712622712
transform 1 0 1388 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4003
timestamp 1712622712
transform 1 0 1364 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4004
timestamp 1712622712
transform 1 0 1356 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4005
timestamp 1712622712
transform 1 0 1276 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4006
timestamp 1712622712
transform 1 0 972 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4007
timestamp 1712622712
transform 1 0 668 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4008
timestamp 1712622712
transform 1 0 628 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4009
timestamp 1712622712
transform 1 0 3012 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4010
timestamp 1712622712
transform 1 0 3004 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4011
timestamp 1712622712
transform 1 0 2964 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4012
timestamp 1712622712
transform 1 0 2876 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4013
timestamp 1712622712
transform 1 0 2876 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4014
timestamp 1712622712
transform 1 0 2716 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1712622712
transform 1 0 2716 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_4016
timestamp 1712622712
transform 1 0 2500 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4017
timestamp 1712622712
transform 1 0 1196 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4018
timestamp 1712622712
transform 1 0 940 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1712622712
transform 1 0 940 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4020
timestamp 1712622712
transform 1 0 940 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4021
timestamp 1712622712
transform 1 0 916 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4022
timestamp 1712622712
transform 1 0 916 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_4023
timestamp 1712622712
transform 1 0 868 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4024
timestamp 1712622712
transform 1 0 860 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1712622712
transform 1 0 860 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4026
timestamp 1712622712
transform 1 0 860 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4027
timestamp 1712622712
transform 1 0 820 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4028
timestamp 1712622712
transform 1 0 820 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4029
timestamp 1712622712
transform 1 0 812 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4030
timestamp 1712622712
transform 1 0 1092 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4031
timestamp 1712622712
transform 1 0 1044 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4032
timestamp 1712622712
transform 1 0 980 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4033
timestamp 1712622712
transform 1 0 1628 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4034
timestamp 1712622712
transform 1 0 1580 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4035
timestamp 1712622712
transform 1 0 1116 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4036
timestamp 1712622712
transform 1 0 1116 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4037
timestamp 1712622712
transform 1 0 1116 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4038
timestamp 1712622712
transform 1 0 1044 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1712622712
transform 1 0 916 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4040
timestamp 1712622712
transform 1 0 1268 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1712622712
transform 1 0 1052 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4042
timestamp 1712622712
transform 1 0 428 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4043
timestamp 1712622712
transform 1 0 396 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4044
timestamp 1712622712
transform 1 0 668 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4045
timestamp 1712622712
transform 1 0 436 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4046
timestamp 1712622712
transform 1 0 1244 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4047
timestamp 1712622712
transform 1 0 668 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4048
timestamp 1712622712
transform 1 0 588 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4049
timestamp 1712622712
transform 1 0 572 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4050
timestamp 1712622712
transform 1 0 524 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4051
timestamp 1712622712
transform 1 0 524 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4052
timestamp 1712622712
transform 1 0 484 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4053
timestamp 1712622712
transform 1 0 484 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4054
timestamp 1712622712
transform 1 0 484 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4055
timestamp 1712622712
transform 1 0 468 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4056
timestamp 1712622712
transform 1 0 468 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4057
timestamp 1712622712
transform 1 0 452 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4058
timestamp 1712622712
transform 1 0 412 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4059
timestamp 1712622712
transform 1 0 316 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4060
timestamp 1712622712
transform 1 0 316 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4061
timestamp 1712622712
transform 1 0 276 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4062
timestamp 1712622712
transform 1 0 644 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4063
timestamp 1712622712
transform 1 0 572 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4064
timestamp 1712622712
transform 1 0 540 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4065
timestamp 1712622712
transform 1 0 540 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4066
timestamp 1712622712
transform 1 0 492 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4067
timestamp 1712622712
transform 1 0 492 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4068
timestamp 1712622712
transform 1 0 468 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4069
timestamp 1712622712
transform 1 0 708 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4070
timestamp 1712622712
transform 1 0 508 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4071
timestamp 1712622712
transform 1 0 380 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4072
timestamp 1712622712
transform 1 0 772 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4073
timestamp 1712622712
transform 1 0 700 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4074
timestamp 1712622712
transform 1 0 700 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1712622712
transform 1 0 668 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4076
timestamp 1712622712
transform 1 0 324 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4077
timestamp 1712622712
transform 1 0 196 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4078
timestamp 1712622712
transform 1 0 1980 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4079
timestamp 1712622712
transform 1 0 1380 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4080
timestamp 1712622712
transform 1 0 1380 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4081
timestamp 1712622712
transform 1 0 1300 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4082
timestamp 1712622712
transform 1 0 796 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4083
timestamp 1712622712
transform 1 0 796 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4084
timestamp 1712622712
transform 1 0 788 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4085
timestamp 1712622712
transform 1 0 740 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4086
timestamp 1712622712
transform 1 0 708 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4087
timestamp 1712622712
transform 1 0 2892 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1712622712
transform 1 0 2892 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4089
timestamp 1712622712
transform 1 0 2836 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4090
timestamp 1712622712
transform 1 0 1868 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4091
timestamp 1712622712
transform 1 0 1828 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4092
timestamp 1712622712
transform 1 0 1820 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4093
timestamp 1712622712
transform 1 0 1740 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4094
timestamp 1712622712
transform 1 0 1500 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1712622712
transform 1 0 1004 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4096
timestamp 1712622712
transform 1 0 2940 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4097
timestamp 1712622712
transform 1 0 2940 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4098
timestamp 1712622712
transform 1 0 2908 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1712622712
transform 1 0 2252 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4100
timestamp 1712622712
transform 1 0 1252 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1712622712
transform 1 0 628 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4102
timestamp 1712622712
transform 1 0 604 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4103
timestamp 1712622712
transform 1 0 604 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1712622712
transform 1 0 2036 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4105
timestamp 1712622712
transform 1 0 1508 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4106
timestamp 1712622712
transform 1 0 1508 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4107
timestamp 1712622712
transform 1 0 1396 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4108
timestamp 1712622712
transform 1 0 748 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4109
timestamp 1712622712
transform 1 0 748 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4110
timestamp 1712622712
transform 1 0 684 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4111
timestamp 1712622712
transform 1 0 684 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1712622712
transform 1 0 652 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4113
timestamp 1712622712
transform 1 0 1100 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4114
timestamp 1712622712
transform 1 0 980 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1712622712
transform 1 0 956 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4116
timestamp 1712622712
transform 1 0 836 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4117
timestamp 1712622712
transform 1 0 724 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4118
timestamp 1712622712
transform 1 0 716 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4119
timestamp 1712622712
transform 1 0 2748 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1712622712
transform 1 0 1340 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4121
timestamp 1712622712
transform 1 0 1300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4122
timestamp 1712622712
transform 1 0 1300 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4123
timestamp 1712622712
transform 1 0 1292 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4124
timestamp 1712622712
transform 1 0 1268 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4125
timestamp 1712622712
transform 1 0 1244 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4126
timestamp 1712622712
transform 1 0 1180 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4127
timestamp 1712622712
transform 1 0 1180 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4128
timestamp 1712622712
transform 1 0 1140 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4129
timestamp 1712622712
transform 1 0 1140 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4130
timestamp 1712622712
transform 1 0 1140 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4131
timestamp 1712622712
transform 1 0 1124 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4132
timestamp 1712622712
transform 1 0 260 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4133
timestamp 1712622712
transform 1 0 188 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4134
timestamp 1712622712
transform 1 0 580 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4135
timestamp 1712622712
transform 1 0 356 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4136
timestamp 1712622712
transform 1 0 924 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4137
timestamp 1712622712
transform 1 0 372 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4138
timestamp 1712622712
transform 1 0 996 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4139
timestamp 1712622712
transform 1 0 820 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4140
timestamp 1712622712
transform 1 0 820 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4141
timestamp 1712622712
transform 1 0 340 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4142
timestamp 1712622712
transform 1 0 340 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1712622712
transform 1 0 268 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1712622712
transform 1 0 212 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4145
timestamp 1712622712
transform 1 0 108 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1712622712
transform 1 0 100 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4147
timestamp 1712622712
transform 1 0 1036 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4148
timestamp 1712622712
transform 1 0 628 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4149
timestamp 1712622712
transform 1 0 628 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4150
timestamp 1712622712
transform 1 0 156 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4151
timestamp 1712622712
transform 1 0 156 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4152
timestamp 1712622712
transform 1 0 68 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1712622712
transform 1 0 1988 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4154
timestamp 1712622712
transform 1 0 1556 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4155
timestamp 1712622712
transform 1 0 1028 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4156
timestamp 1712622712
transform 1 0 1020 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4157
timestamp 1712622712
transform 1 0 1004 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1712622712
transform 1 0 956 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4159
timestamp 1712622712
transform 1 0 956 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4160
timestamp 1712622712
transform 1 0 1068 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4161
timestamp 1712622712
transform 1 0 1036 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4162
timestamp 1712622712
transform 1 0 2812 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4163
timestamp 1712622712
transform 1 0 2516 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4164
timestamp 1712622712
transform 1 0 2516 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4165
timestamp 1712622712
transform 1 0 2444 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4166
timestamp 1712622712
transform 1 0 2444 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1712622712
transform 1 0 2388 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4168
timestamp 1712622712
transform 1 0 1588 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4169
timestamp 1712622712
transform 1 0 876 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4170
timestamp 1712622712
transform 1 0 1900 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4171
timestamp 1712622712
transform 1 0 1780 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4172
timestamp 1712622712
transform 1 0 1780 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4173
timestamp 1712622712
transform 1 0 1700 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4174
timestamp 1712622712
transform 1 0 988 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4175
timestamp 1712622712
transform 1 0 988 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4176
timestamp 1712622712
transform 1 0 980 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4177
timestamp 1712622712
transform 1 0 964 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4178
timestamp 1712622712
transform 1 0 924 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4179
timestamp 1712622712
transform 1 0 1068 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4180
timestamp 1712622712
transform 1 0 924 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4181
timestamp 1712622712
transform 1 0 924 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4182
timestamp 1712622712
transform 1 0 876 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4183
timestamp 1712622712
transform 1 0 564 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1712622712
transform 1 0 276 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4185
timestamp 1712622712
transform 1 0 276 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4186
timestamp 1712622712
transform 1 0 220 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4187
timestamp 1712622712
transform 1 0 220 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4188
timestamp 1712622712
transform 1 0 572 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1712622712
transform 1 0 292 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4190
timestamp 1712622712
transform 1 0 436 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4191
timestamp 1712622712
transform 1 0 308 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4192
timestamp 1712622712
transform 1 0 1228 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4193
timestamp 1712622712
transform 1 0 732 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4194
timestamp 1712622712
transform 1 0 604 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4195
timestamp 1712622712
transform 1 0 364 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1712622712
transform 1 0 364 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4197
timestamp 1712622712
transform 1 0 364 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4198
timestamp 1712622712
transform 1 0 364 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4199
timestamp 1712622712
transform 1 0 332 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4200
timestamp 1712622712
transform 1 0 324 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1712622712
transform 1 0 316 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1712622712
transform 1 0 316 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4203
timestamp 1712622712
transform 1 0 300 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4204
timestamp 1712622712
transform 1 0 804 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4205
timestamp 1712622712
transform 1 0 356 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4206
timestamp 1712622712
transform 1 0 1004 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4207
timestamp 1712622712
transform 1 0 356 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4208
timestamp 1712622712
transform 1 0 268 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4209
timestamp 1712622712
transform 1 0 268 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1712622712
transform 1 0 188 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1712622712
transform 1 0 188 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4212
timestamp 1712622712
transform 1 0 132 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4213
timestamp 1712622712
transform 1 0 892 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1712622712
transform 1 0 596 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1712622712
transform 1 0 620 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4216
timestamp 1712622712
transform 1 0 572 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4217
timestamp 1712622712
transform 1 0 124 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4218
timestamp 1712622712
transform 1 0 116 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4219
timestamp 1712622712
transform 1 0 188 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4220
timestamp 1712622712
transform 1 0 116 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4221
timestamp 1712622712
transform 1 0 284 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4222
timestamp 1712622712
transform 1 0 236 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4223
timestamp 1712622712
transform 1 0 1156 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4224
timestamp 1712622712
transform 1 0 820 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1712622712
transform 1 0 1172 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4226
timestamp 1712622712
transform 1 0 1148 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4227
timestamp 1712622712
transform 1 0 1140 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4228
timestamp 1712622712
transform 1 0 1076 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4229
timestamp 1712622712
transform 1 0 1068 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4230
timestamp 1712622712
transform 1 0 1004 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4231
timestamp 1712622712
transform 1 0 892 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1712622712
transform 1 0 708 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4233
timestamp 1712622712
transform 1 0 1164 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4234
timestamp 1712622712
transform 1 0 980 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4235
timestamp 1712622712
transform 1 0 1124 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4236
timestamp 1712622712
transform 1 0 980 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4237
timestamp 1712622712
transform 1 0 1100 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1712622712
transform 1 0 940 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4239
timestamp 1712622712
transform 1 0 916 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1712622712
transform 1 0 916 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4241
timestamp 1712622712
transform 1 0 916 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4242
timestamp 1712622712
transform 1 0 876 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4243
timestamp 1712622712
transform 1 0 804 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4244
timestamp 1712622712
transform 1 0 804 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4245
timestamp 1712622712
transform 1 0 644 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4246
timestamp 1712622712
transform 1 0 1748 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4247
timestamp 1712622712
transform 1 0 1380 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4248
timestamp 1712622712
transform 1 0 1244 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4249
timestamp 1712622712
transform 1 0 1156 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4250
timestamp 1712622712
transform 1 0 1156 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4251
timestamp 1712622712
transform 1 0 1140 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4252
timestamp 1712622712
transform 1 0 1140 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4253
timestamp 1712622712
transform 1 0 356 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1712622712
transform 1 0 220 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4255
timestamp 1712622712
transform 1 0 572 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4256
timestamp 1712622712
transform 1 0 356 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4257
timestamp 1712622712
transform 1 0 436 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4258
timestamp 1712622712
transform 1 0 420 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4259
timestamp 1712622712
transform 1 0 708 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1712622712
transform 1 0 500 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4261
timestamp 1712622712
transform 1 0 500 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4262
timestamp 1712622712
transform 1 0 452 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4263
timestamp 1712622712
transform 1 0 1204 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_4264
timestamp 1712622712
transform 1 0 692 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4265
timestamp 1712622712
transform 1 0 620 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4266
timestamp 1712622712
transform 1 0 420 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_4267
timestamp 1712622712
transform 1 0 396 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4268
timestamp 1712622712
transform 1 0 324 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4269
timestamp 1712622712
transform 1 0 324 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4270
timestamp 1712622712
transform 1 0 244 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4271
timestamp 1712622712
transform 1 0 228 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4272
timestamp 1712622712
transform 1 0 228 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4273
timestamp 1712622712
transform 1 0 196 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4274
timestamp 1712622712
transform 1 0 92 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4275
timestamp 1712622712
transform 1 0 84 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1712622712
transform 1 0 724 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4277
timestamp 1712622712
transform 1 0 596 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4278
timestamp 1712622712
transform 1 0 836 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1712622712
transform 1 0 772 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4280
timestamp 1712622712
transform 1 0 732 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4281
timestamp 1712622712
transform 1 0 692 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4282
timestamp 1712622712
transform 1 0 212 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4283
timestamp 1712622712
transform 1 0 116 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4284
timestamp 1712622712
transform 1 0 820 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4285
timestamp 1712622712
transform 1 0 308 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4286
timestamp 1712622712
transform 1 0 916 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4287
timestamp 1712622712
transform 1 0 796 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4288
timestamp 1712622712
transform 1 0 852 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4289
timestamp 1712622712
transform 1 0 628 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4290
timestamp 1712622712
transform 1 0 1036 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4291
timestamp 1712622712
transform 1 0 924 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4292
timestamp 1712622712
transform 1 0 2820 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4293
timestamp 1712622712
transform 1 0 2772 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4294
timestamp 1712622712
transform 1 0 1916 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4295
timestamp 1712622712
transform 1 0 1916 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4296
timestamp 1712622712
transform 1 0 1772 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4297
timestamp 1712622712
transform 1 0 1564 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1712622712
transform 1 0 1380 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4299
timestamp 1712622712
transform 1 0 1276 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4300
timestamp 1712622712
transform 1 0 1172 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1712622712
transform 1 0 164 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_4302
timestamp 1712622712
transform 1 0 132 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_4303
timestamp 1712622712
transform 1 0 420 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4304
timestamp 1712622712
transform 1 0 156 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4305
timestamp 1712622712
transform 1 0 564 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1712622712
transform 1 0 460 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4307
timestamp 1712622712
transform 1 0 668 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4308
timestamp 1712622712
transform 1 0 628 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4309
timestamp 1712622712
transform 1 0 692 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4310
timestamp 1712622712
transform 1 0 660 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4311
timestamp 1712622712
transform 1 0 620 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4312
timestamp 1712622712
transform 1 0 140 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4313
timestamp 1712622712
transform 1 0 108 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4314
timestamp 1712622712
transform 1 0 252 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4315
timestamp 1712622712
transform 1 0 188 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4316
timestamp 1712622712
transform 1 0 652 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4317
timestamp 1712622712
transform 1 0 452 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4318
timestamp 1712622712
transform 1 0 740 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4319
timestamp 1712622712
transform 1 0 164 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4320
timestamp 1712622712
transform 1 0 852 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4321
timestamp 1712622712
transform 1 0 716 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4322
timestamp 1712622712
transform 1 0 812 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1712622712
transform 1 0 756 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4324
timestamp 1712622712
transform 1 0 860 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4325
timestamp 1712622712
transform 1 0 804 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4326
timestamp 1712622712
transform 1 0 956 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4327
timestamp 1712622712
transform 1 0 892 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4328
timestamp 1712622712
transform 1 0 892 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4329
timestamp 1712622712
transform 1 0 756 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1712622712
transform 1 0 948 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4331
timestamp 1712622712
transform 1 0 852 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4332
timestamp 1712622712
transform 1 0 276 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1712622712
transform 1 0 116 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4334
timestamp 1712622712
transform 1 0 524 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4335
timestamp 1712622712
transform 1 0 292 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4336
timestamp 1712622712
transform 1 0 428 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4337
timestamp 1712622712
transform 1 0 324 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4338
timestamp 1712622712
transform 1 0 620 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4339
timestamp 1712622712
transform 1 0 476 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4340
timestamp 1712622712
transform 1 0 388 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4341
timestamp 1712622712
transform 1 0 1100 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1712622712
transform 1 0 1076 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4343
timestamp 1712622712
transform 1 0 1004 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1712622712
transform 1 0 900 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4345
timestamp 1712622712
transform 1 0 900 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4346
timestamp 1712622712
transform 1 0 460 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4347
timestamp 1712622712
transform 1 0 460 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4348
timestamp 1712622712
transform 1 0 284 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4349
timestamp 1712622712
transform 1 0 284 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4350
timestamp 1712622712
transform 1 0 252 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4351
timestamp 1712622712
transform 1 0 708 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4352
timestamp 1712622712
transform 1 0 460 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4353
timestamp 1712622712
transform 1 0 804 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4354
timestamp 1712622712
transform 1 0 732 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4355
timestamp 1712622712
transform 1 0 588 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4356
timestamp 1712622712
transform 1 0 116 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4357
timestamp 1712622712
transform 1 0 100 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4358
timestamp 1712622712
transform 1 0 204 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4359
timestamp 1712622712
transform 1 0 116 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4360
timestamp 1712622712
transform 1 0 852 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4361
timestamp 1712622712
transform 1 0 116 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4362
timestamp 1712622712
transform 1 0 116 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4363
timestamp 1712622712
transform 1 0 852 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4364
timestamp 1712622712
transform 1 0 780 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4365
timestamp 1712622712
transform 1 0 892 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4366
timestamp 1712622712
transform 1 0 836 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4367
timestamp 1712622712
transform 1 0 892 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4368
timestamp 1712622712
transform 1 0 868 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4369
timestamp 1712622712
transform 1 0 1316 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4370
timestamp 1712622712
transform 1 0 1236 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4371
timestamp 1712622712
transform 1 0 1140 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1712622712
transform 1 0 1052 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4373
timestamp 1712622712
transform 1 0 1052 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4374
timestamp 1712622712
transform 1 0 1020 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4375
timestamp 1712622712
transform 1 0 940 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4376
timestamp 1712622712
transform 1 0 940 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4377
timestamp 1712622712
transform 1 0 868 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4378
timestamp 1712622712
transform 1 0 948 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4379
timestamp 1712622712
transform 1 0 868 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4380
timestamp 1712622712
transform 1 0 2932 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4381
timestamp 1712622712
transform 1 0 2900 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4382
timestamp 1712622712
transform 1 0 2828 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4383
timestamp 1712622712
transform 1 0 2828 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4384
timestamp 1712622712
transform 1 0 2676 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4385
timestamp 1712622712
transform 1 0 2668 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4386
timestamp 1712622712
transform 1 0 2340 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4387
timestamp 1712622712
transform 1 0 1292 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4388
timestamp 1712622712
transform 1 0 1292 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1712622712
transform 1 0 1124 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4390
timestamp 1712622712
transform 1 0 548 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4391
timestamp 1712622712
transform 1 0 420 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4392
timestamp 1712622712
transform 1 0 420 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4393
timestamp 1712622712
transform 1 0 340 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4394
timestamp 1712622712
transform 1 0 340 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4395
timestamp 1712622712
transform 1 0 300 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4396
timestamp 1712622712
transform 1 0 300 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4397
timestamp 1712622712
transform 1 0 260 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4398
timestamp 1712622712
transform 1 0 212 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4399
timestamp 1712622712
transform 1 0 188 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4400
timestamp 1712622712
transform 1 0 524 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1712622712
transform 1 0 228 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4402
timestamp 1712622712
transform 1 0 580 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4403
timestamp 1712622712
transform 1 0 548 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4404
timestamp 1712622712
transform 1 0 564 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4405
timestamp 1712622712
transform 1 0 500 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4406
timestamp 1712622712
transform 1 0 1356 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4407
timestamp 1712622712
transform 1 0 1356 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4408
timestamp 1712622712
transform 1 0 1220 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1712622712
transform 1 0 1220 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4410
timestamp 1712622712
transform 1 0 1148 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4411
timestamp 1712622712
transform 1 0 1068 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4412
timestamp 1712622712
transform 1 0 660 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4413
timestamp 1712622712
transform 1 0 652 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4414
timestamp 1712622712
transform 1 0 436 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4415
timestamp 1712622712
transform 1 0 404 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4416
timestamp 1712622712
transform 1 0 404 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1712622712
transform 1 0 356 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4418
timestamp 1712622712
transform 1 0 644 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1712622712
transform 1 0 452 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4420
timestamp 1712622712
transform 1 0 380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4421
timestamp 1712622712
transform 1 0 948 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1712622712
transform 1 0 380 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4423
timestamp 1712622712
transform 1 0 348 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4424
timestamp 1712622712
transform 1 0 156 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4425
timestamp 1712622712
transform 1 0 844 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4426
timestamp 1712622712
transform 1 0 652 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1712622712
transform 1 0 860 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4428
timestamp 1712622712
transform 1 0 828 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4429
timestamp 1712622712
transform 1 0 1108 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4430
timestamp 1712622712
transform 1 0 668 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1712622712
transform 1 0 1412 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4432
timestamp 1712622712
transform 1 0 1300 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4433
timestamp 1712622712
transform 1 0 1132 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4434
timestamp 1712622712
transform 1 0 1044 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4435
timestamp 1712622712
transform 1 0 1004 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4436
timestamp 1712622712
transform 1 0 1324 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4437
timestamp 1712622712
transform 1 0 956 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4438
timestamp 1712622712
transform 1 0 1052 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4439
timestamp 1712622712
transform 1 0 972 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4440
timestamp 1712622712
transform 1 0 1716 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4441
timestamp 1712622712
transform 1 0 1556 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4442
timestamp 1712622712
transform 1 0 1348 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4443
timestamp 1712622712
transform 1 0 1020 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4444
timestamp 1712622712
transform 1 0 2916 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4445
timestamp 1712622712
transform 1 0 2876 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1712622712
transform 1 0 2436 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1712622712
transform 1 0 1940 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4448
timestamp 1712622712
transform 1 0 1932 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4449
timestamp 1712622712
transform 1 0 1716 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4450
timestamp 1712622712
transform 1 0 1412 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4451
timestamp 1712622712
transform 1 0 1340 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4452
timestamp 1712622712
transform 1 0 1244 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4453
timestamp 1712622712
transform 1 0 1020 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4454
timestamp 1712622712
transform 1 0 2668 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4455
timestamp 1712622712
transform 1 0 2596 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4456
timestamp 1712622712
transform 1 0 1812 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4457
timestamp 1712622712
transform 1 0 1468 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4458
timestamp 1712622712
transform 1 0 1460 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4459
timestamp 1712622712
transform 1 0 1388 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1712622712
transform 1 0 980 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4461
timestamp 1712622712
transform 1 0 228 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4462
timestamp 1712622712
transform 1 0 76 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4463
timestamp 1712622712
transform 1 0 76 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4464
timestamp 1712622712
transform 1 0 788 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1712622712
transform 1 0 244 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1712622712
transform 1 0 452 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4467
timestamp 1712622712
transform 1 0 300 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4468
timestamp 1712622712
transform 1 0 828 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_4469
timestamp 1712622712
transform 1 0 364 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_4470
timestamp 1712622712
transform 1 0 972 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4471
timestamp 1712622712
transform 1 0 524 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4472
timestamp 1712622712
transform 1 0 516 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1712622712
transform 1 0 276 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4474
timestamp 1712622712
transform 1 0 276 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4475
timestamp 1712622712
transform 1 0 196 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4476
timestamp 1712622712
transform 1 0 1036 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4477
timestamp 1712622712
transform 1 0 980 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4478
timestamp 1712622712
transform 1 0 844 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4479
timestamp 1712622712
transform 1 0 956 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4480
timestamp 1712622712
transform 1 0 716 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4481
timestamp 1712622712
transform 1 0 1188 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1712622712
transform 1 0 956 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4483
timestamp 1712622712
transform 1 0 2868 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4484
timestamp 1712622712
transform 1 0 2836 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4485
timestamp 1712622712
transform 1 0 2524 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1712622712
transform 1 0 2492 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4487
timestamp 1712622712
transform 1 0 2468 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4488
timestamp 1712622712
transform 1 0 1796 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4489
timestamp 1712622712
transform 1 0 1788 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4490
timestamp 1712622712
transform 1 0 1524 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4491
timestamp 1712622712
transform 1 0 1396 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4492
timestamp 1712622712
transform 1 0 1108 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4493
timestamp 1712622712
transform 1 0 1124 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4494
timestamp 1712622712
transform 1 0 684 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4495
timestamp 1712622712
transform 1 0 484 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4496
timestamp 1712622712
transform 1 0 484 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4497
timestamp 1712622712
transform 1 0 348 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4498
timestamp 1712622712
transform 1 0 348 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1712622712
transform 1 0 644 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4500
timestamp 1712622712
transform 1 0 436 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1712622712
transform 1 0 684 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4502
timestamp 1712622712
transform 1 0 652 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4503
timestamp 1712622712
transform 1 0 652 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4504
timestamp 1712622712
transform 1 0 532 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4505
timestamp 1712622712
transform 1 0 596 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4506
timestamp 1712622712
transform 1 0 508 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4507
timestamp 1712622712
transform 1 0 708 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4508
timestamp 1712622712
transform 1 0 588 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1712622712
transform 1 0 588 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4510
timestamp 1712622712
transform 1 0 364 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_4511
timestamp 1712622712
transform 1 0 1244 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4512
timestamp 1712622712
transform 1 0 764 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4513
timestamp 1712622712
transform 1 0 748 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4514
timestamp 1712622712
transform 1 0 676 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4515
timestamp 1712622712
transform 1 0 644 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4516
timestamp 1712622712
transform 1 0 524 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_4517
timestamp 1712622712
transform 1 0 412 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_4518
timestamp 1712622712
transform 1 0 420 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4519
timestamp 1712622712
transform 1 0 340 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4520
timestamp 1712622712
transform 1 0 1556 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4521
timestamp 1712622712
transform 1 0 1492 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4522
timestamp 1712622712
transform 1 0 1260 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4523
timestamp 1712622712
transform 1 0 1260 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4524
timestamp 1712622712
transform 1 0 1196 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4525
timestamp 1712622712
transform 1 0 2684 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4526
timestamp 1712622712
transform 1 0 2404 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4527
timestamp 1712622712
transform 1 0 1332 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4528
timestamp 1712622712
transform 1 0 1268 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4529
timestamp 1712622712
transform 1 0 1188 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4530
timestamp 1712622712
transform 1 0 1084 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4531
timestamp 1712622712
transform 1 0 1396 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4532
timestamp 1712622712
transform 1 0 1316 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4533
timestamp 1712622712
transform 1 0 1316 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1712622712
transform 1 0 932 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4535
timestamp 1712622712
transform 1 0 932 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_4536
timestamp 1712622712
transform 1 0 860 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_4537
timestamp 1712622712
transform 1 0 892 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4538
timestamp 1712622712
transform 1 0 820 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4539
timestamp 1712622712
transform 1 0 980 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4540
timestamp 1712622712
transform 1 0 908 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4541
timestamp 1712622712
transform 1 0 2404 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_4542
timestamp 1712622712
transform 1 0 2364 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_4543
timestamp 1712622712
transform 1 0 2236 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_4544
timestamp 1712622712
transform 1 0 2236 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_4545
timestamp 1712622712
transform 1 0 1476 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4546
timestamp 1712622712
transform 1 0 1220 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4547
timestamp 1712622712
transform 1 0 1220 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4548
timestamp 1712622712
transform 1 0 1028 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4549
timestamp 1712622712
transform 1 0 1028 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4550
timestamp 1712622712
transform 1 0 996 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4551
timestamp 1712622712
transform 1 0 972 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4552
timestamp 1712622712
transform 1 0 900 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4553
timestamp 1712622712
transform 1 0 852 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4554
timestamp 1712622712
transform 1 0 852 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4555
timestamp 1712622712
transform 1 0 828 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4556
timestamp 1712622712
transform 1 0 820 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4557
timestamp 1712622712
transform 1 0 596 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4558
timestamp 1712622712
transform 1 0 940 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4559
timestamp 1712622712
transform 1 0 908 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4560
timestamp 1712622712
transform 1 0 836 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4561
timestamp 1712622712
transform 1 0 772 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_4562
timestamp 1712622712
transform 1 0 1284 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4563
timestamp 1712622712
transform 1 0 1116 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4564
timestamp 1712622712
transform 1 0 988 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4565
timestamp 1712622712
transform 1 0 948 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4566
timestamp 1712622712
transform 1 0 916 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4567
timestamp 1712622712
transform 1 0 1044 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4568
timestamp 1712622712
transform 1 0 988 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4569
timestamp 1712622712
transform 1 0 1852 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4570
timestamp 1712622712
transform 1 0 1708 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1712622712
transform 1 0 1692 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1712622712
transform 1 0 1596 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4573
timestamp 1712622712
transform 1 0 1332 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4574
timestamp 1712622712
transform 1 0 1332 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4575
timestamp 1712622712
transform 1 0 1260 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4576
timestamp 1712622712
transform 1 0 1548 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4577
timestamp 1712622712
transform 1 0 1548 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4578
timestamp 1712622712
transform 1 0 1532 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4579
timestamp 1712622712
transform 1 0 1532 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4580
timestamp 1712622712
transform 1 0 1452 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4581
timestamp 1712622712
transform 1 0 1444 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4582
timestamp 1712622712
transform 1 0 1436 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4583
timestamp 1712622712
transform 1 0 1388 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4584
timestamp 1712622712
transform 1 0 1388 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4585
timestamp 1712622712
transform 1 0 1364 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4586
timestamp 1712622712
transform 1 0 1364 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4587
timestamp 1712622712
transform 1 0 1316 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4588
timestamp 1712622712
transform 1 0 1316 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4589
timestamp 1712622712
transform 1 0 1156 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4590
timestamp 1712622712
transform 1 0 1140 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4591
timestamp 1712622712
transform 1 0 1068 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4592
timestamp 1712622712
transform 1 0 1156 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4593
timestamp 1712622712
transform 1 0 1132 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4594
timestamp 1712622712
transform 1 0 1124 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4595
timestamp 1712622712
transform 1 0 1076 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4596
timestamp 1712622712
transform 1 0 1044 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4597
timestamp 1712622712
transform 1 0 1180 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4598
timestamp 1712622712
transform 1 0 1044 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4599
timestamp 1712622712
transform 1 0 1164 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4600
timestamp 1712622712
transform 1 0 1140 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1712622712
transform 1 0 1196 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1712622712
transform 1 0 1156 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1712622712
transform 1 0 1708 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4604
timestamp 1712622712
transform 1 0 1612 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1712622712
transform 1 0 1524 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1712622712
transform 1 0 1428 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4607
timestamp 1712622712
transform 1 0 1380 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4608
timestamp 1712622712
transform 1 0 1204 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1712622712
transform 1 0 1180 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4610
timestamp 1712622712
transform 1 0 1148 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4611
timestamp 1712622712
transform 1 0 1220 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4612
timestamp 1712622712
transform 1 0 1156 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4613
timestamp 1712622712
transform 1 0 2004 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1712622712
transform 1 0 1908 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4615
timestamp 1712622712
transform 1 0 1724 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4616
timestamp 1712622712
transform 1 0 1668 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1712622712
transform 1 0 1492 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4618
timestamp 1712622712
transform 1 0 1420 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4619
timestamp 1712622712
transform 1 0 1180 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1712622712
transform 1 0 1076 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1712622712
transform 1 0 1500 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1712622712
transform 1 0 1300 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1712622712
transform 1 0 1340 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4624
timestamp 1712622712
transform 1 0 1284 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4625
timestamp 1712622712
transform 1 0 1252 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1712622712
transform 1 0 1468 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4627
timestamp 1712622712
transform 1 0 1348 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1712622712
transform 1 0 1284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4629
timestamp 1712622712
transform 1 0 1284 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4630
timestamp 1712622712
transform 1 0 1244 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4631
timestamp 1712622712
transform 1 0 1500 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1712622712
transform 1 0 1420 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1712622712
transform 1 0 1388 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4634
timestamp 1712622712
transform 1 0 1356 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1712622712
transform 1 0 1396 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4636
timestamp 1712622712
transform 1 0 1372 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4637
timestamp 1712622712
transform 1 0 1492 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4638
timestamp 1712622712
transform 1 0 1412 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4639
timestamp 1712622712
transform 1 0 1636 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4640
timestamp 1712622712
transform 1 0 1572 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4641
timestamp 1712622712
transform 1 0 1876 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4642
timestamp 1712622712
transform 1 0 1844 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4643
timestamp 1712622712
transform 1 0 1844 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4644
timestamp 1712622712
transform 1 0 1844 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4645
timestamp 1712622712
transform 1 0 1780 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4646
timestamp 1712622712
transform 1 0 1700 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4647
timestamp 1712622712
transform 1 0 1796 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4648
timestamp 1712622712
transform 1 0 1772 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4649
timestamp 1712622712
transform 1 0 1676 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4650
timestamp 1712622712
transform 1 0 1628 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4651
timestamp 1712622712
transform 1 0 1988 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4652
timestamp 1712622712
transform 1 0 1884 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4653
timestamp 1712622712
transform 1 0 1884 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4654
timestamp 1712622712
transform 1 0 1772 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4655
timestamp 1712622712
transform 1 0 1676 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4656
timestamp 1712622712
transform 1 0 1404 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4657
timestamp 1712622712
transform 1 0 2108 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4658
timestamp 1712622712
transform 1 0 1812 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4659
timestamp 1712622712
transform 1 0 1804 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4660
timestamp 1712622712
transform 1 0 1804 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4661
timestamp 1712622712
transform 1 0 1692 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4662
timestamp 1712622712
transform 1 0 1692 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4663
timestamp 1712622712
transform 1 0 1660 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4664
timestamp 1712622712
transform 1 0 1652 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4665
timestamp 1712622712
transform 1 0 1636 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4666
timestamp 1712622712
transform 1 0 1628 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4667
timestamp 1712622712
transform 1 0 1612 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4668
timestamp 1712622712
transform 1 0 1612 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4669
timestamp 1712622712
transform 1 0 1604 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4670
timestamp 1712622712
transform 1 0 1596 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4671
timestamp 1712622712
transform 1 0 1596 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4672
timestamp 1712622712
transform 1 0 1564 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4673
timestamp 1712622712
transform 1 0 1564 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4674
timestamp 1712622712
transform 1 0 1548 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4675
timestamp 1712622712
transform 1 0 2164 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4676
timestamp 1712622712
transform 1 0 2060 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1712622712
transform 1 0 1972 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4678
timestamp 1712622712
transform 1 0 1932 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4679
timestamp 1712622712
transform 1 0 2108 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_4680
timestamp 1712622712
transform 1 0 2068 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_4681
timestamp 1712622712
transform 1 0 2052 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4682
timestamp 1712622712
transform 1 0 1900 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4683
timestamp 1712622712
transform 1 0 1900 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4684
timestamp 1712622712
transform 1 0 1852 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4685
timestamp 1712622712
transform 1 0 908 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4686
timestamp 1712622712
transform 1 0 604 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4687
timestamp 1712622712
transform 1 0 1948 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1712622712
transform 1 0 1868 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4689
timestamp 1712622712
transform 1 0 1852 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4690
timestamp 1712622712
transform 1 0 2300 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4691
timestamp 1712622712
transform 1 0 2228 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4692
timestamp 1712622712
transform 1 0 2108 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4693
timestamp 1712622712
transform 1 0 2028 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4694
timestamp 1712622712
transform 1 0 1932 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4695
timestamp 1712622712
transform 1 0 1900 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4696
timestamp 1712622712
transform 1 0 2148 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4697
timestamp 1712622712
transform 1 0 1988 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1712622712
transform 1 0 1908 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4699
timestamp 1712622712
transform 1 0 1868 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4700
timestamp 1712622712
transform 1 0 1868 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4701
timestamp 1712622712
transform 1 0 1540 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4702
timestamp 1712622712
transform 1 0 2764 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4703
timestamp 1712622712
transform 1 0 2764 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4704
timestamp 1712622712
transform 1 0 2732 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4705
timestamp 1712622712
transform 1 0 2732 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4706
timestamp 1712622712
transform 1 0 2732 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4707
timestamp 1712622712
transform 1 0 2732 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1712622712
transform 1 0 2732 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4709
timestamp 1712622712
transform 1 0 2732 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4710
timestamp 1712622712
transform 1 0 2260 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4711
timestamp 1712622712
transform 1 0 1900 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4712
timestamp 1712622712
transform 1 0 2460 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4713
timestamp 1712622712
transform 1 0 2388 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4714
timestamp 1712622712
transform 1 0 2236 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4715
timestamp 1712622712
transform 1 0 2444 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4716
timestamp 1712622712
transform 1 0 2444 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4717
timestamp 1712622712
transform 1 0 2412 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4718
timestamp 1712622712
transform 1 0 2148 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4719
timestamp 1712622712
transform 1 0 2148 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4720
timestamp 1712622712
transform 1 0 2068 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4721
timestamp 1712622712
transform 1 0 1892 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4722
timestamp 1712622712
transform 1 0 2068 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4723
timestamp 1712622712
transform 1 0 1884 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4724
timestamp 1712622712
transform 1 0 1836 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4725
timestamp 1712622712
transform 1 0 1716 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4726
timestamp 1712622712
transform 1 0 2260 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1712622712
transform 1 0 2212 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1712622712
transform 1 0 2180 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4729
timestamp 1712622712
transform 1 0 2052 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1712622712
transform 1 0 2420 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1712622712
transform 1 0 2308 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4732
timestamp 1712622712
transform 1 0 2060 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4733
timestamp 1712622712
transform 1 0 1964 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4734
timestamp 1712622712
transform 1 0 1964 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4735
timestamp 1712622712
transform 1 0 1956 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4736
timestamp 1712622712
transform 1 0 1836 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4737
timestamp 1712622712
transform 1 0 1708 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1712622712
transform 1 0 1788 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1712622712
transform 1 0 1700 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4740
timestamp 1712622712
transform 1 0 1796 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4741
timestamp 1712622712
transform 1 0 1580 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4742
timestamp 1712622712
transform 1 0 1804 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4743
timestamp 1712622712
transform 1 0 1692 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4744
timestamp 1712622712
transform 1 0 1540 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4745
timestamp 1712622712
transform 1 0 1540 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4746
timestamp 1712622712
transform 1 0 1500 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4747
timestamp 1712622712
transform 1 0 2300 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4748
timestamp 1712622712
transform 1 0 2260 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4749
timestamp 1712622712
transform 1 0 2244 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4750
timestamp 1712622712
transform 1 0 2244 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4751
timestamp 1712622712
transform 1 0 2244 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4752
timestamp 1712622712
transform 1 0 2212 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4753
timestamp 1712622712
transform 1 0 2212 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4754
timestamp 1712622712
transform 1 0 2204 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4755
timestamp 1712622712
transform 1 0 2196 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4756
timestamp 1712622712
transform 1 0 2068 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4757
timestamp 1712622712
transform 1 0 2500 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4758
timestamp 1712622712
transform 1 0 2268 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4759
timestamp 1712622712
transform 1 0 2460 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4760
timestamp 1712622712
transform 1 0 2420 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4761
timestamp 1712622712
transform 1 0 2348 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4762
timestamp 1712622712
transform 1 0 2308 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4763
timestamp 1712622712
transform 1 0 2204 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4764
timestamp 1712622712
transform 1 0 2196 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4765
timestamp 1712622712
transform 1 0 2164 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4766
timestamp 1712622712
transform 1 0 2156 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4767
timestamp 1712622712
transform 1 0 2156 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4768
timestamp 1712622712
transform 1 0 2148 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4769
timestamp 1712622712
transform 1 0 2140 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4770
timestamp 1712622712
transform 1 0 2140 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4771
timestamp 1712622712
transform 1 0 2068 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4772
timestamp 1712622712
transform 1 0 2020 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4773
timestamp 1712622712
transform 1 0 2532 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4774
timestamp 1712622712
transform 1 0 2492 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4775
timestamp 1712622712
transform 1 0 2420 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4776
timestamp 1712622712
transform 1 0 2388 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1712622712
transform 1 0 2164 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4778
timestamp 1712622712
transform 1 0 2124 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4779
timestamp 1712622712
transform 1 0 1604 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4780
timestamp 1712622712
transform 1 0 2140 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1712622712
transform 1 0 1660 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4782
timestamp 1712622712
transform 1 0 2308 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4783
timestamp 1712622712
transform 1 0 2212 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4784
timestamp 1712622712
transform 1 0 1540 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4785
timestamp 1712622712
transform 1 0 1500 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1712622712
transform 1 0 1492 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1712622712
transform 1 0 1476 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4788
timestamp 1712622712
transform 1 0 1636 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4789
timestamp 1712622712
transform 1 0 1412 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1712622712
transform 1 0 3084 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4791
timestamp 1712622712
transform 1 0 2932 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4792
timestamp 1712622712
transform 1 0 2884 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4793
timestamp 1712622712
transform 1 0 2764 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4794
timestamp 1712622712
transform 1 0 2764 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4795
timestamp 1712622712
transform 1 0 2700 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1712622712
transform 1 0 2700 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4797
timestamp 1712622712
transform 1 0 2572 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4798
timestamp 1712622712
transform 1 0 1604 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4799
timestamp 1712622712
transform 1 0 2340 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4800
timestamp 1712622712
transform 1 0 2324 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4801
timestamp 1712622712
transform 1 0 2284 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4802
timestamp 1712622712
transform 1 0 2180 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4803
timestamp 1712622712
transform 1 0 2492 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4804
timestamp 1712622712
transform 1 0 2316 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4805
timestamp 1712622712
transform 1 0 2460 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4806
timestamp 1712622712
transform 1 0 2332 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4807
timestamp 1712622712
transform 1 0 2332 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4808
timestamp 1712622712
transform 1 0 2268 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4809
timestamp 1712622712
transform 1 0 2236 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4810
timestamp 1712622712
transform 1 0 2124 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4811
timestamp 1712622712
transform 1 0 2084 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4812
timestamp 1712622712
transform 1 0 2068 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4813
timestamp 1712622712
transform 1 0 2468 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4814
timestamp 1712622712
transform 1 0 2268 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1712622712
transform 1 0 2132 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4816
timestamp 1712622712
transform 1 0 2100 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1712622712
transform 1 0 2108 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4818
timestamp 1712622712
transform 1 0 2052 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4819
timestamp 1712622712
transform 1 0 2140 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4820
timestamp 1712622712
transform 1 0 2092 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4821
timestamp 1712622712
transform 1 0 2564 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4822
timestamp 1712622712
transform 1 0 2444 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1712622712
transform 1 0 2364 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4824
timestamp 1712622712
transform 1 0 2260 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1712622712
transform 1 0 2108 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4826
timestamp 1712622712
transform 1 0 1460 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4827
timestamp 1712622712
transform 1 0 1380 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4828
timestamp 1712622712
transform 1 0 2652 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4829
timestamp 1712622712
transform 1 0 1756 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1712622712
transform 1 0 1420 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1712622712
transform 1 0 2684 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4832
timestamp 1712622712
transform 1 0 2596 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4833
timestamp 1712622712
transform 1 0 2460 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4834
timestamp 1712622712
transform 1 0 2308 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4835
timestamp 1712622712
transform 1 0 2252 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4836
timestamp 1712622712
transform 1 0 1540 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1712622712
transform 1 0 1396 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4838
timestamp 1712622712
transform 1 0 2340 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4839
timestamp 1712622712
transform 1 0 2268 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4840
timestamp 1712622712
transform 1 0 2260 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4841
timestamp 1712622712
transform 1 0 2228 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4842
timestamp 1712622712
transform 1 0 2260 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4843
timestamp 1712622712
transform 1 0 2220 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4844
timestamp 1712622712
transform 1 0 2516 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4845
timestamp 1712622712
transform 1 0 2308 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4846
timestamp 1712622712
transform 1 0 2476 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4847
timestamp 1712622712
transform 1 0 2460 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4848
timestamp 1712622712
transform 1 0 2596 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4849
timestamp 1712622712
transform 1 0 2420 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4850
timestamp 1712622712
transform 1 0 2300 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4851
timestamp 1712622712
transform 1 0 2124 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4852
timestamp 1712622712
transform 1 0 2068 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4853
timestamp 1712622712
transform 1 0 1972 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4854
timestamp 1712622712
transform 1 0 2468 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4855
timestamp 1712622712
transform 1 0 2404 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1712622712
transform 1 0 2404 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4857
timestamp 1712622712
transform 1 0 2364 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4858
timestamp 1712622712
transform 1 0 2036 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4859
timestamp 1712622712
transform 1 0 1980 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4860
timestamp 1712622712
transform 1 0 2236 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4861
timestamp 1712622712
transform 1 0 2220 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4862
timestamp 1712622712
transform 1 0 2500 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4863
timestamp 1712622712
transform 1 0 2468 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1712622712
transform 1 0 2460 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4865
timestamp 1712622712
transform 1 0 2388 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4866
timestamp 1712622712
transform 1 0 2388 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4867
timestamp 1712622712
transform 1 0 2308 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4868
timestamp 1712622712
transform 1 0 2612 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4869
timestamp 1712622712
transform 1 0 1828 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4870
timestamp 1712622712
transform 1 0 1716 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4871
timestamp 1712622712
transform 1 0 1804 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4872
timestamp 1712622712
transform 1 0 1716 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4873
timestamp 1712622712
transform 1 0 1796 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4874
timestamp 1712622712
transform 1 0 1764 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4875
timestamp 1712622712
transform 1 0 1852 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4876
timestamp 1712622712
transform 1 0 1804 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4877
timestamp 1712622712
transform 1 0 1804 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4878
timestamp 1712622712
transform 1 0 1788 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4879
timestamp 1712622712
transform 1 0 1700 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4880
timestamp 1712622712
transform 1 0 1700 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4881
timestamp 1712622712
transform 1 0 1868 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4882
timestamp 1712622712
transform 1 0 1852 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4883
timestamp 1712622712
transform 1 0 1844 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4884
timestamp 1712622712
transform 1 0 1828 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4885
timestamp 1712622712
transform 1 0 1820 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4886
timestamp 1712622712
transform 1 0 1932 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4887
timestamp 1712622712
transform 1 0 1716 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4888
timestamp 1712622712
transform 1 0 1852 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4889
timestamp 1712622712
transform 1 0 1812 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4890
timestamp 1712622712
transform 1 0 1884 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4891
timestamp 1712622712
transform 1 0 1852 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4892
timestamp 1712622712
transform 1 0 3004 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4893
timestamp 1712622712
transform 1 0 2868 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4894
timestamp 1712622712
transform 1 0 2868 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4895
timestamp 1712622712
transform 1 0 2828 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4896
timestamp 1712622712
transform 1 0 2796 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4897
timestamp 1712622712
transform 1 0 2764 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4898
timestamp 1712622712
transform 1 0 2692 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4899
timestamp 1712622712
transform 1 0 2692 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4900
timestamp 1712622712
transform 1 0 2532 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4901
timestamp 1712622712
transform 1 0 2532 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4902
timestamp 1712622712
transform 1 0 2084 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4903
timestamp 1712622712
transform 1 0 1900 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4904
timestamp 1712622712
transform 1 0 1724 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4905
timestamp 1712622712
transform 1 0 2932 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4906
timestamp 1712622712
transform 1 0 2708 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4907
timestamp 1712622712
transform 1 0 2708 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4908
timestamp 1712622712
transform 1 0 2692 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4909
timestamp 1712622712
transform 1 0 2684 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4910
timestamp 1712622712
transform 1 0 2668 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4911
timestamp 1712622712
transform 1 0 2524 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1712622712
transform 1 0 2524 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4913
timestamp 1712622712
transform 1 0 1988 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4914
timestamp 1712622712
transform 1 0 1772 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4915
timestamp 1712622712
transform 1 0 1724 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4916
timestamp 1712622712
transform 1 0 1444 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4917
timestamp 1712622712
transform 1 0 1348 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4918
timestamp 1712622712
transform 1 0 2132 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4919
timestamp 1712622712
transform 1 0 2036 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4920
timestamp 1712622712
transform 1 0 1964 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4921
timestamp 1712622712
transform 1 0 1924 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1712622712
transform 1 0 2028 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4923
timestamp 1712622712
transform 1 0 1972 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4924
timestamp 1712622712
transform 1 0 1988 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4925
timestamp 1712622712
transform 1 0 1932 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4926
timestamp 1712622712
transform 1 0 2364 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4927
timestamp 1712622712
transform 1 0 2260 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4928
timestamp 1712622712
transform 1 0 2260 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4929
timestamp 1712622712
transform 1 0 2188 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4930
timestamp 1712622712
transform 1 0 2292 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4931
timestamp 1712622712
transform 1 0 2188 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4932
timestamp 1712622712
transform 1 0 2036 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4933
timestamp 1712622712
transform 1 0 1988 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4934
timestamp 1712622712
transform 1 0 2052 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4935
timestamp 1712622712
transform 1 0 1964 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4936
timestamp 1712622712
transform 1 0 2172 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4937
timestamp 1712622712
transform 1 0 2068 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1712622712
transform 1 0 2220 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4939
timestamp 1712622712
transform 1 0 2148 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4940
timestamp 1712622712
transform 1 0 2284 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4941
timestamp 1712622712
transform 1 0 2268 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4942
timestamp 1712622712
transform 1 0 2268 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4943
timestamp 1712622712
transform 1 0 2236 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1712622712
transform 1 0 2436 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4945
timestamp 1712622712
transform 1 0 2236 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1712622712
transform 1 0 3036 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4947
timestamp 1712622712
transform 1 0 2988 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4948
timestamp 1712622712
transform 1 0 2764 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4949
timestamp 1712622712
transform 1 0 2484 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4950
timestamp 1712622712
transform 1 0 2452 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4951
timestamp 1712622712
transform 1 0 2452 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4952
timestamp 1712622712
transform 1 0 2452 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4953
timestamp 1712622712
transform 1 0 2428 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4954
timestamp 1712622712
transform 1 0 2396 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4955
timestamp 1712622712
transform 1 0 2212 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4956
timestamp 1712622712
transform 1 0 2132 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4957
timestamp 1712622712
transform 1 0 2388 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4958
timestamp 1712622712
transform 1 0 2228 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1712622712
transform 1 0 2276 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4960
timestamp 1712622712
transform 1 0 2180 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4961
timestamp 1712622712
transform 1 0 2332 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4962
timestamp 1712622712
transform 1 0 2284 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4963
timestamp 1712622712
transform 1 0 2308 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4964
timestamp 1712622712
transform 1 0 2164 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4965
timestamp 1712622712
transform 1 0 2468 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4966
timestamp 1712622712
transform 1 0 2276 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4967
timestamp 1712622712
transform 1 0 2332 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4968
timestamp 1712622712
transform 1 0 2308 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4969
timestamp 1712622712
transform 1 0 2364 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4970
timestamp 1712622712
transform 1 0 2356 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4971
timestamp 1712622712
transform 1 0 2348 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4972
timestamp 1712622712
transform 1 0 2284 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4973
timestamp 1712622712
transform 1 0 2420 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4974
timestamp 1712622712
transform 1 0 2372 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1712622712
transform 1 0 2348 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4976
timestamp 1712622712
transform 1 0 2348 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4977
timestamp 1712622712
transform 1 0 2340 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4978
timestamp 1712622712
transform 1 0 2244 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4979
timestamp 1712622712
transform 1 0 2460 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4980
timestamp 1712622712
transform 1 0 2308 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4981
timestamp 1712622712
transform 1 0 2444 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1712622712
transform 1 0 2348 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1712622712
transform 1 0 2500 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4984
timestamp 1712622712
transform 1 0 2436 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4985
timestamp 1712622712
transform 1 0 2924 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4986
timestamp 1712622712
transform 1 0 2796 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4987
timestamp 1712622712
transform 1 0 2564 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4988
timestamp 1712622712
transform 1 0 2460 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4989
timestamp 1712622712
transform 1 0 2412 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4990
timestamp 1712622712
transform 1 0 2404 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4991
timestamp 1712622712
transform 1 0 2348 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4992
timestamp 1712622712
transform 1 0 2476 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4993
timestamp 1712622712
transform 1 0 2356 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4994
timestamp 1712622712
transform 1 0 2980 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4995
timestamp 1712622712
transform 1 0 2940 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4996
timestamp 1712622712
transform 1 0 2764 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4997
timestamp 1712622712
transform 1 0 2668 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4998
timestamp 1712622712
transform 1 0 2500 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4999
timestamp 1712622712
transform 1 0 2468 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5000
timestamp 1712622712
transform 1 0 2468 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5001
timestamp 1712622712
transform 1 0 2452 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5002
timestamp 1712622712
transform 1 0 2436 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5003
timestamp 1712622712
transform 1 0 2436 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5004
timestamp 1712622712
transform 1 0 2396 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5005
timestamp 1712622712
transform 1 0 2612 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5006
timestamp 1712622712
transform 1 0 2468 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5007
timestamp 1712622712
transform 1 0 2596 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5008
timestamp 1712622712
transform 1 0 2556 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5009
timestamp 1712622712
transform 1 0 2612 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5010
timestamp 1712622712
transform 1 0 2500 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5011
timestamp 1712622712
transform 1 0 2620 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5012
timestamp 1712622712
transform 1 0 2580 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5013
timestamp 1712622712
transform 1 0 2596 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5014
timestamp 1712622712
transform 1 0 2492 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5015
timestamp 1712622712
transform 1 0 2764 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_5016
timestamp 1712622712
transform 1 0 2764 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5017
timestamp 1712622712
transform 1 0 2740 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5018
timestamp 1712622712
transform 1 0 2724 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5019
timestamp 1712622712
transform 1 0 2724 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5020
timestamp 1712622712
transform 1 0 2644 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_5021
timestamp 1712622712
transform 1 0 2516 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5022
timestamp 1712622712
transform 1 0 2124 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_5023
timestamp 1712622712
transform 1 0 2668 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5024
timestamp 1712622712
transform 1 0 2564 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5025
timestamp 1712622712
transform 1 0 2684 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5026
timestamp 1712622712
transform 1 0 2644 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5027
timestamp 1712622712
transform 1 0 2620 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5028
timestamp 1712622712
transform 1 0 2572 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5029
timestamp 1712622712
transform 1 0 2724 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5030
timestamp 1712622712
transform 1 0 2668 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5031
timestamp 1712622712
transform 1 0 2892 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5032
timestamp 1712622712
transform 1 0 2852 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5033
timestamp 1712622712
transform 1 0 2780 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5034
timestamp 1712622712
transform 1 0 2716 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5035
timestamp 1712622712
transform 1 0 2684 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5036
timestamp 1712622712
transform 1 0 2116 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_5037
timestamp 1712622712
transform 1 0 2052 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_5038
timestamp 1712622712
transform 1 0 3308 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1712622712
transform 1 0 3164 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5040
timestamp 1712622712
transform 1 0 3116 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5041
timestamp 1712622712
transform 1 0 2612 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5042
timestamp 1712622712
transform 1 0 2684 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5043
timestamp 1712622712
transform 1 0 2468 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5044
timestamp 1712622712
transform 1 0 2012 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5045
timestamp 1712622712
transform 1 0 2012 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5046
timestamp 1712622712
transform 1 0 1948 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5047
timestamp 1712622712
transform 1 0 1908 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5048
timestamp 1712622712
transform 1 0 3228 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5049
timestamp 1712622712
transform 1 0 3180 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5050
timestamp 1712622712
transform 1 0 3284 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5051
timestamp 1712622712
transform 1 0 3212 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5052
timestamp 1712622712
transform 1 0 3212 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5053
timestamp 1712622712
transform 1 0 3180 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5054
timestamp 1712622712
transform 1 0 2692 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5055
timestamp 1712622712
transform 1 0 2652 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5056
timestamp 1712622712
transform 1 0 2764 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5057
timestamp 1712622712
transform 1 0 2692 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5058
timestamp 1712622712
transform 1 0 2740 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5059
timestamp 1712622712
transform 1 0 2668 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5060
timestamp 1712622712
transform 1 0 3004 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5061
timestamp 1712622712
transform 1 0 2868 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5062
timestamp 1712622712
transform 1 0 3060 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5063
timestamp 1712622712
transform 1 0 3020 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5064
timestamp 1712622712
transform 1 0 3060 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5065
timestamp 1712622712
transform 1 0 3020 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5066
timestamp 1712622712
transform 1 0 3020 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5067
timestamp 1712622712
transform 1 0 2980 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5068
timestamp 1712622712
transform 1 0 3236 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5069
timestamp 1712622712
transform 1 0 3140 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5070
timestamp 1712622712
transform 1 0 3124 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5071
timestamp 1712622712
transform 1 0 2996 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5072
timestamp 1712622712
transform 1 0 3060 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5073
timestamp 1712622712
transform 1 0 3044 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5074
timestamp 1712622712
transform 1 0 3060 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5075
timestamp 1712622712
transform 1 0 3012 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5076
timestamp 1712622712
transform 1 0 2996 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5077
timestamp 1712622712
transform 1 0 2924 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5078
timestamp 1712622712
transform 1 0 2908 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5079
timestamp 1712622712
transform 1 0 3116 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5080
timestamp 1712622712
transform 1 0 3044 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5081
timestamp 1712622712
transform 1 0 3060 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5082
timestamp 1712622712
transform 1 0 2820 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5083
timestamp 1712622712
transform 1 0 3116 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5084
timestamp 1712622712
transform 1 0 2972 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5085
timestamp 1712622712
transform 1 0 3060 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5086
timestamp 1712622712
transform 1 0 3060 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5087
timestamp 1712622712
transform 1 0 3020 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5088
timestamp 1712622712
transform 1 0 2996 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5089
timestamp 1712622712
transform 1 0 3028 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5090
timestamp 1712622712
transform 1 0 2884 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5091
timestamp 1712622712
transform 1 0 2988 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5092
timestamp 1712622712
transform 1 0 2932 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5093
timestamp 1712622712
transform 1 0 2884 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5094
timestamp 1712622712
transform 1 0 3060 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_5095
timestamp 1712622712
transform 1 0 3012 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_5096
timestamp 1712622712
transform 1 0 3268 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5097
timestamp 1712622712
transform 1 0 3268 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5098
timestamp 1712622712
transform 1 0 3212 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1712622712
transform 1 0 3204 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5100
timestamp 1712622712
transform 1 0 3204 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5101
timestamp 1712622712
transform 1 0 3180 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5102
timestamp 1712622712
transform 1 0 3180 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5103
timestamp 1712622712
transform 1 0 3156 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5104
timestamp 1712622712
transform 1 0 3148 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5105
timestamp 1712622712
transform 1 0 2980 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5106
timestamp 1712622712
transform 1 0 2924 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5107
timestamp 1712622712
transform 1 0 2836 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5108
timestamp 1712622712
transform 1 0 3060 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5109
timestamp 1712622712
transform 1 0 3044 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5110
timestamp 1712622712
transform 1 0 3076 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5111
timestamp 1712622712
transform 1 0 3044 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5112
timestamp 1712622712
transform 1 0 3172 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5113
timestamp 1712622712
transform 1 0 3036 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5114
timestamp 1712622712
transform 1 0 3116 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5115
timestamp 1712622712
transform 1 0 3060 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5116
timestamp 1712622712
transform 1 0 3204 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5117
timestamp 1712622712
transform 1 0 3132 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5118
timestamp 1712622712
transform 1 0 2692 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5119
timestamp 1712622712
transform 1 0 2660 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5120
timestamp 1712622712
transform 1 0 2612 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5121
timestamp 1712622712
transform 1 0 2564 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5122
timestamp 1712622712
transform 1 0 2508 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5123
timestamp 1712622712
transform 1 0 2500 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5124
timestamp 1712622712
transform 1 0 2492 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5125
timestamp 1712622712
transform 1 0 2484 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5126
timestamp 1712622712
transform 1 0 3100 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5127
timestamp 1712622712
transform 1 0 3044 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5128
timestamp 1712622712
transform 1 0 3004 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5129
timestamp 1712622712
transform 1 0 3004 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5130
timestamp 1712622712
transform 1 0 3084 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5131
timestamp 1712622712
transform 1 0 3044 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5132
timestamp 1712622712
transform 1 0 2972 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5133
timestamp 1712622712
transform 1 0 3044 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5134
timestamp 1712622712
transform 1 0 2748 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5135
timestamp 1712622712
transform 1 0 2988 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5136
timestamp 1712622712
transform 1 0 2908 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5137
timestamp 1712622712
transform 1 0 3108 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5138
timestamp 1712622712
transform 1 0 3100 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5139
timestamp 1712622712
transform 1 0 3076 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5140
timestamp 1712622712
transform 1 0 2924 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5141
timestamp 1712622712
transform 1 0 3188 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5142
timestamp 1712622712
transform 1 0 2988 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5143
timestamp 1712622712
transform 1 0 2988 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5144
timestamp 1712622712
transform 1 0 2948 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5145
timestamp 1712622712
transform 1 0 2580 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_5146
timestamp 1712622712
transform 1 0 2516 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_5147
timestamp 1712622712
transform 1 0 3092 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5148
timestamp 1712622712
transform 1 0 2964 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5149
timestamp 1712622712
transform 1 0 2972 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5150
timestamp 1712622712
transform 1 0 2924 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5151
timestamp 1712622712
transform 1 0 2876 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5152
timestamp 1712622712
transform 1 0 2812 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5153
timestamp 1712622712
transform 1 0 3068 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5154
timestamp 1712622712
transform 1 0 2916 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5155
timestamp 1712622712
transform 1 0 3100 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5156
timestamp 1712622712
transform 1 0 3044 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5157
timestamp 1712622712
transform 1 0 2636 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1712622712
transform 1 0 2564 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5159
timestamp 1712622712
transform 1 0 2988 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5160
timestamp 1712622712
transform 1 0 2940 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5161
timestamp 1712622712
transform 1 0 3100 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5162
timestamp 1712622712
transform 1 0 2932 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5163
timestamp 1712622712
transform 1 0 2836 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5164
timestamp 1712622712
transform 1 0 3228 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5165
timestamp 1712622712
transform 1 0 3132 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5166
timestamp 1712622712
transform 1 0 2892 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5167
timestamp 1712622712
transform 1 0 2964 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5168
timestamp 1712622712
transform 1 0 2748 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5169
timestamp 1712622712
transform 1 0 2908 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5170
timestamp 1712622712
transform 1 0 2836 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5171
timestamp 1712622712
transform 1 0 2868 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5172
timestamp 1712622712
transform 1 0 2828 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5173
timestamp 1712622712
transform 1 0 2876 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5174
timestamp 1712622712
transform 1 0 2852 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5175
timestamp 1712622712
transform 1 0 2740 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5176
timestamp 1712622712
transform 1 0 2660 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5177
timestamp 1712622712
transform 1 0 2876 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1712622712
transform 1 0 2804 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5179
timestamp 1712622712
transform 1 0 2796 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5180
timestamp 1712622712
transform 1 0 2756 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5181
timestamp 1712622712
transform 1 0 2908 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5182
timestamp 1712622712
transform 1 0 2804 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5183
timestamp 1712622712
transform 1 0 2980 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5184
timestamp 1712622712
transform 1 0 2892 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5185
timestamp 1712622712
transform 1 0 3228 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5186
timestamp 1712622712
transform 1 0 3188 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5187
timestamp 1712622712
transform 1 0 2628 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5188
timestamp 1712622712
transform 1 0 2500 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_5189
timestamp 1712622712
transform 1 0 2916 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5190
timestamp 1712622712
transform 1 0 2804 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1712622712
transform 1 0 2812 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5192
timestamp 1712622712
transform 1 0 2700 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5193
timestamp 1712622712
transform 1 0 2828 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5194
timestamp 1712622712
transform 1 0 2812 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5195
timestamp 1712622712
transform 1 0 2804 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5196
timestamp 1712622712
transform 1 0 2772 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5197
timestamp 1712622712
transform 1 0 2724 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5198
timestamp 1712622712
transform 1 0 2868 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5199
timestamp 1712622712
transform 1 0 2836 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5200
timestamp 1712622712
transform 1 0 2804 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5201
timestamp 1712622712
transform 1 0 2756 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5202
timestamp 1712622712
transform 1 0 2668 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5203
timestamp 1712622712
transform 1 0 2516 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5204
timestamp 1712622712
transform 1 0 3220 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5205
timestamp 1712622712
transform 1 0 3188 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5206
timestamp 1712622712
transform 1 0 3380 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_5207
timestamp 1712622712
transform 1 0 3332 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_5208
timestamp 1712622712
transform 1 0 3180 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_5209
timestamp 1712622712
transform 1 0 3092 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_5210
timestamp 1712622712
transform 1 0 3332 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5211
timestamp 1712622712
transform 1 0 3196 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5212
timestamp 1712622712
transform 1 0 3436 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5213
timestamp 1712622712
transform 1 0 3324 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5214
timestamp 1712622712
transform 1 0 3068 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5215
timestamp 1712622712
transform 1 0 2892 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5216
timestamp 1712622712
transform 1 0 3292 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5217
timestamp 1712622712
transform 1 0 3244 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5218
timestamp 1712622712
transform 1 0 3348 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5219
timestamp 1712622712
transform 1 0 3300 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5220
timestamp 1712622712
transform 1 0 3196 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5221
timestamp 1712622712
transform 1 0 3196 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5222
timestamp 1712622712
transform 1 0 3340 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5223
timestamp 1712622712
transform 1 0 3340 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5224
timestamp 1712622712
transform 1 0 3324 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5225
timestamp 1712622712
transform 1 0 3284 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5226
timestamp 1712622712
transform 1 0 3396 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5227
timestamp 1712622712
transform 1 0 3372 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5228
timestamp 1712622712
transform 1 0 3412 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5229
timestamp 1712622712
transform 1 0 3388 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5230
timestamp 1712622712
transform 1 0 3364 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5231
timestamp 1712622712
transform 1 0 3348 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5232
timestamp 1712622712
transform 1 0 3300 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5233
timestamp 1712622712
transform 1 0 3044 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5234
timestamp 1712622712
transform 1 0 2964 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5235
timestamp 1712622712
transform 1 0 2932 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5236
timestamp 1712622712
transform 1 0 3404 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_5237
timestamp 1712622712
transform 1 0 3260 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5238
timestamp 1712622712
transform 1 0 3100 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5239
timestamp 1712622712
transform 1 0 2996 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5240
timestamp 1712622712
transform 1 0 2940 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5241
timestamp 1712622712
transform 1 0 3316 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5242
timestamp 1712622712
transform 1 0 3244 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5243
timestamp 1712622712
transform 1 0 3156 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5244
timestamp 1712622712
transform 1 0 3364 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5245
timestamp 1712622712
transform 1 0 3308 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5246
timestamp 1712622712
transform 1 0 3284 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5247
timestamp 1712622712
transform 1 0 3380 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5248
timestamp 1712622712
transform 1 0 3300 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5249
timestamp 1712622712
transform 1 0 3356 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5250
timestamp 1712622712
transform 1 0 3260 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5251
timestamp 1712622712
transform 1 0 3324 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_5252
timestamp 1712622712
transform 1 0 3292 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_5253
timestamp 1712622712
transform 1 0 3404 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5254
timestamp 1712622712
transform 1 0 3356 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5255
timestamp 1712622712
transform 1 0 3380 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5256
timestamp 1712622712
transform 1 0 3348 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5257
timestamp 1712622712
transform 1 0 3292 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5258
timestamp 1712622712
transform 1 0 3228 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5259
timestamp 1712622712
transform 1 0 3188 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5260
timestamp 1712622712
transform 1 0 3132 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5261
timestamp 1712622712
transform 1 0 3188 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1712622712
transform 1 0 3124 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5263
timestamp 1712622712
transform 1 0 3268 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5264
timestamp 1712622712
transform 1 0 3156 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5265
timestamp 1712622712
transform 1 0 3196 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5266
timestamp 1712622712
transform 1 0 3060 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5267
timestamp 1712622712
transform 1 0 3076 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5268
timestamp 1712622712
transform 1 0 2988 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5269
timestamp 1712622712
transform 1 0 2732 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5270
timestamp 1712622712
transform 1 0 2580 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5271
timestamp 1712622712
transform 1 0 1996 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1712622712
transform 1 0 1956 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5273
timestamp 1712622712
transform 1 0 2308 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5274
timestamp 1712622712
transform 1 0 2268 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5275
timestamp 1712622712
transform 1 0 1836 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5276
timestamp 1712622712
transform 1 0 1804 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1712622712
transform 1 0 1940 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5278
timestamp 1712622712
transform 1 0 1836 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5279
timestamp 1712622712
transform 1 0 1148 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1712622712
transform 1 0 1052 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1712622712
transform 1 0 356 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5282
timestamp 1712622712
transform 1 0 292 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5283
timestamp 1712622712
transform 1 0 452 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5284
timestamp 1712622712
transform 1 0 364 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1712622712
transform 1 0 468 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1712622712
transform 1 0 428 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1712622712
transform 1 0 908 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_5288
timestamp 1712622712
transform 1 0 844 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_5289
timestamp 1712622712
transform 1 0 3036 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5290
timestamp 1712622712
transform 1 0 2948 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5291
timestamp 1712622712
transform 1 0 3076 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5292
timestamp 1712622712
transform 1 0 3052 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5293
timestamp 1712622712
transform 1 0 3164 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5294
timestamp 1712622712
transform 1 0 2972 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1712622712
transform 1 0 3044 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5296
timestamp 1712622712
transform 1 0 2956 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5297
timestamp 1712622712
transform 1 0 2908 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1712622712
transform 1 0 2828 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1712622712
transform 1 0 2988 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1712622712
transform 1 0 2876 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1712622712
transform 1 0 2820 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5302
timestamp 1712622712
transform 1 0 2676 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1712622712
transform 1 0 2660 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5304
timestamp 1712622712
transform 1 0 2612 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5305
timestamp 1712622712
transform 1 0 2276 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5306
timestamp 1712622712
transform 1 0 2172 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5307
timestamp 1712622712
transform 1 0 2124 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5308
timestamp 1712622712
transform 1 0 1124 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5309
timestamp 1712622712
transform 1 0 2452 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5310
timestamp 1712622712
transform 1 0 2388 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5311
timestamp 1712622712
transform 1 0 2180 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5312
timestamp 1712622712
transform 1 0 1764 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5313
timestamp 1712622712
transform 1 0 1652 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5314
timestamp 1712622712
transform 1 0 1324 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5315
timestamp 1712622712
transform 1 0 1228 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5316
timestamp 1712622712
transform 1 0 1076 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5317
timestamp 1712622712
transform 1 0 996 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5318
timestamp 1712622712
transform 1 0 1076 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5319
timestamp 1712622712
transform 1 0 932 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5320
timestamp 1712622712
transform 1 0 924 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5321
timestamp 1712622712
transform 1 0 868 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5322
timestamp 1712622712
transform 1 0 1148 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5323
timestamp 1712622712
transform 1 0 948 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5324
timestamp 1712622712
transform 1 0 1164 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5325
timestamp 1712622712
transform 1 0 1132 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1712622712
transform 1 0 908 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_5327
timestamp 1712622712
transform 1 0 908 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5328
timestamp 1712622712
transform 1 0 788 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1712622712
transform 1 0 564 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5330
timestamp 1712622712
transform 1 0 2092 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5331
timestamp 1712622712
transform 1 0 1980 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5332
timestamp 1712622712
transform 1 0 1860 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5333
timestamp 1712622712
transform 1 0 1756 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5334
timestamp 1712622712
transform 1 0 2100 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5335
timestamp 1712622712
transform 1 0 1988 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5336
timestamp 1712622712
transform 1 0 1940 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5337
timestamp 1712622712
transform 1 0 1756 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5338
timestamp 1712622712
transform 1 0 1564 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5339
timestamp 1712622712
transform 1 0 1564 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5340
timestamp 1712622712
transform 1 0 1484 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5341
timestamp 1712622712
transform 1 0 2436 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5342
timestamp 1712622712
transform 1 0 2412 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5343
timestamp 1712622712
transform 1 0 2084 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5344
timestamp 1712622712
transform 1 0 2068 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5345
timestamp 1712622712
transform 1 0 1956 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5346
timestamp 1712622712
transform 1 0 3156 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5347
timestamp 1712622712
transform 1 0 3084 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5348
timestamp 1712622712
transform 1 0 2836 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5349
timestamp 1712622712
transform 1 0 2828 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5350
timestamp 1712622712
transform 1 0 2652 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5351
timestamp 1712622712
transform 1 0 2436 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5352
timestamp 1712622712
transform 1 0 2372 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5353
timestamp 1712622712
transform 1 0 2868 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5354
timestamp 1712622712
transform 1 0 2828 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5355
timestamp 1712622712
transform 1 0 2676 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5356
timestamp 1712622712
transform 1 0 2676 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5357
timestamp 1712622712
transform 1 0 956 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5358
timestamp 1712622712
transform 1 0 860 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5359
timestamp 1712622712
transform 1 0 564 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5360
timestamp 1712622712
transform 1 0 524 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5361
timestamp 1712622712
transform 1 0 524 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5362
timestamp 1712622712
transform 1 0 436 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5363
timestamp 1712622712
transform 1 0 404 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5364
timestamp 1712622712
transform 1 0 404 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5365
timestamp 1712622712
transform 1 0 388 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5366
timestamp 1712622712
transform 1 0 372 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5367
timestamp 1712622712
transform 1 0 220 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5368
timestamp 1712622712
transform 1 0 2940 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5369
timestamp 1712622712
transform 1 0 2852 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5370
timestamp 1712622712
transform 1 0 2780 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5371
timestamp 1712622712
transform 1 0 2740 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5372
timestamp 1712622712
transform 1 0 2724 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5373
timestamp 1712622712
transform 1 0 2556 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5374
timestamp 1712622712
transform 1 0 3036 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5375
timestamp 1712622712
transform 1 0 2972 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5376
timestamp 1712622712
transform 1 0 3020 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5377
timestamp 1712622712
transform 1 0 2996 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5378
timestamp 1712622712
transform 1 0 2556 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5379
timestamp 1712622712
transform 1 0 2524 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5380
timestamp 1712622712
transform 1 0 2596 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5381
timestamp 1712622712
transform 1 0 2580 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5382
timestamp 1712622712
transform 1 0 2548 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5383
timestamp 1712622712
transform 1 0 2508 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5384
timestamp 1712622712
transform 1 0 2508 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1712622712
transform 1 0 2508 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5386
timestamp 1712622712
transform 1 0 2460 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5387
timestamp 1712622712
transform 1 0 2892 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5388
timestamp 1712622712
transform 1 0 2788 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5389
timestamp 1712622712
transform 1 0 2740 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5390
timestamp 1712622712
transform 1 0 2764 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5391
timestamp 1712622712
transform 1 0 2644 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5392
timestamp 1712622712
transform 1 0 2628 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5393
timestamp 1712622712
transform 1 0 2572 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5394
timestamp 1712622712
transform 1 0 2468 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5395
timestamp 1712622712
transform 1 0 2204 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5396
timestamp 1712622712
transform 1 0 2772 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5397
timestamp 1712622712
transform 1 0 2668 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5398
timestamp 1712622712
transform 1 0 2684 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5399
timestamp 1712622712
transform 1 0 2620 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5400
timestamp 1712622712
transform 1 0 2188 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5401
timestamp 1712622712
transform 1 0 2116 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5402
timestamp 1712622712
transform 1 0 2012 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5403
timestamp 1712622712
transform 1 0 2372 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5404
timestamp 1712622712
transform 1 0 2332 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5405
timestamp 1712622712
transform 1 0 2324 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5406
timestamp 1712622712
transform 1 0 2212 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5407
timestamp 1712622712
transform 1 0 2036 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5408
timestamp 1712622712
transform 1 0 2412 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5409
timestamp 1712622712
transform 1 0 2380 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5410
timestamp 1712622712
transform 1 0 2260 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5411
timestamp 1712622712
transform 1 0 2068 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5412
timestamp 1712622712
transform 1 0 2004 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5413
timestamp 1712622712
transform 1 0 2300 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5414
timestamp 1712622712
transform 1 0 2132 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5415
timestamp 1712622712
transform 1 0 2036 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5416
timestamp 1712622712
transform 1 0 1900 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5417
timestamp 1712622712
transform 1 0 2316 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5418
timestamp 1712622712
transform 1 0 2076 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5419
timestamp 1712622712
transform 1 0 2356 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5420
timestamp 1712622712
transform 1 0 2308 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5421
timestamp 1712622712
transform 1 0 2276 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5422
timestamp 1712622712
transform 1 0 2172 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5423
timestamp 1712622712
transform 1 0 1980 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5424
timestamp 1712622712
transform 1 0 2340 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_5425
timestamp 1712622712
transform 1 0 2292 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_5426
timestamp 1712622712
transform 1 0 2356 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5427
timestamp 1712622712
transform 1 0 2284 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5428
timestamp 1712622712
transform 1 0 2324 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5429
timestamp 1712622712
transform 1 0 2196 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5430
timestamp 1712622712
transform 1 0 1916 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5431
timestamp 1712622712
transform 1 0 1788 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5432
timestamp 1712622712
transform 1 0 2028 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1712622712
transform 1 0 1844 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5434
timestamp 1712622712
transform 1 0 2268 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5435
timestamp 1712622712
transform 1 0 2036 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5436
timestamp 1712622712
transform 1 0 1940 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5437
timestamp 1712622712
transform 1 0 1980 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5438
timestamp 1712622712
transform 1 0 1900 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5439
timestamp 1712622712
transform 1 0 1860 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5440
timestamp 1712622712
transform 1 0 1756 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5441
timestamp 1712622712
transform 1 0 1724 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5442
timestamp 1712622712
transform 1 0 1692 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5443
timestamp 1712622712
transform 1 0 1908 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5444
timestamp 1712622712
transform 1 0 1804 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5445
timestamp 1712622712
transform 1 0 1916 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5446
timestamp 1712622712
transform 1 0 1828 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5447
timestamp 1712622712
transform 1 0 1908 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5448
timestamp 1712622712
transform 1 0 1852 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5449
timestamp 1712622712
transform 1 0 1788 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5450
timestamp 1712622712
transform 1 0 1732 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5451
timestamp 1712622712
transform 1 0 1652 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5452
timestamp 1712622712
transform 1 0 1948 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5453
timestamp 1712622712
transform 1 0 1884 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5454
timestamp 1712622712
transform 1 0 1772 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5455
timestamp 1712622712
transform 1 0 1700 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5456
timestamp 1712622712
transform 1 0 1716 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5457
timestamp 1712622712
transform 1 0 1628 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5458
timestamp 1712622712
transform 1 0 1716 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5459
timestamp 1712622712
transform 1 0 1660 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5460
timestamp 1712622712
transform 1 0 1892 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5461
timestamp 1712622712
transform 1 0 1820 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5462
timestamp 1712622712
transform 1 0 1772 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5463
timestamp 1712622712
transform 1 0 1812 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5464
timestamp 1712622712
transform 1 0 1652 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5465
timestamp 1712622712
transform 1 0 1580 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5466
timestamp 1712622712
transform 1 0 1572 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5467
timestamp 1712622712
transform 1 0 1556 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1712622712
transform 1 0 1548 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5469
timestamp 1712622712
transform 1 0 1748 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5470
timestamp 1712622712
transform 1 0 1644 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5471
timestamp 1712622712
transform 1 0 1540 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5472
timestamp 1712622712
transform 1 0 1436 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5473
timestamp 1712622712
transform 1 0 1676 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5474
timestamp 1712622712
transform 1 0 1468 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5475
timestamp 1712622712
transform 1 0 1452 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5476
timestamp 1712622712
transform 1 0 1420 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5477
timestamp 1712622712
transform 1 0 1420 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5478
timestamp 1712622712
transform 1 0 1276 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5479
timestamp 1712622712
transform 1 0 1244 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5480
timestamp 1712622712
transform 1 0 1644 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1712622712
transform 1 0 1548 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5482
timestamp 1712622712
transform 1 0 1444 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1712622712
transform 1 0 1348 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5484
timestamp 1712622712
transform 1 0 1572 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1712622712
transform 1 0 1452 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1712622712
transform 1 0 1308 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5487
timestamp 1712622712
transform 1 0 1252 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5488
timestamp 1712622712
transform 1 0 1588 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1712622712
transform 1 0 1332 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1712622712
transform 1 0 1268 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5491
timestamp 1712622712
transform 1 0 1188 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5492
timestamp 1712622712
transform 1 0 1532 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5493
timestamp 1712622712
transform 1 0 1276 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5494
timestamp 1712622712
transform 1 0 1596 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1712622712
transform 1 0 1476 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5496
timestamp 1712622712
transform 1 0 1364 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5497
timestamp 1712622712
transform 1 0 1252 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5498
timestamp 1712622712
transform 1 0 1148 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1712622712
transform 1 0 1036 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5500
timestamp 1712622712
transform 1 0 1324 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1712622712
transform 1 0 1132 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5502
timestamp 1712622712
transform 1 0 1356 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5503
timestamp 1712622712
transform 1 0 1332 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1712622712
transform 1 0 1460 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5505
timestamp 1712622712
transform 1 0 1340 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5506
timestamp 1712622712
transform 1 0 1228 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5507
timestamp 1712622712
transform 1 0 1124 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5508
timestamp 1712622712
transform 1 0 1012 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5509
timestamp 1712622712
transform 1 0 956 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1712622712
transform 1 0 260 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5511
timestamp 1712622712
transform 1 0 1212 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5512
timestamp 1712622712
transform 1 0 932 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5513
timestamp 1712622712
transform 1 0 548 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5514
timestamp 1712622712
transform 1 0 244 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5515
timestamp 1712622712
transform 1 0 1108 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5516
timestamp 1712622712
transform 1 0 548 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5517
timestamp 1712622712
transform 1 0 1140 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5518
timestamp 1712622712
transform 1 0 1116 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5519
timestamp 1712622712
transform 1 0 660 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5520
timestamp 1712622712
transform 1 0 292 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5521
timestamp 1712622712
transform 1 0 1028 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5522
timestamp 1712622712
transform 1 0 628 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5523
timestamp 1712622712
transform 1 0 964 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5524
timestamp 1712622712
transform 1 0 932 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5525
timestamp 1712622712
transform 1 0 1036 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5526
timestamp 1712622712
transform 1 0 844 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5527
timestamp 1712622712
transform 1 0 756 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5528
timestamp 1712622712
transform 1 0 1060 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5529
timestamp 1712622712
transform 1 0 900 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5530
timestamp 1712622712
transform 1 0 892 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5531
timestamp 1712622712
transform 1 0 580 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5532
timestamp 1712622712
transform 1 0 532 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5533
timestamp 1712622712
transform 1 0 420 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5534
timestamp 1712622712
transform 1 0 660 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5535
timestamp 1712622712
transform 1 0 524 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5536
timestamp 1712622712
transform 1 0 756 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5537
timestamp 1712622712
transform 1 0 660 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5538
timestamp 1712622712
transform 1 0 956 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5539
timestamp 1712622712
transform 1 0 900 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5540
timestamp 1712622712
transform 1 0 716 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5541
timestamp 1712622712
transform 1 0 716 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5542
timestamp 1712622712
transform 1 0 692 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5543
timestamp 1712622712
transform 1 0 644 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1712622712
transform 1 0 468 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5545
timestamp 1712622712
transform 1 0 452 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5546
timestamp 1712622712
transform 1 0 604 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5547
timestamp 1712622712
transform 1 0 452 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5548
timestamp 1712622712
transform 1 0 700 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5549
timestamp 1712622712
transform 1 0 628 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5550
timestamp 1712622712
transform 1 0 596 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5551
timestamp 1712622712
transform 1 0 452 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5552
timestamp 1712622712
transform 1 0 596 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5553
timestamp 1712622712
transform 1 0 492 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5554
timestamp 1712622712
transform 1 0 700 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5555
timestamp 1712622712
transform 1 0 636 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5556
timestamp 1712622712
transform 1 0 916 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5557
timestamp 1712622712
transform 1 0 836 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5558
timestamp 1712622712
transform 1 0 852 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5559
timestamp 1712622712
transform 1 0 788 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5560
timestamp 1712622712
transform 1 0 892 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5561
timestamp 1712622712
transform 1 0 796 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5562
timestamp 1712622712
transform 1 0 796 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5563
timestamp 1712622712
transform 1 0 708 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5564
timestamp 1712622712
transform 1 0 668 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5565
timestamp 1712622712
transform 1 0 620 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5566
timestamp 1712622712
transform 1 0 788 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5567
timestamp 1712622712
transform 1 0 596 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5568
timestamp 1712622712
transform 1 0 916 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5569
timestamp 1712622712
transform 1 0 892 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5570
timestamp 1712622712
transform 1 0 892 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5571
timestamp 1712622712
transform 1 0 780 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5572
timestamp 1712622712
transform 1 0 748 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5573
timestamp 1712622712
transform 1 0 668 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5574
timestamp 1712622712
transform 1 0 620 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5575
timestamp 1712622712
transform 1 0 740 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5576
timestamp 1712622712
transform 1 0 660 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5577
timestamp 1712622712
transform 1 0 740 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5578
timestamp 1712622712
transform 1 0 692 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5579
timestamp 1712622712
transform 1 0 884 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5580
timestamp 1712622712
transform 1 0 852 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5581
timestamp 1712622712
transform 1 0 804 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5582
timestamp 1712622712
transform 1 0 644 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5583
timestamp 1712622712
transform 1 0 924 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5584
timestamp 1712622712
transform 1 0 724 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5585
timestamp 1712622712
transform 1 0 940 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5586
timestamp 1712622712
transform 1 0 900 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5587
timestamp 1712622712
transform 1 0 820 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5588
timestamp 1712622712
transform 1 0 772 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5589
timestamp 1712622712
transform 1 0 1884 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5590
timestamp 1712622712
transform 1 0 1788 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5591
timestamp 1712622712
transform 1 0 1692 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5592
timestamp 1712622712
transform 1 0 1196 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5593
timestamp 1712622712
transform 1 0 1964 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5594
timestamp 1712622712
transform 1 0 1924 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5595
timestamp 1712622712
transform 1 0 3148 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_5596
timestamp 1712622712
transform 1 0 2948 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_5597
timestamp 1712622712
transform 1 0 2820 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_5598
timestamp 1712622712
transform 1 0 2772 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5599
timestamp 1712622712
transform 1 0 2396 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5600
timestamp 1712622712
transform 1 0 2332 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5601
timestamp 1712622712
transform 1 0 2180 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5602
timestamp 1712622712
transform 1 0 2084 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5603
timestamp 1712622712
transform 1 0 1820 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5604
timestamp 1712622712
transform 1 0 1132 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5605
timestamp 1712622712
transform 1 0 1132 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5606
timestamp 1712622712
transform 1 0 916 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5607
timestamp 1712622712
transform 1 0 692 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5608
timestamp 1712622712
transform 1 0 620 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5609
timestamp 1712622712
transform 1 0 492 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5610
timestamp 1712622712
transform 1 0 492 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5611
timestamp 1712622712
transform 1 0 468 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5612
timestamp 1712622712
transform 1 0 3244 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5613
timestamp 1712622712
transform 1 0 3156 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5614
timestamp 1712622712
transform 1 0 3124 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5615
timestamp 1712622712
transform 1 0 3156 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5616
timestamp 1712622712
transform 1 0 3092 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5617
timestamp 1712622712
transform 1 0 3092 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5618
timestamp 1712622712
transform 1 0 3028 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5619
timestamp 1712622712
transform 1 0 2908 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5620
timestamp 1712622712
transform 1 0 2620 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5621
timestamp 1712622712
transform 1 0 2412 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5622
timestamp 1712622712
transform 1 0 2340 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5623
timestamp 1712622712
transform 1 0 1988 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5624
timestamp 1712622712
transform 1 0 1988 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5625
timestamp 1712622712
transform 1 0 1860 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5626
timestamp 1712622712
transform 1 0 1684 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5627
timestamp 1712622712
transform 1 0 1524 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5628
timestamp 1712622712
transform 1 0 1252 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5629
timestamp 1712622712
transform 1 0 2508 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5630
timestamp 1712622712
transform 1 0 2372 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5631
timestamp 1712622712
transform 1 0 916 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5632
timestamp 1712622712
transform 1 0 852 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5633
timestamp 1712622712
transform 1 0 2052 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5634
timestamp 1712622712
transform 1 0 1884 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5635
timestamp 1712622712
transform 1 0 2724 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5636
timestamp 1712622712
transform 1 0 2652 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5637
timestamp 1712622712
transform 1 0 2844 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5638
timestamp 1712622712
transform 1 0 2764 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5639
timestamp 1712622712
transform 1 0 2636 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5640
timestamp 1712622712
transform 1 0 2556 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5641
timestamp 1712622712
transform 1 0 2452 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5642
timestamp 1712622712
transform 1 0 2420 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5643
timestamp 1712622712
transform 1 0 2092 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5644
timestamp 1712622712
transform 1 0 2020 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5645
timestamp 1712622712
transform 1 0 2348 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5646
timestamp 1712622712
transform 1 0 2308 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5647
timestamp 1712622712
transform 1 0 2116 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5648
timestamp 1712622712
transform 1 0 2036 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5649
timestamp 1712622712
transform 1 0 1812 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5650
timestamp 1712622712
transform 1 0 1740 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5651
timestamp 1712622712
transform 1 0 1956 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1712622712
transform 1 0 1892 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5653
timestamp 1712622712
transform 1 0 1660 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5654
timestamp 1712622712
transform 1 0 1580 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5655
timestamp 1712622712
transform 1 0 1604 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5656
timestamp 1712622712
transform 1 0 1532 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5657
timestamp 1712622712
transform 1 0 1412 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5658
timestamp 1712622712
transform 1 0 1340 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5659
timestamp 1712622712
transform 1 0 1172 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1712622712
transform 1 0 1076 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5661
timestamp 1712622712
transform 1 0 1180 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5662
timestamp 1712622712
transform 1 0 1116 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5663
timestamp 1712622712
transform 1 0 236 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5664
timestamp 1712622712
transform 1 0 140 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5665
timestamp 1712622712
transform 1 0 268 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5666
timestamp 1712622712
transform 1 0 140 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5667
timestamp 1712622712
transform 1 0 396 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5668
timestamp 1712622712
transform 1 0 260 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5669
timestamp 1712622712
transform 1 0 428 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5670
timestamp 1712622712
transform 1 0 324 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5671
timestamp 1712622712
transform 1 0 412 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5672
timestamp 1712622712
transform 1 0 308 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5673
timestamp 1712622712
transform 1 0 452 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5674
timestamp 1712622712
transform 1 0 364 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5675
timestamp 1712622712
transform 1 0 572 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5676
timestamp 1712622712
transform 1 0 524 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5677
timestamp 1712622712
transform 1 0 588 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5678
timestamp 1712622712
transform 1 0 484 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5679
timestamp 1712622712
transform 1 0 884 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5680
timestamp 1712622712
transform 1 0 820 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5681
timestamp 1712622712
transform 1 0 3356 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5682
timestamp 1712622712
transform 1 0 3308 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5683
timestamp 1712622712
transform 1 0 3196 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5684
timestamp 1712622712
transform 1 0 3060 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5685
timestamp 1712622712
transform 1 0 3164 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5686
timestamp 1712622712
transform 1 0 3068 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5687
timestamp 1712622712
transform 1 0 3436 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_5688
timestamp 1712622712
transform 1 0 3348 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1712622712
transform 1 0 3364 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5690
timestamp 1712622712
transform 1 0 3228 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5691
timestamp 1712622712
transform 1 0 3348 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1712622712
transform 1 0 3324 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1712622712
transform 1 0 3396 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1712622712
transform 1 0 3364 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5695
timestamp 1712622712
transform 1 0 3428 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5696
timestamp 1712622712
transform 1 0 3388 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5697
timestamp 1712622712
transform 1 0 3436 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5698
timestamp 1712622712
transform 1 0 3436 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5699
timestamp 1712622712
transform 1 0 3380 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5700
timestamp 1712622712
transform 1 0 3380 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5701
timestamp 1712622712
transform 1 0 3348 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5702
timestamp 1712622712
transform 1 0 3348 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1712622712
transform 1 0 3324 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5704
timestamp 1712622712
transform 1 0 3292 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5705
timestamp 1712622712
transform 1 0 3268 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5706
timestamp 1712622712
transform 1 0 3076 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5707
timestamp 1712622712
transform 1 0 3076 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1712622712
transform 1 0 2900 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5709
timestamp 1712622712
transform 1 0 2340 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5710
timestamp 1712622712
transform 1 0 2332 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1712622712
transform 1 0 2300 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5712
timestamp 1712622712
transform 1 0 2300 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5713
timestamp 1712622712
transform 1 0 2244 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1712622712
transform 1 0 2228 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5715
timestamp 1712622712
transform 1 0 3188 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1712622712
transform 1 0 2692 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5717
timestamp 1712622712
transform 1 0 2532 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5718
timestamp 1712622712
transform 1 0 2436 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5719
timestamp 1712622712
transform 1 0 2436 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5720
timestamp 1712622712
transform 1 0 2244 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5721
timestamp 1712622712
transform 1 0 2180 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5722
timestamp 1712622712
transform 1 0 2164 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5723
timestamp 1712622712
transform 1 0 2092 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5724
timestamp 1712622712
transform 1 0 1780 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1712622712
transform 1 0 1612 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5726
timestamp 1712622712
transform 1 0 1468 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5727
timestamp 1712622712
transform 1 0 980 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5728
timestamp 1712622712
transform 1 0 868 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5729
timestamp 1712622712
transform 1 0 2044 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5730
timestamp 1712622712
transform 1 0 2028 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5731
timestamp 1712622712
transform 1 0 2012 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_5732
timestamp 1712622712
transform 1 0 2004 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1712622712
transform 1 0 1980 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_5734
timestamp 1712622712
transform 1 0 1972 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5735
timestamp 1712622712
transform 1 0 1924 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_5736
timestamp 1712622712
transform 1 0 2204 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5737
timestamp 1712622712
transform 1 0 2156 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5738
timestamp 1712622712
transform 1 0 2116 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5739
timestamp 1712622712
transform 1 0 2108 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5740
timestamp 1712622712
transform 1 0 1708 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5741
timestamp 1712622712
transform 1 0 2364 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5742
timestamp 1712622712
transform 1 0 1756 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5743
timestamp 1712622712
transform 1 0 2500 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5744
timestamp 1712622712
transform 1 0 2420 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1712622712
transform 1 0 2268 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5746
timestamp 1712622712
transform 1 0 1932 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5747
timestamp 1712622712
transform 1 0 2612 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5748
timestamp 1712622712
transform 1 0 2492 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5749
timestamp 1712622712
transform 1 0 2492 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1712622712
transform 1 0 2444 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5751
timestamp 1712622712
transform 1 0 2244 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1712622712
transform 1 0 2244 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5753
timestamp 1712622712
transform 1 0 1892 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5754
timestamp 1712622712
transform 1 0 2772 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_5755
timestamp 1712622712
transform 1 0 2476 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5756
timestamp 1712622712
transform 1 0 2476 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_5757
timestamp 1712622712
transform 1 0 2420 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5758
timestamp 1712622712
transform 1 0 1316 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5759
timestamp 1712622712
transform 1 0 1164 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5760
timestamp 1712622712
transform 1 0 1164 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5761
timestamp 1712622712
transform 1 0 1004 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5762
timestamp 1712622712
transform 1 0 1004 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5763
timestamp 1712622712
transform 1 0 908 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5764
timestamp 1712622712
transform 1 0 876 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5765
timestamp 1712622712
transform 1 0 788 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5766
timestamp 1712622712
transform 1 0 2996 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5767
timestamp 1712622712
transform 1 0 2964 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5768
timestamp 1712622712
transform 1 0 2908 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5769
timestamp 1712622712
transform 1 0 2844 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5770
timestamp 1712622712
transform 1 0 2844 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5771
timestamp 1712622712
transform 1 0 844 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5772
timestamp 1712622712
transform 1 0 708 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5773
timestamp 1712622712
transform 1 0 980 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5774
timestamp 1712622712
transform 1 0 964 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5775
timestamp 1712622712
transform 1 0 948 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5776
timestamp 1712622712
transform 1 0 756 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5777
timestamp 1712622712
transform 1 0 652 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5778
timestamp 1712622712
transform 1 0 620 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5779
timestamp 1712622712
transform 1 0 860 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5780
timestamp 1712622712
transform 1 0 564 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5781
timestamp 1712622712
transform 1 0 564 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5782
timestamp 1712622712
transform 1 0 516 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5783
timestamp 1712622712
transform 1 0 468 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5784
timestamp 1712622712
transform 1 0 468 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5785
timestamp 1712622712
transform 1 0 676 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5786
timestamp 1712622712
transform 1 0 516 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5787
timestamp 1712622712
transform 1 0 428 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_5788
timestamp 1712622712
transform 1 0 420 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5789
timestamp 1712622712
transform 1 0 388 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_5790
timestamp 1712622712
transform 1 0 372 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5791
timestamp 1712622712
transform 1 0 572 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5792
timestamp 1712622712
transform 1 0 556 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5793
timestamp 1712622712
transform 1 0 548 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5794
timestamp 1712622712
transform 1 0 468 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5795
timestamp 1712622712
transform 1 0 356 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5796
timestamp 1712622712
transform 1 0 348 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5797
timestamp 1712622712
transform 1 0 324 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5798
timestamp 1712622712
transform 1 0 660 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5799
timestamp 1712622712
transform 1 0 540 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5800
timestamp 1712622712
transform 1 0 364 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5801
timestamp 1712622712
transform 1 0 364 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5802
timestamp 1712622712
transform 1 0 324 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5803
timestamp 1712622712
transform 1 0 276 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5804
timestamp 1712622712
transform 1 0 684 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5805
timestamp 1712622712
transform 1 0 676 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5806
timestamp 1712622712
transform 1 0 660 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5807
timestamp 1712622712
transform 1 0 588 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5808
timestamp 1712622712
transform 1 0 316 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5809
timestamp 1712622712
transform 1 0 316 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5810
timestamp 1712622712
transform 1 0 268 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5811
timestamp 1712622712
transform 1 0 252 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5812
timestamp 1712622712
transform 1 0 612 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5813
timestamp 1712622712
transform 1 0 580 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5814
timestamp 1712622712
transform 1 0 548 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5815
timestamp 1712622712
transform 1 0 420 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5816
timestamp 1712622712
transform 1 0 420 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5817
timestamp 1712622712
transform 1 0 92 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5818
timestamp 1712622712
transform 1 0 84 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5819
timestamp 1712622712
transform 1 0 804 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5820
timestamp 1712622712
transform 1 0 756 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5821
timestamp 1712622712
transform 1 0 732 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5822
timestamp 1712622712
transform 1 0 588 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5823
timestamp 1712622712
transform 1 0 556 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5824
timestamp 1712622712
transform 1 0 548 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5825
timestamp 1712622712
transform 1 0 340 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5826
timestamp 1712622712
transform 1 0 340 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5827
timestamp 1712622712
transform 1 0 324 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1712622712
transform 1 0 316 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5829
timestamp 1712622712
transform 1 0 172 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5830
timestamp 1712622712
transform 1 0 124 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5831
timestamp 1712622712
transform 1 0 92 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_5832
timestamp 1712622712
transform 1 0 868 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5833
timestamp 1712622712
transform 1 0 852 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5834
timestamp 1712622712
transform 1 0 828 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5835
timestamp 1712622712
transform 1 0 820 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5836
timestamp 1712622712
transform 1 0 780 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5837
timestamp 1712622712
transform 1 0 644 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5838
timestamp 1712622712
transform 1 0 636 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5839
timestamp 1712622712
transform 1 0 628 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5840
timestamp 1712622712
transform 1 0 532 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5841
timestamp 1712622712
transform 1 0 3076 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5842
timestamp 1712622712
transform 1 0 3044 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5843
timestamp 1712622712
transform 1 0 3044 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5844
timestamp 1712622712
transform 1 0 2988 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5845
timestamp 1712622712
transform 1 0 2908 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5846
timestamp 1712622712
transform 1 0 2900 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5847
timestamp 1712622712
transform 1 0 2868 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5848
timestamp 1712622712
transform 1 0 2868 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5849
timestamp 1712622712
transform 1 0 2644 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5850
timestamp 1712622712
transform 1 0 2644 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5851
timestamp 1712622712
transform 1 0 2540 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5852
timestamp 1712622712
transform 1 0 1220 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5853
timestamp 1712622712
transform 1 0 1052 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_5854
timestamp 1712622712
transform 1 0 1044 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5855
timestamp 1712622712
transform 1 0 1012 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5856
timestamp 1712622712
transform 1 0 972 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_5857
timestamp 1712622712
transform 1 0 964 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5858
timestamp 1712622712
transform 1 0 1292 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5859
timestamp 1712622712
transform 1 0 1284 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_5860
timestamp 1712622712
transform 1 0 1276 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1712622712
transform 1 0 1268 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1712622712
transform 1 0 1260 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1712622712
transform 1 0 1236 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5864
timestamp 1712622712
transform 1 0 1236 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5865
timestamp 1712622712
transform 1 0 1212 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_5866
timestamp 1712622712
transform 1 0 1204 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5867
timestamp 1712622712
transform 1 0 1204 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5868
timestamp 1712622712
transform 1 0 1204 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5869
timestamp 1712622712
transform 1 0 1204 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5870
timestamp 1712622712
transform 1 0 1156 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5871
timestamp 1712622712
transform 1 0 1156 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5872
timestamp 1712622712
transform 1 0 1108 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5873
timestamp 1712622712
transform 1 0 1108 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5874
timestamp 1712622712
transform 1 0 1460 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5875
timestamp 1712622712
transform 1 0 1404 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5876
timestamp 1712622712
transform 1 0 1404 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5877
timestamp 1712622712
transform 1 0 1300 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5878
timestamp 1712622712
transform 1 0 1292 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5879
timestamp 1712622712
transform 1 0 1284 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5880
timestamp 1712622712
transform 1 0 1252 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5881
timestamp 1712622712
transform 1 0 1252 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5882
timestamp 1712622712
transform 1 0 1252 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5883
timestamp 1712622712
transform 1 0 1204 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5884
timestamp 1712622712
transform 1 0 1204 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5885
timestamp 1712622712
transform 1 0 1204 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5886
timestamp 1712622712
transform 1 0 1516 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5887
timestamp 1712622712
transform 1 0 1516 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5888
timestamp 1712622712
transform 1 0 1516 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5889
timestamp 1712622712
transform 1 0 1484 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5890
timestamp 1712622712
transform 1 0 1460 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_5891
timestamp 1712622712
transform 1 0 1420 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5892
timestamp 1712622712
transform 1 0 1412 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5893
timestamp 1712622712
transform 1 0 1316 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5894
timestamp 1712622712
transform 1 0 1604 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5895
timestamp 1712622712
transform 1 0 1604 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5896
timestamp 1712622712
transform 1 0 1556 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5897
timestamp 1712622712
transform 1 0 1548 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5898
timestamp 1712622712
transform 1 0 1532 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5899
timestamp 1712622712
transform 1 0 1468 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5900
timestamp 1712622712
transform 1 0 1468 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_5901
timestamp 1712622712
transform 1 0 1796 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5902
timestamp 1712622712
transform 1 0 1780 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5903
timestamp 1712622712
transform 1 0 1780 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5904
timestamp 1712622712
transform 1 0 1780 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5905
timestamp 1712622712
transform 1 0 1708 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5906
timestamp 1712622712
transform 1 0 1684 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5907
timestamp 1712622712
transform 1 0 1660 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5908
timestamp 1712622712
transform 1 0 1660 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5909
timestamp 1712622712
transform 1 0 1964 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5910
timestamp 1712622712
transform 1 0 1940 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5911
timestamp 1712622712
transform 1 0 1892 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_5912
timestamp 1712622712
transform 1 0 1892 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5913
timestamp 1712622712
transform 1 0 1892 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5914
timestamp 1712622712
transform 1 0 1892 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5915
timestamp 1712622712
transform 1 0 1852 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_5916
timestamp 1712622712
transform 1 0 1852 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5917
timestamp 1712622712
transform 1 0 2148 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5918
timestamp 1712622712
transform 1 0 2100 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5919
timestamp 1712622712
transform 1 0 2052 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_5920
timestamp 1712622712
transform 1 0 2004 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_5921
timestamp 1712622712
transform 1 0 2284 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5922
timestamp 1712622712
transform 1 0 2252 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5923
timestamp 1712622712
transform 1 0 2236 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5924
timestamp 1712622712
transform 1 0 2196 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5925
timestamp 1712622712
transform 1 0 2180 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5926
timestamp 1712622712
transform 1 0 2172 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5927
timestamp 1712622712
transform 1 0 2068 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5928
timestamp 1712622712
transform 1 0 2852 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5929
timestamp 1712622712
transform 1 0 2732 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5930
timestamp 1712622712
transform 1 0 2708 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5931
timestamp 1712622712
transform 1 0 2684 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5932
timestamp 1712622712
transform 1 0 2580 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5933
timestamp 1712622712
transform 1 0 2580 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5934
timestamp 1712622712
transform 1 0 2492 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5935
timestamp 1712622712
transform 1 0 3340 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5936
timestamp 1712622712
transform 1 0 3084 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5937
timestamp 1712622712
transform 1 0 2468 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5938
timestamp 1712622712
transform 1 0 2388 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5939
timestamp 1712622712
transform 1 0 2300 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5940
timestamp 1712622712
transform 1 0 2564 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5941
timestamp 1712622712
transform 1 0 2548 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5942
timestamp 1712622712
transform 1 0 2484 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5943
timestamp 1712622712
transform 1 0 2348 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5944
timestamp 1712622712
transform 1 0 2780 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5945
timestamp 1712622712
transform 1 0 2596 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5946
timestamp 1712622712
transform 1 0 2588 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_5947
timestamp 1712622712
transform 1 0 2364 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_5948
timestamp 1712622712
transform 1 0 2364 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5949
timestamp 1712622712
transform 1 0 2300 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5950
timestamp 1712622712
transform 1 0 2388 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5951
timestamp 1712622712
transform 1 0 2340 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5952
timestamp 1712622712
transform 1 0 2204 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5953
timestamp 1712622712
transform 1 0 2556 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5954
timestamp 1712622712
transform 1 0 2452 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_5955
timestamp 1712622712
transform 1 0 2452 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5956
timestamp 1712622712
transform 1 0 2348 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_5957
timestamp 1712622712
transform 1 0 2620 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5958
timestamp 1712622712
transform 1 0 2580 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5959
timestamp 1712622712
transform 1 0 2500 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5960
timestamp 1712622712
transform 1 0 2412 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5961
timestamp 1712622712
transform 1 0 2588 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5962
timestamp 1712622712
transform 1 0 2564 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5963
timestamp 1712622712
transform 1 0 2436 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5964
timestamp 1712622712
transform 1 0 2428 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5965
timestamp 1712622712
transform 1 0 2340 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5966
timestamp 1712622712
transform 1 0 2252 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5967
timestamp 1712622712
transform 1 0 2468 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5968
timestamp 1712622712
transform 1 0 2220 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5969
timestamp 1712622712
transform 1 0 2020 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5970
timestamp 1712622712
transform 1 0 1956 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5971
timestamp 1712622712
transform 1 0 1852 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5972
timestamp 1712622712
transform 1 0 1844 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5973
timestamp 1712622712
transform 1 0 1628 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5974
timestamp 1712622712
transform 1 0 2300 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5975
timestamp 1712622712
transform 1 0 2236 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5976
timestamp 1712622712
transform 1 0 2236 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5977
timestamp 1712622712
transform 1 0 1972 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5978
timestamp 1712622712
transform 1 0 1908 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5979
timestamp 1712622712
transform 1 0 1868 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5980
timestamp 1712622712
transform 1 0 1868 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5981
timestamp 1712622712
transform 1 0 1556 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5982
timestamp 1712622712
transform 1 0 2164 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5983
timestamp 1712622712
transform 1 0 1940 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5984
timestamp 1712622712
transform 1 0 1780 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5985
timestamp 1712622712
transform 1 0 1772 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_5986
timestamp 1712622712
transform 1 0 1572 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5987
timestamp 1712622712
transform 1 0 2140 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5988
timestamp 1712622712
transform 1 0 2060 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5989
timestamp 1712622712
transform 1 0 1860 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5990
timestamp 1712622712
transform 1 0 1668 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5991
timestamp 1712622712
transform 1 0 1524 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5992
timestamp 1712622712
transform 1 0 1804 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_5993
timestamp 1712622712
transform 1 0 1804 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5994
timestamp 1712622712
transform 1 0 1684 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5995
timestamp 1712622712
transform 1 0 1652 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_5996
timestamp 1712622712
transform 1 0 1388 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_5997
timestamp 1712622712
transform 1 0 1948 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5998
timestamp 1712622712
transform 1 0 1868 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5999
timestamp 1712622712
transform 1 0 1796 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_6000
timestamp 1712622712
transform 1 0 1796 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6001
timestamp 1712622712
transform 1 0 1636 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_6002
timestamp 1712622712
transform 1 0 1636 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_6003
timestamp 1712622712
transform 1 0 1588 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_6004
timestamp 1712622712
transform 1 0 1396 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_6005
timestamp 1712622712
transform 1 0 1308 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_6006
timestamp 1712622712
transform 1 0 1724 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6007
timestamp 1712622712
transform 1 0 1620 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_6008
timestamp 1712622712
transform 1 0 1620 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6009
timestamp 1712622712
transform 1 0 1556 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_6010
timestamp 1712622712
transform 1 0 1428 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_6011
timestamp 1712622712
transform 1 0 1428 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6012
timestamp 1712622712
transform 1 0 1196 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6013
timestamp 1712622712
transform 1 0 1628 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6014
timestamp 1712622712
transform 1 0 1564 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6015
timestamp 1712622712
transform 1 0 1460 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_6016
timestamp 1712622712
transform 1 0 1420 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_6017
timestamp 1712622712
transform 1 0 1412 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_6018
timestamp 1712622712
transform 1 0 1412 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6019
timestamp 1712622712
transform 1 0 1036 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_6020
timestamp 1712622712
transform 1 0 1476 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_6021
timestamp 1712622712
transform 1 0 1300 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6022
timestamp 1712622712
transform 1 0 1188 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_6023
timestamp 1712622712
transform 1 0 1188 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_6024
timestamp 1712622712
transform 1 0 780 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_6025
timestamp 1712622712
transform 1 0 1380 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_6026
timestamp 1712622712
transform 1 0 1236 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_6027
timestamp 1712622712
transform 1 0 1108 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_6028
timestamp 1712622712
transform 1 0 1092 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_6029
timestamp 1712622712
transform 1 0 716 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_6030
timestamp 1712622712
transform 1 0 1308 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_6031
timestamp 1712622712
transform 1 0 1212 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_6032
timestamp 1712622712
transform 1 0 1084 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_6033
timestamp 1712622712
transform 1 0 1068 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_6034
timestamp 1712622712
transform 1 0 676 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_6035
timestamp 1712622712
transform 1 0 1204 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_6036
timestamp 1712622712
transform 1 0 1164 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6037
timestamp 1712622712
transform 1 0 1052 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6038
timestamp 1712622712
transform 1 0 1052 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_6039
timestamp 1712622712
transform 1 0 716 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_6040
timestamp 1712622712
transform 1 0 1340 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_6041
timestamp 1712622712
transform 1 0 1148 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6042
timestamp 1712622712
transform 1 0 1076 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6043
timestamp 1712622712
transform 1 0 1076 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_6044
timestamp 1712622712
transform 1 0 1076 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6045
timestamp 1712622712
transform 1 0 1044 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6046
timestamp 1712622712
transform 1 0 860 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6047
timestamp 1712622712
transform 1 0 860 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6048
timestamp 1712622712
transform 1 0 764 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6049
timestamp 1712622712
transform 1 0 1212 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6050
timestamp 1712622712
transform 1 0 988 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6051
timestamp 1712622712
transform 1 0 972 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6052
timestamp 1712622712
transform 1 0 964 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6053
timestamp 1712622712
transform 1 0 916 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6054
timestamp 1712622712
transform 1 0 772 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_6055
timestamp 1712622712
transform 1 0 700 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_6056
timestamp 1712622712
transform 1 0 1124 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6057
timestamp 1712622712
transform 1 0 836 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6058
timestamp 1712622712
transform 1 0 748 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6059
timestamp 1712622712
transform 1 0 652 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6060
timestamp 1712622712
transform 1 0 564 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6061
timestamp 1712622712
transform 1 0 1012 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6062
timestamp 1712622712
transform 1 0 812 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6063
timestamp 1712622712
transform 1 0 764 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6064
timestamp 1712622712
transform 1 0 732 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6065
timestamp 1712622712
transform 1 0 668 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6066
timestamp 1712622712
transform 1 0 748 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6067
timestamp 1712622712
transform 1 0 724 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_6068
timestamp 1712622712
transform 1 0 620 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_6069
timestamp 1712622712
transform 1 0 548 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6070
timestamp 1712622712
transform 1 0 524 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_6071
timestamp 1712622712
transform 1 0 500 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_6072
timestamp 1712622712
transform 1 0 684 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6073
timestamp 1712622712
transform 1 0 684 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6074
timestamp 1712622712
transform 1 0 580 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6075
timestamp 1712622712
transform 1 0 508 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6076
timestamp 1712622712
transform 1 0 508 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6077
timestamp 1712622712
transform 1 0 500 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6078
timestamp 1712622712
transform 1 0 628 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_6079
timestamp 1712622712
transform 1 0 596 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6080
timestamp 1712622712
transform 1 0 548 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6081
timestamp 1712622712
transform 1 0 532 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_6082
timestamp 1712622712
transform 1 0 492 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6083
timestamp 1712622712
transform 1 0 732 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6084
timestamp 1712622712
transform 1 0 684 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6085
timestamp 1712622712
transform 1 0 604 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6086
timestamp 1712622712
transform 1 0 564 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_6087
timestamp 1712622712
transform 1 0 540 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_6088
timestamp 1712622712
transform 1 0 508 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_6089
timestamp 1712622712
transform 1 0 804 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6090
timestamp 1712622712
transform 1 0 804 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6091
timestamp 1712622712
transform 1 0 740 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6092
timestamp 1712622712
transform 1 0 700 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6093
timestamp 1712622712
transform 1 0 700 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6094
timestamp 1712622712
transform 1 0 980 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6095
timestamp 1712622712
transform 1 0 892 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6096
timestamp 1712622712
transform 1 0 3420 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_6097
timestamp 1712622712
transform 1 0 3388 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_6098
timestamp 1712622712
transform 1 0 3300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_6099
timestamp 1712622712
transform 1 0 3260 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_6100
timestamp 1712622712
transform 1 0 3428 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_6101
timestamp 1712622712
transform 1 0 2092 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6102
timestamp 1712622712
transform 1 0 2084 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6103
timestamp 1712622712
transform 1 0 2004 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6104
timestamp 1712622712
transform 1 0 1916 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_6105
timestamp 1712622712
transform 1 0 3108 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6106
timestamp 1712622712
transform 1 0 2900 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6107
timestamp 1712622712
transform 1 0 2876 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6108
timestamp 1712622712
transform 1 0 2820 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_6109
timestamp 1712622712
transform 1 0 2692 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_6110
timestamp 1712622712
transform 1 0 2692 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_6111
timestamp 1712622712
transform 1 0 2612 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_6112
timestamp 1712622712
transform 1 0 2604 0 1 2815
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1712622712
transform 1 0 3200 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1712622712
transform 1 0 2104 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1712622712
transform 1 0 1488 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1712622712
transform 1 0 1800 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1712622712
transform 1 0 2600 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1712622712
transform 1 0 624 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1712622712
transform 1 0 2328 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1712622712
transform 1 0 784 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1712622712
transform 1 0 2040 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1712622712
transform 1 0 1904 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1712622712
transform 1 0 168 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1712622712
transform 1 0 288 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1712622712
transform 1 0 2464 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1712622712
transform 1 0 2488 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1712622712
transform 1 0 2488 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1712622712
transform 1 0 1272 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1712622712
transform 1 0 1096 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1712622712
transform 1 0 1136 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1712622712
transform 1 0 1064 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1712622712
transform 1 0 848 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1712622712
transform 1 0 1352 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1712622712
transform 1 0 1288 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1712622712
transform 1 0 784 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1712622712
transform 1 0 736 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1712622712
transform 1 0 712 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1712622712
transform 1 0 584 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1712622712
transform 1 0 736 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1712622712
transform 1 0 512 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1712622712
transform 1 0 1024 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1712622712
transform 1 0 456 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1712622712
transform 1 0 448 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1712622712
transform 1 0 344 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1712622712
transform 1 0 544 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1712622712
transform 1 0 320 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1712622712
transform 1 0 1224 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1712622712
transform 1 0 352 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1712622712
transform 1 0 352 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1712622712
transform 1 0 168 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1712622712
transform 1 0 328 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1712622712
transform 1 0 88 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1712622712
transform 1 0 192 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1712622712
transform 1 0 1160 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1712622712
transform 1 0 288 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1712622712
transform 1 0 344 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1712622712
transform 1 0 216 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1712622712
transform 1 0 328 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1712622712
transform 1 0 816 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1712622712
transform 1 0 112 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1712622712
transform 1 0 144 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1712622712
transform 1 0 1104 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1712622712
transform 1 0 360 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1712622712
transform 1 0 208 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1712622712
transform 1 0 144 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1712622712
transform 1 0 136 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1712622712
transform 1 0 824 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1712622712
transform 1 0 1112 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1712622712
transform 1 0 448 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1712622712
transform 1 0 424 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1712622712
transform 1 0 152 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1712622712
transform 1 0 248 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1712622712
transform 1 0 96 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1712622712
transform 1 0 704 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1712622712
transform 1 0 1336 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1712622712
transform 1 0 296 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1712622712
transform 1 0 96 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1712622712
transform 1 0 192 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1712622712
transform 1 0 576 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1712622712
transform 1 0 1120 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1712622712
transform 1 0 544 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1712622712
transform 1 0 432 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1712622712
transform 1 0 136 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1712622712
transform 1 0 328 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1712622712
transform 1 0 664 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1712622712
transform 1 0 136 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1712622712
transform 1 0 96 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1712622712
transform 1 0 1240 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1712622712
transform 1 0 240 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1712622712
transform 1 0 344 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1712622712
transform 1 0 176 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1712622712
transform 1 0 304 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1712622712
transform 1 0 496 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1712622712
transform 1 0 160 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1712622712
transform 1 0 640 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1712622712
transform 1 0 576 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1712622712
transform 1 0 408 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1712622712
transform 1 0 440 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1712622712
transform 1 0 568 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1712622712
transform 1 0 568 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_88
timestamp 1712622712
transform 1 0 1224 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_89
timestamp 1712622712
transform 1 0 912 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1712622712
transform 1 0 864 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_91
timestamp 1712622712
transform 1 0 816 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_92
timestamp 1712622712
transform 1 0 864 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1712622712
transform 1 0 808 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_94
timestamp 1712622712
transform 1 0 744 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_95
timestamp 1712622712
transform 1 0 1200 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1712622712
transform 1 0 1160 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_97
timestamp 1712622712
transform 1 0 1032 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_98
timestamp 1712622712
transform 1 0 1096 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1712622712
transform 1 0 1040 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_100
timestamp 1712622712
transform 1 0 1152 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_101
timestamp 1712622712
transform 1 0 1056 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1712622712
transform 1 0 984 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_103
timestamp 1712622712
transform 1 0 1464 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1712622712
transform 1 0 1416 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1712622712
transform 1 0 1392 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_106
timestamp 1712622712
transform 1 0 1232 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_107
timestamp 1712622712
transform 1 0 1088 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_108
timestamp 1712622712
transform 1 0 1824 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_109
timestamp 1712622712
transform 1 0 1712 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_110
timestamp 1712622712
transform 1 0 1768 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_111
timestamp 1712622712
transform 1 0 1640 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_112
timestamp 1712622712
transform 1 0 1656 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1712622712
transform 1 0 1648 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_114
timestamp 1712622712
transform 1 0 1600 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_115
timestamp 1712622712
transform 1 0 1344 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_116
timestamp 1712622712
transform 1 0 2024 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_117
timestamp 1712622712
transform 1 0 2056 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1712622712
transform 1 0 2168 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_119
timestamp 1712622712
transform 1 0 2120 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_120
timestamp 1712622712
transform 1 0 1984 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1712622712
transform 1 0 1872 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_122
timestamp 1712622712
transform 1 0 2320 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1712622712
transform 1 0 2440 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1712622712
transform 1 0 2264 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1712622712
transform 1 0 2368 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_126
timestamp 1712622712
transform 1 0 2216 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_127
timestamp 1712622712
transform 1 0 2128 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_128
timestamp 1712622712
transform 1 0 2048 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_129
timestamp 1712622712
transform 1 0 1280 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_130
timestamp 1712622712
transform 1 0 2488 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_131
timestamp 1712622712
transform 1 0 2512 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_132
timestamp 1712622712
transform 1 0 2304 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_133
timestamp 1712622712
transform 1 0 2440 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_134
timestamp 1712622712
transform 1 0 2096 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_135
timestamp 1712622712
transform 1 0 2144 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_136
timestamp 1712622712
transform 1 0 2400 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_137
timestamp 1712622712
transform 1 0 2504 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_138
timestamp 1712622712
transform 1 0 2440 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_139
timestamp 1712622712
transform 1 0 2152 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_140
timestamp 1712622712
transform 1 0 2304 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_141
timestamp 1712622712
transform 1 0 2024 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_142
timestamp 1712622712
transform 1 0 2104 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_143
timestamp 1712622712
transform 1 0 2456 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_144
timestamp 1712622712
transform 1 0 2536 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_145
timestamp 1712622712
transform 1 0 2560 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_146
timestamp 1712622712
transform 1 0 2176 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_147
timestamp 1712622712
transform 1 0 2280 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_148
timestamp 1712622712
transform 1 0 2040 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_149
timestamp 1712622712
transform 1 0 1952 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_150
timestamp 1712622712
transform 1 0 1784 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_151
timestamp 1712622712
transform 1 0 1728 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_152
timestamp 1712622712
transform 1 0 1832 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_153
timestamp 1712622712
transform 1 0 1776 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_154
timestamp 1712622712
transform 1 0 1840 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_155
timestamp 1712622712
transform 1 0 1816 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_156
timestamp 1712622712
transform 1 0 1816 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_157
timestamp 1712622712
transform 1 0 1360 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_158
timestamp 1712622712
transform 1 0 2304 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_159
timestamp 1712622712
transform 1 0 1968 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_160
timestamp 1712622712
transform 1 0 1960 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_161
timestamp 1712622712
transform 1 0 1912 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_162
timestamp 1712622712
transform 1 0 1960 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_163
timestamp 1712622712
transform 1 0 1824 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_164
timestamp 1712622712
transform 1 0 1840 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_165
timestamp 1712622712
transform 1 0 1976 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_166
timestamp 1712622712
transform 1 0 2280 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_167
timestamp 1712622712
transform 1 0 2128 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_168
timestamp 1712622712
transform 1 0 2168 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_169
timestamp 1712622712
transform 1 0 2128 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_170
timestamp 1712622712
transform 1 0 2128 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_171
timestamp 1712622712
transform 1 0 2184 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_172
timestamp 1712622712
transform 1 0 2344 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_173
timestamp 1712622712
transform 1 0 2480 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_174
timestamp 1712622712
transform 1 0 2456 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_175
timestamp 1712622712
transform 1 0 2408 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_176
timestamp 1712622712
transform 1 0 2336 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_177
timestamp 1712622712
transform 1 0 2376 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_178
timestamp 1712622712
transform 1 0 2320 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_179
timestamp 1712622712
transform 1 0 2296 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_180
timestamp 1712622712
transform 1 0 2544 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_181
timestamp 1712622712
transform 1 0 2488 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_182
timestamp 1712622712
transform 1 0 2544 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_183
timestamp 1712622712
transform 1 0 2664 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_184
timestamp 1712622712
transform 1 0 2096 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_185
timestamp 1712622712
transform 1 0 1928 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_186
timestamp 1712622712
transform 1 0 2400 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_187
timestamp 1712622712
transform 1 0 2592 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_188
timestamp 1712622712
transform 1 0 2496 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_189
timestamp 1712622712
transform 1 0 2840 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_190
timestamp 1712622712
transform 1 0 2608 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_191
timestamp 1712622712
transform 1 0 2488 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_192
timestamp 1712622712
transform 1 0 2664 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_193
timestamp 1712622712
transform 1 0 2560 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_194
timestamp 1712622712
transform 1 0 2512 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_195
timestamp 1712622712
transform 1 0 2832 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_196
timestamp 1712622712
transform 1 0 2600 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_197
timestamp 1712622712
transform 1 0 3168 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_198
timestamp 1712622712
transform 1 0 2744 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_199
timestamp 1712622712
transform 1 0 2904 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_200
timestamp 1712622712
transform 1 0 3072 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_201
timestamp 1712622712
transform 1 0 3232 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_202
timestamp 1712622712
transform 1 0 3352 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_203
timestamp 1712622712
transform 1 0 3312 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_204
timestamp 1712622712
transform 1 0 3288 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_205
timestamp 1712622712
transform 1 0 3016 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_206
timestamp 1712622712
transform 1 0 3056 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_207
timestamp 1712622712
transform 1 0 2928 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_208
timestamp 1712622712
transform 1 0 3048 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_209
timestamp 1712622712
transform 1 0 3016 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_210
timestamp 1712622712
transform 1 0 2560 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_211
timestamp 1712622712
transform 1 0 2608 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_212
timestamp 1712622712
transform 1 0 2880 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_213
timestamp 1712622712
transform 1 0 952 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_214
timestamp 1712622712
transform 1 0 1448 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_215
timestamp 1712622712
transform 1 0 1584 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_216
timestamp 1712622712
transform 1 0 1896 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_217
timestamp 1712622712
transform 1 0 3152 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_218
timestamp 1712622712
transform 1 0 2392 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_219
timestamp 1712622712
transform 1 0 1144 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_220
timestamp 1712622712
transform 1 0 3264 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_221
timestamp 1712622712
transform 1 0 3272 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_222
timestamp 1712622712
transform 1 0 3240 0 -1 2370
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1712622712
transform 1 0 2648 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1712622712
transform 1 0 1520 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1712622712
transform 1 0 1440 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1712622712
transform 1 0 960 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1712622712
transform 1 0 224 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1712622712
transform 1 0 1512 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1712622712
transform 1 0 408 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1712622712
transform 1 0 400 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1712622712
transform 1 0 856 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1712622712
transform 1 0 1624 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1712622712
transform 1 0 760 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1712622712
transform 1 0 2016 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1712622712
transform 1 0 1640 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1712622712
transform 1 0 1592 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1712622712
transform 1 0 1520 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1712622712
transform 1 0 344 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1712622712
transform 1 0 1304 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1712622712
transform 1 0 1976 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1712622712
transform 1 0 1408 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1712622712
transform 1 0 1792 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1712622712
transform 1 0 96 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1712622712
transform 1 0 1752 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1712622712
transform 1 0 1112 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1712622712
transform 1 0 960 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1712622712
transform 1 0 496 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1712622712
transform 1 0 696 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1712622712
transform 1 0 400 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1712622712
transform 1 0 512 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1712622712
transform 1 0 320 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1712622712
transform 1 0 632 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1712622712
transform 1 0 272 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1712622712
transform 1 0 360 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1712622712
transform 1 0 592 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1712622712
transform 1 0 864 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1712622712
transform 1 0 296 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1712622712
transform 1 0 320 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1712622712
transform 1 0 608 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1712622712
transform 1 0 696 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1712622712
transform 1 0 224 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1712622712
transform 1 0 720 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1712622712
transform 1 0 800 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1712622712
transform 1 0 288 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1712622712
transform 1 0 624 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1712622712
transform 1 0 624 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1712622712
transform 1 0 304 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1712622712
transform 1 0 688 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1712622712
transform 1 0 784 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1712622712
transform 1 0 264 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_48
timestamp 1712622712
transform 1 0 448 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_49
timestamp 1712622712
transform 1 0 696 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_50
timestamp 1712622712
transform 1 0 280 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_51
timestamp 1712622712
transform 1 0 632 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_52
timestamp 1712622712
transform 1 0 848 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_53
timestamp 1712622712
transform 1 0 384 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_54
timestamp 1712622712
transform 1 0 640 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1712622712
transform 1 0 816 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_56
timestamp 1712622712
transform 1 0 352 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_57
timestamp 1712622712
transform 1 0 304 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_58
timestamp 1712622712
transform 1 0 712 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_59
timestamp 1712622712
transform 1 0 184 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_60
timestamp 1712622712
transform 1 0 1088 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_61
timestamp 1712622712
transform 1 0 384 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_62
timestamp 1712622712
transform 1 0 728 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_63
timestamp 1712622712
transform 1 0 328 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_64
timestamp 1712622712
transform 1 0 896 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_65
timestamp 1712622712
transform 1 0 976 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_66
timestamp 1712622712
transform 1 0 968 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_67
timestamp 1712622712
transform 1 0 1088 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_68
timestamp 1712622712
transform 1 0 1032 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_69
timestamp 1712622712
transform 1 0 1152 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_70
timestamp 1712622712
transform 1 0 1136 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_71
timestamp 1712622712
transform 1 0 1344 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_72
timestamp 1712622712
transform 1 0 1528 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_73
timestamp 1712622712
transform 1 0 1512 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_74
timestamp 1712622712
transform 1 0 1400 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_75
timestamp 1712622712
transform 1 0 1360 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_76
timestamp 1712622712
transform 1 0 1392 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_77
timestamp 1712622712
transform 1 0 1616 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_78
timestamp 1712622712
transform 1 0 1736 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_79
timestamp 1712622712
transform 1 0 1768 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_80
timestamp 1712622712
transform 1 0 1664 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_81
timestamp 1712622712
transform 1 0 1632 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_82
timestamp 1712622712
transform 1 0 1712 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_83
timestamp 1712622712
transform 1 0 2152 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_84
timestamp 1712622712
transform 1 0 1848 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_85
timestamp 1712622712
transform 1 0 1808 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_86
timestamp 1712622712
transform 1 0 2224 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_87
timestamp 1712622712
transform 1 0 1944 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_88
timestamp 1712622712
transform 1 0 1904 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_89
timestamp 1712622712
transform 1 0 2392 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_90
timestamp 1712622712
transform 1 0 2096 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_91
timestamp 1712622712
transform 1 0 1856 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_92
timestamp 1712622712
transform 1 0 2448 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_93
timestamp 1712622712
transform 1 0 2432 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_94
timestamp 1712622712
transform 1 0 2152 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_95
timestamp 1712622712
transform 1 0 2376 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_96
timestamp 1712622712
transform 1 0 1448 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_97
timestamp 1712622712
transform 1 0 1456 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_98
timestamp 1712622712
transform 1 0 2272 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_99
timestamp 1712622712
transform 1 0 2120 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_100
timestamp 1712622712
transform 1 0 2272 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_101
timestamp 1712622712
transform 1 0 2184 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_102
timestamp 1712622712
transform 1 0 2064 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_103
timestamp 1712622712
transform 1 0 2168 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_104
timestamp 1712622712
transform 1 0 1800 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_105
timestamp 1712622712
transform 1 0 1704 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_106
timestamp 1712622712
transform 1 0 1904 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_107
timestamp 1712622712
transform 1 0 1832 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_108
timestamp 1712622712
transform 1 0 1936 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_109
timestamp 1712622712
transform 1 0 2184 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_110
timestamp 1712622712
transform 1 0 2336 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_111
timestamp 1712622712
transform 1 0 2008 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_112
timestamp 1712622712
transform 1 0 2144 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_113
timestamp 1712622712
transform 1 0 2248 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_114
timestamp 1712622712
transform 1 0 2136 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_115
timestamp 1712622712
transform 1 0 2272 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_116
timestamp 1712622712
transform 1 0 2448 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_117
timestamp 1712622712
transform 1 0 2240 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_118
timestamp 1712622712
transform 1 0 2384 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_119
timestamp 1712622712
transform 1 0 2416 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_120
timestamp 1712622712
transform 1 0 2384 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_121
timestamp 1712622712
transform 1 0 2456 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_122
timestamp 1712622712
transform 1 0 2584 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_123
timestamp 1712622712
transform 1 0 2440 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_124
timestamp 1712622712
transform 1 0 2544 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_125
timestamp 1712622712
transform 1 0 2640 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_126
timestamp 1712622712
transform 1 0 2544 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_127
timestamp 1712622712
transform 1 0 2640 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_128
timestamp 1712622712
transform 1 0 2016 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_129
timestamp 1712622712
transform 1 0 1896 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_130
timestamp 1712622712
transform 1 0 1312 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_131
timestamp 1712622712
transform 1 0 2696 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_132
timestamp 1712622712
transform 1 0 3000 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_133
timestamp 1712622712
transform 1 0 3024 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_134
timestamp 1712622712
transform 1 0 2632 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_135
timestamp 1712622712
transform 1 0 1728 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_136
timestamp 1712622712
transform 1 0 2976 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_137
timestamp 1712622712
transform 1 0 2552 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_138
timestamp 1712622712
transform 1 0 2904 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_139
timestamp 1712622712
transform 1 0 2960 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_140
timestamp 1712622712
transform 1 0 3064 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_141
timestamp 1712622712
transform 1 0 2608 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_142
timestamp 1712622712
transform 1 0 1800 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_143
timestamp 1712622712
transform 1 0 2792 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_144
timestamp 1712622712
transform 1 0 2712 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_145
timestamp 1712622712
transform 1 0 2904 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_146
timestamp 1712622712
transform 1 0 2840 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_147
timestamp 1712622712
transform 1 0 2784 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_148
timestamp 1712622712
transform 1 0 2600 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_149
timestamp 1712622712
transform 1 0 2864 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_150
timestamp 1712622712
transform 1 0 2528 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_151
timestamp 1712622712
transform 1 0 2640 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_152
timestamp 1712622712
transform 1 0 2848 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_153
timestamp 1712622712
transform 1 0 2792 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_154
timestamp 1712622712
transform 1 0 2576 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_155
timestamp 1712622712
transform 1 0 2840 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_156
timestamp 1712622712
transform 1 0 3176 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_157
timestamp 1712622712
transform 1 0 3344 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_158
timestamp 1712622712
transform 1 0 3376 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_159
timestamp 1712622712
transform 1 0 3256 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_160
timestamp 1712622712
transform 1 0 3160 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_161
timestamp 1712622712
transform 1 0 3392 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_162
timestamp 1712622712
transform 1 0 3368 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_163
timestamp 1712622712
transform 1 0 3312 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_164
timestamp 1712622712
transform 1 0 2872 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_165
timestamp 1712622712
transform 1 0 896 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_166
timestamp 1712622712
transform 1 0 1640 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_167
timestamp 1712622712
transform 1 0 1760 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_168
timestamp 1712622712
transform 1 0 1976 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_169
timestamp 1712622712
transform 1 0 2840 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_170
timestamp 1712622712
transform 1 0 3120 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_171
timestamp 1712622712
transform 1 0 3128 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_172
timestamp 1712622712
transform 1 0 3216 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_173
timestamp 1712622712
transform 1 0 2352 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_174
timestamp 1712622712
transform 1 0 1928 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_175
timestamp 1712622712
transform 1 0 536 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_176
timestamp 1712622712
transform 1 0 888 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_177
timestamp 1712622712
transform 1 0 824 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_178
timestamp 1712622712
transform 1 0 1864 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_179
timestamp 1712622712
transform 1 0 1200 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_180
timestamp 1712622712
transform 1 0 1416 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_181
timestamp 1712622712
transform 1 0 2240 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_182
timestamp 1712622712
transform 1 0 3024 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_183
timestamp 1712622712
transform 1 0 3392 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_184
timestamp 1712622712
transform 1 0 3328 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_185
timestamp 1712622712
transform 1 0 3128 0 1 2570
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1712622712
transform 1 0 2984 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1712622712
transform 1 0 3184 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1712622712
transform 1 0 968 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1712622712
transform 1 0 992 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1712622712
transform 1 0 2112 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1712622712
transform 1 0 1424 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1712622712
transform 1 0 384 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1712622712
transform 1 0 776 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1712622712
transform 1 0 1680 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1712622712
transform 1 0 1896 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1712622712
transform 1 0 872 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1712622712
transform 1 0 1776 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1712622712
transform 1 0 776 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1712622712
transform 1 0 744 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1712622712
transform 1 0 2016 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1712622712
transform 1 0 2504 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1712622712
transform 1 0 2064 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1712622712
transform 1 0 1504 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1712622712
transform 1 0 1848 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1712622712
transform 1 0 1528 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1712622712
transform 1 0 1704 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1712622712
transform 1 0 616 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1712622712
transform 1 0 160 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1712622712
transform 1 0 352 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1712622712
transform 1 0 1496 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1712622712
transform 1 0 1808 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1712622712
transform 1 0 128 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1712622712
transform 1 0 1928 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1712622712
transform 1 0 1512 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1712622712
transform 1 0 1536 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1712622712
transform 1 0 1352 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1712622712
transform 1 0 1264 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1712622712
transform 1 0 1384 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1712622712
transform 1 0 3232 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1712622712
transform 1 0 1368 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1712622712
transform 1 0 1168 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1712622712
transform 1 0 1536 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1712622712
transform 1 0 1304 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1712622712
transform 1 0 1192 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1712622712
transform 1 0 1176 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1712622712
transform 1 0 1272 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1712622712
transform 1 0 784 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1712622712
transform 1 0 992 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1712622712
transform 1 0 656 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1712622712
transform 1 0 904 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1712622712
transform 1 0 1192 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1712622712
transform 1 0 616 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1712622712
transform 1 0 832 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1712622712
transform 1 0 1144 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1712622712
transform 1 0 608 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1712622712
transform 1 0 112 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1712622712
transform 1 0 872 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1712622712
transform 1 0 1248 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1712622712
transform 1 0 920 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1712622712
transform 1 0 96 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1712622712
transform 1 0 912 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1712622712
transform 1 0 1120 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1712622712
transform 1 0 944 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1712622712
transform 1 0 872 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1712622712
transform 1 0 1024 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1712622712
transform 1 0 1368 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1712622712
transform 1 0 1288 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1712622712
transform 1 0 904 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1712622712
transform 1 0 936 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1712622712
transform 1 0 1128 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1712622712
transform 1 0 1160 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1712622712
transform 1 0 832 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1712622712
transform 1 0 2744 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1712622712
transform 1 0 760 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1712622712
transform 1 0 976 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1712622712
transform 1 0 664 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1712622712
transform 1 0 1048 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1712622712
transform 1 0 504 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1712622712
transform 1 0 1128 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1712622712
transform 1 0 1200 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1712622712
transform 1 0 472 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1712622712
transform 1 0 1280 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1712622712
transform 1 0 1344 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1712622712
transform 1 0 1512 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1712622712
transform 1 0 1256 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1712622712
transform 1 0 216 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1712622712
transform 1 0 1736 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1712622712
transform 1 0 1296 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1712622712
transform 1 0 880 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1712622712
transform 1 0 2080 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1712622712
transform 1 0 1912 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1712622712
transform 1 0 1272 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1712622712
transform 1 0 536 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1712622712
transform 1 0 1704 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1712622712
transform 1 0 1336 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1712622712
transform 1 0 1808 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1712622712
transform 1 0 592 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1712622712
transform 1 0 1640 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1712622712
transform 1 0 1376 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1712622712
transform 1 0 1640 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1712622712
transform 1 0 1400 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1712622712
transform 1 0 1256 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1712622712
transform 1 0 544 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1712622712
transform 1 0 2704 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1712622712
transform 1 0 1992 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1712622712
transform 1 0 1848 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1712622712
transform 1 0 1304 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1712622712
transform 1 0 656 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1712622712
transform 1 0 2016 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1712622712
transform 1 0 1520 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1712622712
transform 1 0 856 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1712622712
transform 1 0 1944 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1712622712
transform 1 0 1712 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1712622712
transform 1 0 1664 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1712622712
transform 1 0 1352 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1712622712
transform 1 0 2464 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1712622712
transform 1 0 1888 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1712622712
transform 1 0 1560 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1712622712
transform 1 0 2504 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1712622712
transform 1 0 2304 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1712622712
transform 1 0 1760 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1712622712
transform 1 0 2688 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1712622712
transform 1 0 2400 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1712622712
transform 1 0 2024 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1712622712
transform 1 0 2672 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1712622712
transform 1 0 2280 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1712622712
transform 1 0 2432 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1712622712
transform 1 0 2560 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1712622712
transform 1 0 2672 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1712622712
transform 1 0 2760 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1712622712
transform 1 0 2520 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_126
timestamp 1712622712
transform 1 0 1496 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_127
timestamp 1712622712
transform 1 0 3080 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_128
timestamp 1712622712
transform 1 0 2688 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_129
timestamp 1712622712
transform 1 0 2736 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_130
timestamp 1712622712
transform 1 0 2848 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_131
timestamp 1712622712
transform 1 0 2928 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_132
timestamp 1712622712
transform 1 0 3096 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_133
timestamp 1712622712
transform 1 0 3040 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_134
timestamp 1712622712
transform 1 0 2712 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_135
timestamp 1712622712
transform 1 0 2736 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_136
timestamp 1712622712
transform 1 0 2760 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_137
timestamp 1712622712
transform 1 0 3144 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_138
timestamp 1712622712
transform 1 0 2912 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_139
timestamp 1712622712
transform 1 0 2872 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_140
timestamp 1712622712
transform 1 0 2736 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_141
timestamp 1712622712
transform 1 0 3280 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_142
timestamp 1712622712
transform 1 0 3256 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_143
timestamp 1712622712
transform 1 0 2800 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_144
timestamp 1712622712
transform 1 0 2664 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_145
timestamp 1712622712
transform 1 0 3216 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_146
timestamp 1712622712
transform 1 0 3280 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_147
timestamp 1712622712
transform 1 0 3328 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_148
timestamp 1712622712
transform 1 0 2072 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_149
timestamp 1712622712
transform 1 0 2848 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_150
timestamp 1712622712
transform 1 0 2752 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_151
timestamp 1712622712
transform 1 0 2696 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_152
timestamp 1712622712
transform 1 0 2824 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_153
timestamp 1712622712
transform 1 0 2768 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_154
timestamp 1712622712
transform 1 0 3144 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_155
timestamp 1712622712
transform 1 0 3320 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_156
timestamp 1712622712
transform 1 0 3048 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_157
timestamp 1712622712
transform 1 0 3280 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_158
timestamp 1712622712
transform 1 0 3256 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_159
timestamp 1712622712
transform 1 0 3400 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_160
timestamp 1712622712
transform 1 0 3160 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_161
timestamp 1712622712
transform 1 0 3232 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_162
timestamp 1712622712
transform 1 0 2824 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_163
timestamp 1712622712
transform 1 0 2560 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_164
timestamp 1712622712
transform 1 0 2464 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_165
timestamp 1712622712
transform 1 0 768 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_166
timestamp 1712622712
transform 1 0 792 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_167
timestamp 1712622712
transform 1 0 896 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_168
timestamp 1712622712
transform 1 0 1672 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_169
timestamp 1712622712
transform 1 0 1800 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_170
timestamp 1712622712
transform 1 0 1904 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_171
timestamp 1712622712
transform 1 0 1112 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_172
timestamp 1712622712
transform 1 0 896 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_173
timestamp 1712622712
transform 1 0 688 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_174
timestamp 1712622712
transform 1 0 600 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_175
timestamp 1712622712
transform 1 0 472 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_176
timestamp 1712622712
transform 1 0 424 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_177
timestamp 1712622712
transform 1 0 448 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_178
timestamp 1712622712
transform 1 0 344 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_179
timestamp 1712622712
transform 1 0 144 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_180
timestamp 1712622712
transform 1 0 88 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_181
timestamp 1712622712
transform 1 0 120 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_182
timestamp 1712622712
transform 1 0 928 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_183
timestamp 1712622712
transform 1 0 1136 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_184
timestamp 1712622712
transform 1 0 1240 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_185
timestamp 1712622712
transform 1 0 1320 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_186
timestamp 1712622712
transform 1 0 1344 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_187
timestamp 1712622712
transform 1 0 1560 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_188
timestamp 1712622712
transform 1 0 1648 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_189
timestamp 1712622712
transform 1 0 1824 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_190
timestamp 1712622712
transform 1 0 1776 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_191
timestamp 1712622712
transform 1 0 2064 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_192
timestamp 1712622712
transform 1 0 2160 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_193
timestamp 1712622712
transform 1 0 2312 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_194
timestamp 1712622712
transform 1 0 2016 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_195
timestamp 1712622712
transform 1 0 2376 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_196
timestamp 1712622712
transform 1 0 2528 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_197
timestamp 1712622712
transform 1 0 2752 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_198
timestamp 1712622712
transform 1 0 2552 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_199
timestamp 1712622712
transform 1 0 2800 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_200
timestamp 1712622712
transform 1 0 3064 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_201
timestamp 1712622712
transform 1 0 2704 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_202
timestamp 1712622712
transform 1 0 3152 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_203
timestamp 1712622712
transform 1 0 2496 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_204
timestamp 1712622712
transform 1 0 824 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_205
timestamp 1712622712
transform 1 0 784 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_206
timestamp 1712622712
transform 1 0 1728 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_207
timestamp 1712622712
transform 1 0 2064 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_208
timestamp 1712622712
transform 1 0 1272 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_209
timestamp 1712622712
transform 1 0 2248 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_210
timestamp 1712622712
transform 1 0 3400 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_211
timestamp 1712622712
transform 1 0 3296 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_212
timestamp 1712622712
transform 1 0 3400 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_213
timestamp 1712622712
transform 1 0 3280 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_214
timestamp 1712622712
transform 1 0 3272 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_215
timestamp 1712622712
transform 1 0 3312 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_216
timestamp 1712622712
transform 1 0 3392 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_217
timestamp 1712622712
transform 1 0 3296 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_218
timestamp 1712622712
transform 1 0 3312 0 1 770
box -8 -3 32 105
use NOR3X1  NOR3X1_0
timestamp 1712622712
transform 1 0 3168 0 -1 1970
box -7 -3 68 105
use OAI21X1  OAI21X1_0
timestamp 1712622712
transform 1 0 3152 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1712622712
transform 1 0 1728 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1712622712
transform 1 0 2184 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1712622712
transform 1 0 1016 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1712622712
transform 1 0 1640 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1712622712
transform 1 0 1872 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1712622712
transform 1 0 1400 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1712622712
transform 1 0 1640 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1712622712
transform 1 0 1792 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1712622712
transform 1 0 1528 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1712622712
transform 1 0 896 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1712622712
transform 1 0 1424 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1712622712
transform 1 0 2576 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1712622712
transform 1 0 2696 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1712622712
transform 1 0 1224 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1712622712
transform 1 0 1968 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1712622712
transform 1 0 1592 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1712622712
transform 1 0 2144 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1712622712
transform 1 0 240 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1712622712
transform 1 0 608 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1712622712
transform 1 0 112 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1712622712
transform 1 0 1608 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1712622712
transform 1 0 312 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1712622712
transform 1 0 1424 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1712622712
transform 1 0 1288 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1712622712
transform 1 0 1912 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1712622712
transform 1 0 1640 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1712622712
transform 1 0 96 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1712622712
transform 1 0 656 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1712622712
transform 1 0 1240 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1712622712
transform 1 0 1928 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1712622712
transform 1 0 2040 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1712622712
transform 1 0 1336 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1712622712
transform 1 0 1496 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1712622712
transform 1 0 1448 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1712622712
transform 1 0 1568 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1712622712
transform 1 0 1312 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1712622712
transform 1 0 1336 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1712622712
transform 1 0 1312 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1712622712
transform 1 0 896 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1712622712
transform 1 0 1256 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1712622712
transform 1 0 1208 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1712622712
transform 1 0 1328 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1712622712
transform 1 0 1136 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1712622712
transform 1 0 1040 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1712622712
transform 1 0 864 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1712622712
transform 1 0 720 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1712622712
transform 1 0 1080 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1712622712
transform 1 0 1136 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1712622712
transform 1 0 1384 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1712622712
transform 1 0 1152 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1712622712
transform 1 0 1088 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1712622712
transform 1 0 784 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1712622712
transform 1 0 656 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1712622712
transform 1 0 840 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1712622712
transform 1 0 1176 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1712622712
transform 1 0 1344 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1712622712
transform 1 0 992 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1712622712
transform 1 0 1328 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1712622712
transform 1 0 1392 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1712622712
transform 1 0 456 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1712622712
transform 1 0 584 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1712622712
transform 1 0 1200 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1712622712
transform 1 0 856 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1712622712
transform 1 0 1040 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1712622712
transform 1 0 856 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1712622712
transform 1 0 1232 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1712622712
transform 1 0 392 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1712622712
transform 1 0 392 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1712622712
transform 1 0 752 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1712622712
transform 1 0 624 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1712622712
transform 1 0 664 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1712622712
transform 1 0 720 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1712622712
transform 1 0 312 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1712622712
transform 1 0 280 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1712622712
transform 1 0 1008 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1712622712
transform 1 0 888 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1712622712
transform 1 0 952 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1712622712
transform 1 0 560 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1712622712
transform 1 0 264 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1712622712
transform 1 0 240 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1712622712
transform 1 0 976 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1712622712
transform 1 0 640 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1712622712
transform 1 0 1096 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1712622712
transform 1 0 216 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1712622712
transform 1 0 208 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1712622712
transform 1 0 680 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1712622712
transform 1 0 792 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1712622712
transform 1 0 704 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1712622712
transform 1 0 88 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1712622712
transform 1 0 144 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1712622712
transform 1 0 624 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1712622712
transform 1 0 720 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1712622712
transform 1 0 624 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1712622712
transform 1 0 144 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1712622712
transform 1 0 136 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1712622712
transform 1 0 592 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1712622712
transform 1 0 792 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1712622712
transform 1 0 752 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1712622712
transform 1 0 520 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1712622712
transform 1 0 216 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1712622712
transform 1 0 952 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1712622712
transform 1 0 872 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1712622712
transform 1 0 960 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1712622712
transform 1 0 960 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1712622712
transform 1 0 200 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1712622712
transform 1 0 936 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1712622712
transform 1 0 800 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1712622712
transform 1 0 944 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1712622712
transform 1 0 1000 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1712622712
transform 1 0 1144 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1712622712
transform 1 0 1096 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1712622712
transform 1 0 664 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1712622712
transform 1 0 704 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1712622712
transform 1 0 592 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1712622712
transform 1 0 648 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1712622712
transform 1 0 1200 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1712622712
transform 1 0 1288 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1712622712
transform 1 0 816 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1712622712
transform 1 0 1016 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1712622712
transform 1 0 864 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1712622712
transform 1 0 920 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1712622712
transform 1 0 1248 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1712622712
transform 1 0 1408 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1712622712
transform 1 0 1128 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1712622712
transform 1 0 1144 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1712622712
transform 1 0 1448 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1712622712
transform 1 0 1192 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1712622712
transform 1 0 1456 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1712622712
transform 1 0 1488 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1712622712
transform 1 0 1320 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1712622712
transform 1 0 1336 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1712622712
transform 1 0 1456 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1712622712
transform 1 0 1656 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1712622712
transform 1 0 1744 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1712622712
transform 1 0 1640 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1712622712
transform 1 0 1696 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1712622712
transform 1 0 1656 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1712622712
transform 1 0 1784 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1712622712
transform 1 0 2072 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1712622712
transform 1 0 1976 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1712622712
transform 1 0 1960 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1712622712
transform 1 0 1792 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1712622712
transform 1 0 1848 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1712622712
transform 1 0 2224 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1712622712
transform 1 0 1864 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1712622712
transform 1 0 1864 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1712622712
transform 1 0 1688 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1712622712
transform 1 0 2040 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1712622712
transform 1 0 2272 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1712622712
transform 1 0 1600 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1712622712
transform 1 0 2488 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1712622712
transform 1 0 1584 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1712622712
transform 1 0 1968 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1712622712
transform 1 0 1504 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1712622712
transform 1 0 1600 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1712622712
transform 1 0 2296 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1712622712
transform 1 0 2304 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1712622712
transform 1 0 1984 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1712622712
transform 1 0 2240 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1712622712
transform 1 0 2056 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1712622712
transform 1 0 2256 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1712622712
transform 1 0 1368 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_163
timestamp 1712622712
transform 1 0 2232 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_164
timestamp 1712622712
transform 1 0 2304 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_165
timestamp 1712622712
transform 1 0 1984 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_166
timestamp 1712622712
transform 1 0 2376 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_167
timestamp 1712622712
transform 1 0 1920 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_168
timestamp 1712622712
transform 1 0 2320 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_169
timestamp 1712622712
transform 1 0 1664 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_170
timestamp 1712622712
transform 1 0 1608 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_171
timestamp 1712622712
transform 1 0 1912 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_172
timestamp 1712622712
transform 1 0 1840 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_173
timestamp 1712622712
transform 1 0 1760 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_174
timestamp 1712622712
transform 1 0 2024 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_175
timestamp 1712622712
transform 1 0 1720 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_176
timestamp 1712622712
transform 1 0 2104 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_177
timestamp 1712622712
transform 1 0 1976 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_178
timestamp 1712622712
transform 1 0 2024 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_179
timestamp 1712622712
transform 1 0 2192 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_180
timestamp 1712622712
transform 1 0 2080 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_181
timestamp 1712622712
transform 1 0 2360 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_182
timestamp 1712622712
transform 1 0 2176 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_183
timestamp 1712622712
transform 1 0 2336 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_184
timestamp 1712622712
transform 1 0 2312 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_185
timestamp 1712622712
transform 1 0 2400 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_186
timestamp 1712622712
transform 1 0 2480 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_187
timestamp 1712622712
transform 1 0 2424 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_188
timestamp 1712622712
transform 1 0 2584 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_189
timestamp 1712622712
transform 1 0 2568 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_190
timestamp 1712622712
transform 1 0 2520 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_191
timestamp 1712622712
transform 1 0 2600 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_192
timestamp 1712622712
transform 1 0 2544 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_193
timestamp 1712622712
transform 1 0 2648 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_194
timestamp 1712622712
transform 1 0 2640 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_195
timestamp 1712622712
transform 1 0 2704 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_196
timestamp 1712622712
transform 1 0 2824 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_197
timestamp 1712622712
transform 1 0 2856 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_198
timestamp 1712622712
transform 1 0 2976 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_199
timestamp 1712622712
transform 1 0 3024 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_200
timestamp 1712622712
transform 1 0 3024 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_201
timestamp 1712622712
transform 1 0 3032 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_202
timestamp 1712622712
transform 1 0 2824 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_203
timestamp 1712622712
transform 1 0 2888 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_204
timestamp 1712622712
transform 1 0 2952 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_205
timestamp 1712622712
transform 1 0 2984 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_206
timestamp 1712622712
transform 1 0 3048 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_207
timestamp 1712622712
transform 1 0 3096 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_208
timestamp 1712622712
transform 1 0 3168 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_209
timestamp 1712622712
transform 1 0 3080 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_210
timestamp 1712622712
transform 1 0 3016 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_211
timestamp 1712622712
transform 1 0 3160 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_212
timestamp 1712622712
transform 1 0 3016 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_213
timestamp 1712622712
transform 1 0 2896 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_214
timestamp 1712622712
transform 1 0 2896 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_215
timestamp 1712622712
transform 1 0 2904 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_216
timestamp 1712622712
transform 1 0 3024 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_217
timestamp 1712622712
transform 1 0 3032 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_218
timestamp 1712622712
transform 1 0 2968 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_219
timestamp 1712622712
transform 1 0 2944 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_220
timestamp 1712622712
transform 1 0 2792 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_221
timestamp 1712622712
transform 1 0 3080 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_222
timestamp 1712622712
transform 1 0 2800 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_223
timestamp 1712622712
transform 1 0 2696 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_224
timestamp 1712622712
transform 1 0 2760 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_225
timestamp 1712622712
transform 1 0 2760 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_226
timestamp 1712622712
transform 1 0 2880 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_227
timestamp 1712622712
transform 1 0 2888 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_228
timestamp 1712622712
transform 1 0 2648 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_229
timestamp 1712622712
transform 1 0 2768 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_230
timestamp 1712622712
transform 1 0 2712 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_231
timestamp 1712622712
transform 1 0 2712 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_232
timestamp 1712622712
transform 1 0 2840 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_233
timestamp 1712622712
transform 1 0 3184 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_234
timestamp 1712622712
transform 1 0 3232 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_235
timestamp 1712622712
transform 1 0 3336 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_236
timestamp 1712622712
transform 1 0 3296 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_237
timestamp 1712622712
transform 1 0 2736 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_238
timestamp 1712622712
transform 1 0 2896 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_239
timestamp 1712622712
transform 1 0 3096 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_240
timestamp 1712622712
transform 1 0 3176 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_241
timestamp 1712622712
transform 1 0 3320 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_242
timestamp 1712622712
transform 1 0 3320 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_243
timestamp 1712622712
transform 1 0 3336 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_244
timestamp 1712622712
transform 1 0 2864 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_245
timestamp 1712622712
transform 1 0 2944 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_246
timestamp 1712622712
transform 1 0 3064 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_247
timestamp 1712622712
transform 1 0 3272 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_248
timestamp 1712622712
transform 1 0 3392 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_249
timestamp 1712622712
transform 1 0 3192 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_250
timestamp 1712622712
transform 1 0 3064 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_251
timestamp 1712622712
transform 1 0 3240 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_252
timestamp 1712622712
transform 1 0 3040 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_253
timestamp 1712622712
transform 1 0 2920 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_254
timestamp 1712622712
transform 1 0 2960 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_255
timestamp 1712622712
transform 1 0 2632 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_256
timestamp 1712622712
transform 1 0 2552 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_257
timestamp 1712622712
transform 1 0 2144 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_258
timestamp 1712622712
transform 1 0 2088 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_259
timestamp 1712622712
transform 1 0 2016 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_260
timestamp 1712622712
transform 1 0 3096 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_261
timestamp 1712622712
transform 1 0 2936 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_262
timestamp 1712622712
transform 1 0 2528 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_263
timestamp 1712622712
transform 1 0 2648 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_264
timestamp 1712622712
transform 1 0 2664 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_265
timestamp 1712622712
transform 1 0 2400 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_266
timestamp 1712622712
transform 1 0 2432 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_267
timestamp 1712622712
transform 1 0 2176 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_268
timestamp 1712622712
transform 1 0 1984 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_269
timestamp 1712622712
transform 1 0 2040 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_270
timestamp 1712622712
transform 1 0 2312 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_271
timestamp 1712622712
transform 1 0 2328 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_272
timestamp 1712622712
transform 1 0 2176 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_273
timestamp 1712622712
transform 1 0 2296 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_274
timestamp 1712622712
transform 1 0 2088 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_275
timestamp 1712622712
transform 1 0 2136 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_276
timestamp 1712622712
transform 1 0 1992 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_277
timestamp 1712622712
transform 1 0 1944 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_278
timestamp 1712622712
transform 1 0 1784 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_279
timestamp 1712622712
transform 1 0 1880 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_280
timestamp 1712622712
transform 1 0 1928 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_281
timestamp 1712622712
transform 1 0 1920 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_282
timestamp 1712622712
transform 1 0 1632 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_283
timestamp 1712622712
transform 1 0 1744 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_284
timestamp 1712622712
transform 1 0 1584 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_285
timestamp 1712622712
transform 1 0 1688 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_286
timestamp 1712622712
transform 1 0 1400 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_287
timestamp 1712622712
transform 1 0 1512 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_288
timestamp 1712622712
transform 1 0 1312 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_289
timestamp 1712622712
transform 1 0 1416 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_290
timestamp 1712622712
transform 1 0 1208 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_291
timestamp 1712622712
transform 1 0 1280 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_292
timestamp 1712622712
transform 1 0 1144 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_293
timestamp 1712622712
transform 1 0 1232 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_294
timestamp 1712622712
transform 1 0 1520 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_295
timestamp 1712622712
transform 1 0 1480 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_296
timestamp 1712622712
transform 1 0 1152 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_297
timestamp 1712622712
transform 1 0 1304 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_298
timestamp 1712622712
transform 1 0 208 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_299
timestamp 1712622712
transform 1 0 1192 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_300
timestamp 1712622712
transform 1 0 216 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_301
timestamp 1712622712
transform 1 0 1088 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_302
timestamp 1712622712
transform 1 0 248 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_303
timestamp 1712622712
transform 1 0 1008 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_304
timestamp 1712622712
transform 1 0 992 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_305
timestamp 1712622712
transform 1 0 1024 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_306
timestamp 1712622712
transform 1 0 368 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_307
timestamp 1712622712
transform 1 0 632 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_308
timestamp 1712622712
transform 1 0 400 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_309
timestamp 1712622712
transform 1 0 576 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_310
timestamp 1712622712
transform 1 0 384 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_311
timestamp 1712622712
transform 1 0 568 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_312
timestamp 1712622712
transform 1 0 432 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_313
timestamp 1712622712
transform 1 0 576 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_314
timestamp 1712622712
transform 1 0 536 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_315
timestamp 1712622712
transform 1 0 760 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_316
timestamp 1712622712
transform 1 0 560 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_317
timestamp 1712622712
transform 1 0 712 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_318
timestamp 1712622712
transform 1 0 856 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_319
timestamp 1712622712
transform 1 0 776 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_320
timestamp 1712622712
transform 1 0 952 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_321
timestamp 1712622712
transform 1 0 896 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_322
timestamp 1712622712
transform 1 0 3120 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_323
timestamp 1712622712
transform 1 0 2872 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_324
timestamp 1712622712
transform 1 0 3328 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_325
timestamp 1712622712
transform 1 0 3368 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_326
timestamp 1712622712
transform 1 0 3136 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_327
timestamp 1712622712
transform 1 0 3168 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_328
timestamp 1712622712
transform 1 0 3160 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_329
timestamp 1712622712
transform 1 0 3360 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_330
timestamp 1712622712
transform 1 0 3272 0 -1 2370
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1712622712
transform 1 0 1552 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1712622712
transform 1 0 792 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1712622712
transform 1 0 2112 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1712622712
transform 1 0 1488 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1712622712
transform 1 0 1136 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1712622712
transform 1 0 1016 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1712622712
transform 1 0 928 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1712622712
transform 1 0 928 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1712622712
transform 1 0 1088 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1712622712
transform 1 0 1032 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1712622712
transform 1 0 1176 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1712622712
transform 1 0 1288 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1712622712
transform 1 0 1376 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1712622712
transform 1 0 1512 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1712622712
transform 1 0 2024 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1712622712
transform 1 0 1560 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1712622712
transform 1 0 1472 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1712622712
transform 1 0 1864 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1712622712
transform 1 0 1424 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1712622712
transform 1 0 2112 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1712622712
transform 1 0 2392 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1712622712
transform 1 0 2528 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1712622712
transform 1 0 2600 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1712622712
transform 1 0 2704 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1712622712
transform 1 0 2960 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1712622712
transform 1 0 2952 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1712622712
transform 1 0 1176 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1712622712
transform 1 0 3088 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1712622712
transform 1 0 2888 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1712622712
transform 1 0 1232 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1712622712
transform 1 0 3080 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1712622712
transform 1 0 2808 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1712622712
transform 1 0 1560 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1712622712
transform 1 0 2960 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1712622712
transform 1 0 3240 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1712622712
transform 1 0 3280 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_36
timestamp 1712622712
transform 1 0 2776 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_37
timestamp 1712622712
transform 1 0 2992 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_38
timestamp 1712622712
transform 1 0 3112 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1712622712
transform 1 0 3368 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_40
timestamp 1712622712
transform 1 0 3248 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_41
timestamp 1712622712
transform 1 0 3264 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1712622712
transform 1 0 3168 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_43
timestamp 1712622712
transform 1 0 1104 0 1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_44
timestamp 1712622712
transform 1 0 2704 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_45
timestamp 1712622712
transform 1 0 2744 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_46
timestamp 1712622712
transform 1 0 2736 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_47
timestamp 1712622712
transform 1 0 2744 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_48
timestamp 1712622712
transform 1 0 3208 0 1 2570
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1712622712
transform 1 0 3368 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1712622712
transform 1 0 3336 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1712622712
transform 1 0 3248 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1712622712
transform 1 0 2968 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1712622712
transform 1 0 3248 0 -1 1770
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1712622712
transform 1 0 3024 0 -1 2970
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1712622712
transform 1 0 3216 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1712622712
transform 1 0 3304 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_8
timestamp 1712622712
transform 1 0 3168 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_9
timestamp 1712622712
transform 1 0 1696 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_10
timestamp 1712622712
transform 1 0 1240 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_11
timestamp 1712622712
transform 1 0 992 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_12
timestamp 1712622712
transform 1 0 896 0 1 1970
box -8 -3 40 105
use OR2X1  OR2X1_13
timestamp 1712622712
transform 1 0 1312 0 1 1770
box -8 -3 40 105
use OR2X1  OR2X1_14
timestamp 1712622712
transform 1 0 464 0 -1 1570
box -8 -3 40 105
use OR2X1  OR2X1_15
timestamp 1712622712
transform 1 0 496 0 1 1570
box -8 -3 40 105
use OR2X1  OR2X1_16
timestamp 1712622712
transform 1 0 400 0 -1 970
box -8 -3 40 105
use OR2X1  OR2X1_17
timestamp 1712622712
transform 1 0 488 0 1 970
box -8 -3 40 105
use OR2X1  OR2X1_18
timestamp 1712622712
transform 1 0 1248 0 1 370
box -8 -3 40 105
use OR2X1  OR2X1_19
timestamp 1712622712
transform 1 0 2648 0 -1 1370
box -8 -3 40 105
use OR2X1  OR2X1_20
timestamp 1712622712
transform 1 0 3128 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_21
timestamp 1712622712
transform 1 0 3056 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_22
timestamp 1712622712
transform 1 0 3216 0 -1 970
box -8 -3 40 105
use OR2X2  OR2X2_0
timestamp 1712622712
transform 1 0 3376 0 1 770
box -7 -3 35 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1712622712
transform 1 0 3480 0 1 3317
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1712622712
transform 1 0 3480 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1712622712
transform 1 0 24 0 1 3317
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1712622712
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1712622712
transform 1 0 3456 0 1 3293
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1712622712
transform 1 0 3456 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1712622712
transform 1 0 48 0 1 3293
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1712622712
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1712622712
transform 1 0 3480 0 1 3270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1712622712
transform 1 0 3480 0 1 3070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1712622712
transform 1 0 3480 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1712622712
transform 1 0 3480 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1712622712
transform 1 0 3480 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1712622712
transform 1 0 3480 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1712622712
transform 1 0 3480 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1712622712
transform 1 0 3480 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1712622712
transform 1 0 3480 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1712622712
transform 1 0 3480 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1712622712
transform 1 0 3480 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1712622712
transform 1 0 3480 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1712622712
transform 1 0 3480 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1712622712
transform 1 0 3480 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1712622712
transform 1 0 3480 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1712622712
transform 1 0 3480 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1712622712
transform 1 0 3480 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1712622712
transform 1 0 24 0 1 3270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1712622712
transform 1 0 24 0 1 3070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1712622712
transform 1 0 24 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1712622712
transform 1 0 24 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1712622712
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1712622712
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1712622712
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1712622712
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1712622712
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1712622712
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1712622712
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1712622712
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1712622712
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1712622712
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1712622712
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1712622712
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1712622712
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1712622712
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1712622712
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1712622712
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1712622712
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1712622712
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1712622712
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1712622712
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1712622712
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1712622712
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1712622712
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1712622712
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1712622712
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1712622712
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1712622712
transform 1 0 48 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1712622712
transform 1 0 48 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1712622712
transform 1 0 48 0 1 3170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_50
timestamp 1712622712
transform 1 0 3456 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_51
timestamp 1712622712
transform 1 0 3456 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_52
timestamp 1712622712
transform 1 0 3456 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_53
timestamp 1712622712
transform 1 0 3456 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_54
timestamp 1712622712
transform 1 0 3456 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_55
timestamp 1712622712
transform 1 0 3456 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_56
timestamp 1712622712
transform 1 0 3456 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_57
timestamp 1712622712
transform 1 0 3456 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_58
timestamp 1712622712
transform 1 0 3456 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_59
timestamp 1712622712
transform 1 0 3456 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_60
timestamp 1712622712
transform 1 0 3456 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_61
timestamp 1712622712
transform 1 0 3456 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_62
timestamp 1712622712
transform 1 0 3456 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_63
timestamp 1712622712
transform 1 0 3456 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_64
timestamp 1712622712
transform 1 0 3456 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_65
timestamp 1712622712
transform 1 0 3456 0 1 3170
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1712622712
transform 1 0 3032 0 -1 770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1712622712
transform 1 0 3264 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1712622712
transform 1 0 3376 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_3
timestamp 1712622712
transform 1 0 3096 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_4
timestamp 1712622712
transform 1 0 2808 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_5
timestamp 1712622712
transform 1 0 2976 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1712622712
transform 1 0 2824 0 1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1712622712
transform 1 0 2888 0 -1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1712622712
transform 1 0 2784 0 -1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_3
timestamp 1712622712
transform 1 0 2952 0 -1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1712622712
transform 1 0 2992 0 1 3170
box -8 -3 64 105
<< labels >>
rlabel metal2 2876 3338 2876 3338 4 in_clka
rlabel metal2 2004 3338 2004 3338 4 in_clkb
rlabel metal3 3501 1925 3501 1925 4 in_restart
rlabel metal3 3501 795 3501 795 4 in_move[1]
rlabel metal3 3501 815 3501 815 4 in_move[0]
rlabel metal2 956 3338 956 3338 4 board_out[31]
rlabel metal2 884 3338 884 3338 4 board_out[30]
rlabel metal2 700 3338 700 3338 4 board_out[29]
rlabel metal2 636 3338 636 3338 4 board_out[28]
rlabel metal2 604 3338 604 3338 4 board_out[27]
rlabel metal2 564 3338 564 3338 4 board_out[26]
rlabel metal2 580 3338 580 3338 4 board_out[25]
rlabel metal2 620 3338 620 3338 4 board_out[24]
rlabel metal2 780 3338 780 3338 4 board_out[23]
rlabel metal2 748 3338 748 3338 4 board_out[22]
rlabel metal2 916 3338 916 3338 4 board_out[21]
rlabel metal2 1036 3338 1036 3338 4 board_out[20]
rlabel metal2 1052 3338 1052 3338 4 board_out[19]
rlabel metal2 1068 3338 1068 3338 4 board_out[18]
rlabel metal2 1108 3338 1108 3338 4 board_out[17]
rlabel metal2 1188 3338 1188 3338 4 board_out[16]
rlabel metal2 1476 3338 1476 3338 4 board_out[15]
rlabel metal2 1556 3338 1556 3338 4 board_out[14]
rlabel metal2 1636 3338 1636 3338 4 board_out[13]
rlabel metal2 1652 3338 1652 3338 4 board_out[12]
rlabel metal2 1860 3338 1860 3338 4 board_out[11]
rlabel metal2 1940 3338 1940 3338 4 board_out[10]
rlabel metal2 1972 3338 1972 3338 4 board_out[9]
rlabel metal2 1876 3338 1876 3338 4 board_out[8]
rlabel metal2 2292 3338 2292 3338 4 board_out[7]
rlabel metal2 2436 3338 2436 3338 4 board_out[6]
rlabel metal2 2500 3338 2500 3338 4 board_out[5]
rlabel metal2 2452 3338 2452 3338 4 board_out[4]
rlabel metal2 2332 3338 2332 3338 4 board_out[3]
rlabel metal2 2588 3338 2588 3338 4 board_out[2]
rlabel metal2 2484 3338 2484 3338 4 board_out[1]
rlabel metal2 2388 3338 2388 3338 4 board_out[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 28836.002 6345.000 28836.002 6435.000 
<< end >>
