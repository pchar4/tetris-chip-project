magic
tech scmos
timestamp 1710841341
<< metal1 >>
rect 14 2507 2730 2527
rect 38 2483 2706 2503
rect 14 2467 2730 2473
rect 226 2423 236 2426
rect 266 2423 276 2426
rect 1292 2423 1301 2426
rect 1356 2423 1365 2426
rect 226 2416 229 2423
rect 154 2406 157 2414
rect 188 2413 213 2416
rect 220 2413 229 2416
rect 306 2413 316 2416
rect 380 2413 397 2416
rect 500 2413 509 2416
rect 516 2413 525 2416
rect 564 2413 589 2416
rect 620 2413 637 2416
rect 692 2413 717 2416
rect 796 2413 813 2416
rect 908 2413 933 2416
rect 956 2413 981 2416
rect 1076 2413 1085 2416
rect 1132 2413 1157 2416
rect 1188 2413 1213 2416
rect 1236 2413 1245 2416
rect 1290 2413 1333 2416
rect 1354 2413 1389 2416
rect 100 2403 117 2406
rect 154 2403 164 2406
rect 194 2403 212 2406
rect 364 2403 372 2406
rect 506 2405 509 2413
rect 626 2403 644 2406
rect 754 2403 772 2406
rect 930 2405 933 2413
rect 1082 2405 1085 2413
rect 1194 2403 1212 2406
rect 1290 2405 1293 2413
rect 1386 2405 1389 2413
rect 1562 2403 1565 2414
rect 1588 2413 1613 2416
rect 1652 2413 1677 2416
rect 1722 2413 1732 2416
rect 1804 2413 1821 2416
rect 1850 2413 1884 2416
rect 1948 2413 1981 2416
rect 2010 2406 2013 2414
rect 2036 2413 2053 2416
rect 2202 2413 2228 2416
rect 2300 2413 2317 2416
rect 2338 2406 2341 2414
rect 2346 2413 2364 2416
rect 2388 2413 2405 2416
rect 2500 2413 2517 2416
rect 2540 2413 2549 2416
rect 2570 2413 2612 2416
rect 1754 2403 1789 2406
rect 1796 2403 1829 2406
rect 1836 2403 1861 2406
rect 1914 2403 1940 2406
rect 1996 2403 2013 2406
rect 2188 2403 2213 2406
rect 2266 2403 2292 2406
rect 2338 2403 2357 2406
rect 2532 2403 2541 2406
rect 2556 2403 2604 2406
rect 106 2393 140 2396
rect 1754 2395 1757 2403
rect 1762 2393 1788 2396
rect 1946 2393 1988 2396
rect 2266 2393 2284 2396
rect 2306 2393 2324 2396
rect 38 2367 2706 2373
rect 2618 2346 2621 2356
rect 802 2343 837 2346
rect 2108 2343 2156 2346
rect 2618 2343 2636 2346
rect 802 2336 805 2343
rect 146 2333 172 2336
rect 266 2333 284 2336
rect 298 2333 324 2336
rect 338 2333 348 2336
rect 372 2333 397 2336
rect 402 2326 405 2335
rect 428 2333 437 2336
rect 458 2333 484 2336
rect 516 2333 524 2336
rect 796 2333 805 2336
rect 810 2333 844 2336
rect 1066 2333 1084 2336
rect 1172 2333 1189 2336
rect 1242 2333 1260 2336
rect 1340 2333 1365 2336
rect 1546 2333 1564 2336
rect 1580 2333 1605 2336
rect 1626 2333 1652 2336
rect 1722 2333 1740 2336
rect 1754 2333 1772 2336
rect 1778 2333 1820 2336
rect 1884 2333 1924 2336
rect 1242 2326 1245 2333
rect 130 2323 221 2326
rect 130 2313 133 2323
rect 218 2316 221 2323
rect 188 2313 213 2316
rect 218 2313 236 2316
rect 210 2306 213 2313
rect 242 2306 245 2325
rect 292 2323 325 2326
rect 332 2323 349 2326
rect 370 2323 405 2326
rect 426 2323 452 2326
rect 482 2323 492 2326
rect 522 2323 532 2326
rect 692 2323 701 2326
rect 1002 2323 1028 2326
rect 1202 2323 1220 2326
rect 1234 2323 1245 2326
rect 1402 2323 1428 2326
rect 1442 2323 1492 2326
rect 1530 2323 1556 2326
rect 1588 2323 1597 2326
rect 1620 2323 1653 2326
rect 1828 2323 1868 2326
rect 1932 2323 1941 2326
rect 2114 2323 2117 2343
rect 2204 2333 2245 2336
rect 2282 2333 2292 2336
rect 2322 2333 2340 2336
rect 2474 2333 2500 2336
rect 2538 2333 2564 2336
rect 2634 2333 2644 2336
rect 2178 2323 2188 2326
rect 2202 2323 2260 2326
rect 2300 2323 2341 2326
rect 2524 2323 2565 2326
rect 260 2313 277 2316
rect 868 2313 893 2316
rect 1044 2313 1077 2316
rect 1236 2313 1253 2316
rect 1444 2313 1485 2316
rect 1836 2313 1853 2316
rect 1972 2313 1989 2316
rect 210 2303 245 2306
rect 14 2267 2730 2273
rect 234 2233 260 2236
rect 2154 2233 2173 2236
rect 2194 2233 2244 2236
rect 2586 2233 2605 2236
rect 2154 2226 2157 2233
rect 290 2223 308 2226
rect 714 2223 741 2226
rect 714 2216 717 2223
rect 114 2213 124 2216
rect 138 2213 164 2216
rect 338 2213 364 2216
rect 378 2213 388 2216
rect 394 2213 428 2216
rect 452 2213 485 2216
rect 500 2213 509 2216
rect 628 2213 645 2216
rect 100 2203 109 2206
rect 130 2203 156 2206
rect 370 2203 380 2206
rect 444 2203 453 2206
rect 482 2195 485 2213
rect 506 2205 509 2213
rect 642 2196 645 2213
rect 650 2206 653 2216
rect 708 2213 717 2216
rect 722 2213 781 2216
rect 810 2206 813 2225
rect 964 2223 997 2226
rect 1116 2223 1133 2226
rect 1164 2223 1173 2226
rect 1284 2223 1301 2226
rect 1332 2223 1341 2226
rect 1604 2223 1613 2226
rect 1660 2223 1685 2226
rect 1842 2223 1868 2226
rect 1892 2223 1917 2226
rect 1946 2223 1973 2226
rect 2140 2223 2157 2226
rect 930 2213 948 2216
rect 962 2213 1012 2216
rect 1074 2213 1100 2216
rect 1178 2213 1204 2216
rect 1282 2213 1316 2216
rect 1404 2213 1452 2216
rect 1490 2213 1524 2216
rect 1556 2213 1581 2216
rect 1602 2213 1637 2216
rect 1700 2213 1709 2216
rect 1716 2213 1757 2216
rect 1898 2213 1957 2216
rect 1994 2213 2028 2216
rect 2058 2213 2117 2216
rect 2132 2213 2157 2216
rect 2170 2215 2173 2233
rect 2252 2223 2269 2226
rect 2284 2223 2309 2226
rect 2524 2223 2533 2226
rect 2580 2223 2597 2226
rect 2602 2225 2605 2233
rect 2258 2213 2276 2216
rect 2282 2213 2332 2216
rect 2364 2213 2373 2216
rect 2396 2213 2421 2216
rect 2436 2213 2445 2216
rect 2476 2213 2508 2216
rect 2530 2213 2564 2216
rect 650 2203 684 2206
rect 714 2203 748 2206
rect 762 2203 796 2206
rect 810 2203 821 2206
rect 828 2203 869 2206
rect 908 2203 925 2206
rect 930 2203 940 2206
rect 1028 2203 1037 2206
rect 1042 2203 1052 2206
rect 1116 2203 1125 2206
rect 1130 2203 1140 2206
rect 1220 2203 1229 2206
rect 1234 2203 1260 2206
rect 1284 2203 1293 2206
rect 1354 2203 1380 2206
rect 1476 2203 1516 2206
rect 1578 2205 1581 2213
rect 1604 2203 1621 2206
rect 1634 2205 1637 2213
rect 1660 2203 1692 2206
rect 1722 2203 1756 2206
rect 1788 2203 1828 2206
rect 2010 2203 2020 2206
rect 2034 2203 2044 2206
rect 2074 2203 2100 2206
rect 2338 2203 2356 2206
rect 2362 2203 2388 2206
rect 642 2193 677 2196
rect 818 2195 821 2203
rect 1346 2193 1372 2196
rect 1794 2193 1820 2196
rect 2338 2193 2348 2196
rect 2418 2195 2421 2213
rect 2428 2203 2461 2206
rect 2490 2203 2500 2206
rect 2538 2203 2556 2206
rect 2610 2203 2613 2214
rect 38 2167 2706 2173
rect 1114 2143 1132 2146
rect 1450 2143 1460 2146
rect 1612 2143 1637 2146
rect 2018 2143 2044 2146
rect 2218 2143 2228 2146
rect 2314 2143 2332 2146
rect 2506 2143 2524 2146
rect 1634 2136 1637 2143
rect 2218 2136 2221 2143
rect 114 2126 117 2134
rect 138 2133 172 2136
rect 188 2133 205 2136
rect 724 2133 749 2136
rect 780 2133 789 2136
rect 794 2133 804 2136
rect 834 2126 837 2134
rect 858 2133 876 2136
rect 946 2133 964 2136
rect 1130 2133 1140 2136
rect 1234 2133 1244 2136
rect 1266 2133 1308 2136
rect 1380 2133 1389 2136
rect 1394 2133 1420 2136
rect 1436 2133 1477 2136
rect 1514 2133 1524 2136
rect 1548 2133 1589 2136
rect 1634 2133 1644 2136
rect 1668 2133 1685 2136
rect 74 2123 92 2126
rect 106 2123 117 2126
rect 124 2123 164 2126
rect 234 2123 252 2126
rect 338 2106 341 2125
rect 362 2123 372 2126
rect 442 2123 452 2126
rect 516 2123 541 2126
rect 690 2123 700 2126
rect 778 2123 812 2126
rect 826 2123 837 2126
rect 850 2123 884 2126
rect 988 2123 997 2126
rect 1026 2123 1052 2126
rect 1066 2123 1084 2126
rect 1476 2123 1485 2126
rect 1532 2123 1541 2126
rect 1586 2125 1589 2133
rect 1738 2126 1741 2134
rect 1762 2126 1765 2134
rect 1788 2133 1805 2136
rect 1828 2133 1837 2136
rect 1884 2133 1909 2136
rect 1956 2133 1973 2136
rect 2012 2133 2029 2136
rect 2052 2133 2084 2136
rect 2122 2133 2148 2136
rect 2170 2126 2173 2134
rect 2196 2133 2221 2136
rect 2236 2133 2276 2136
rect 2340 2133 2373 2136
rect 2450 2126 2453 2134
rect 2532 2133 2541 2136
rect 2610 2133 2644 2136
rect 1612 2123 1621 2126
rect 1634 2123 1652 2126
rect 1666 2123 1677 2126
rect 388 2113 405 2116
rect 468 2113 477 2116
rect 892 2113 909 2116
rect 940 2113 957 2116
rect 314 2103 341 2106
rect 402 2106 405 2113
rect 1674 2106 1677 2123
rect 1730 2123 1741 2126
rect 1748 2123 1765 2126
rect 1842 2123 1868 2126
rect 1898 2123 1940 2126
rect 2066 2123 2092 2126
rect 2156 2123 2173 2126
rect 2258 2123 2284 2126
rect 2420 2123 2453 2126
rect 2546 2123 2564 2126
rect 2570 2123 2604 2126
rect 1730 2116 1733 2123
rect 1716 2113 1733 2116
rect 2354 2113 2380 2116
rect 402 2103 421 2106
rect 1674 2103 1708 2106
rect 2354 2103 2396 2106
rect 14 2067 2730 2073
rect 1842 2033 1884 2036
rect 2154 2033 2196 2036
rect 100 2023 109 2026
rect 140 2023 157 2026
rect 298 2016 301 2026
rect 1396 2023 1413 2026
rect 1436 2023 1469 2026
rect 1604 2023 1637 2026
rect 1794 2023 1812 2026
rect 1836 2023 1861 2026
rect 1892 2023 1901 2026
rect 2106 2023 2124 2026
rect 2148 2023 2173 2026
rect 2314 2023 2332 2026
rect 2458 2023 2500 2026
rect 2524 2023 2533 2026
rect 1634 2016 1637 2023
rect 202 2013 212 2016
rect 226 2013 244 2016
rect 298 2013 332 2016
rect 436 2013 453 2016
rect 562 2013 588 2016
rect 724 2013 733 2016
rect 764 2013 773 2016
rect 810 2006 813 2014
rect 914 2013 940 2016
rect 946 2013 964 2016
rect 146 2003 172 2006
rect 218 2003 252 2006
rect 266 2003 284 2006
rect 290 2003 324 2006
rect 610 2003 620 2006
rect 644 2003 661 2006
rect 746 2003 756 2006
rect 780 2003 813 2006
rect 946 2003 949 2013
rect 1002 2003 1005 2014
rect 1036 2013 1053 2016
rect 1058 2013 1068 2016
rect 1100 2013 1133 2016
rect 1242 2013 1260 2016
rect 1274 2007 1277 2016
rect 1324 2013 1356 2016
rect 1388 2013 1405 2016
rect 1428 2013 1437 2016
rect 1450 2013 1484 2016
rect 1564 2013 1573 2016
rect 1634 2013 1645 2016
rect 1652 2013 1661 2016
rect 1684 2013 1717 2016
rect 1754 2013 1788 2016
rect 1906 2013 1916 2016
rect 1922 2013 1956 2016
rect 1986 2013 2020 2016
rect 2060 2013 2077 2016
rect 2154 2013 2188 2016
rect 2210 2013 2236 2016
rect 2300 2013 2309 2016
rect 2372 2013 2381 2016
rect 2394 2013 2428 2016
rect 2612 2013 2637 2016
rect 2668 2013 2677 2016
rect 1642 2007 1645 2013
rect 1034 2003 1076 2006
rect 1114 2003 1132 2006
rect 1156 2003 1165 2006
rect 1204 2003 1221 2006
rect 1226 2003 1252 2006
rect 1282 2003 1316 2006
rect 1338 2003 1348 2006
rect 1394 2003 1420 2006
rect 1514 2003 1540 2006
rect 1676 2003 1716 2006
rect 1898 2003 1908 2006
rect 1994 2003 2012 2006
rect 2052 2003 2061 2006
rect 2084 2003 2117 2006
rect 2260 2003 2277 2006
rect 2282 2003 2292 2006
rect 2444 2003 2477 2006
rect 2530 2003 2548 2006
rect 266 1995 269 2003
rect 1218 1996 1221 2003
rect 1218 1993 1245 1996
rect 1282 1993 1308 1996
rect 2058 1993 2076 1996
rect 2242 1993 2252 1996
rect 38 1967 2706 1973
rect 714 1943 724 1946
rect 876 1943 901 1946
rect 1434 1943 1444 1946
rect 1586 1943 1604 1946
rect 1818 1943 1836 1946
rect 1908 1943 1917 1946
rect 2164 1943 2173 1946
rect 2394 1943 2420 1946
rect 146 1933 157 1936
rect 186 1933 196 1936
rect 250 1933 260 1936
rect 674 1933 684 1936
rect 722 1933 732 1936
rect 738 1933 748 1936
rect 778 1933 804 1936
rect 828 1933 837 1936
rect 916 1933 933 1936
rect 1124 1933 1141 1936
rect 1282 1933 1300 1936
rect 1426 1933 1452 1936
rect 1634 1933 1652 1936
rect 1676 1933 1693 1936
rect 1698 1933 1708 1936
rect 1732 1933 1780 1936
rect 1812 1933 1821 1936
rect 1844 1933 1885 1936
rect 2034 1933 2052 1936
rect 2098 1933 2148 1936
rect 2290 1933 2300 1936
rect 2386 1933 2428 1936
rect 2442 1933 2476 1936
rect 2500 1933 2509 1936
rect 74 1923 77 1933
rect 154 1925 157 1933
rect 218 1923 236 1926
rect 250 1923 268 1926
rect 282 1923 300 1926
rect 644 1923 661 1926
rect 700 1923 717 1926
rect 738 1925 741 1933
rect 772 1923 805 1926
rect 834 1923 852 1926
rect 876 1923 885 1926
rect 140 1913 149 1916
rect 218 1915 221 1923
rect 250 1916 253 1923
rect 244 1913 253 1916
rect 828 1913 845 1916
rect 930 1906 933 1933
rect 1146 1926 1149 1933
rect 1130 1923 1149 1926
rect 1170 1926 1173 1933
rect 1170 1923 1181 1926
rect 964 1913 996 1916
rect 1068 1913 1085 1916
rect 1178 1906 1181 1923
rect 1196 1913 1205 1916
rect 1234 1913 1252 1916
rect 1258 1906 1261 1925
rect 1282 1923 1293 1926
rect 1460 1923 1469 1926
rect 1484 1923 1493 1926
rect 1498 1923 1524 1926
rect 1674 1923 1716 1926
rect 1740 1923 1757 1926
rect 1882 1925 1885 1933
rect 2242 1926 2245 1933
rect 2522 1926 2525 1933
rect 1908 1923 1917 1926
rect 2034 1923 2044 1926
rect 2068 1923 2077 1926
rect 2082 1923 2092 1926
rect 2098 1923 2140 1926
rect 2164 1923 2189 1926
rect 2204 1923 2245 1926
rect 2282 1923 2325 1926
rect 2330 1923 2356 1926
rect 2506 1923 2525 1926
rect 2532 1923 2557 1926
rect 2562 1923 2572 1926
rect 2596 1923 2605 1926
rect 1282 1916 1285 1923
rect 1276 1913 1285 1916
rect 1364 1913 1373 1916
rect 1378 1913 1388 1916
rect 1540 1913 1549 1916
rect 1676 1913 1685 1916
rect 2500 1913 2517 1916
rect 2562 1906 2565 1923
rect 930 1903 956 1906
rect 1178 1903 1212 1906
rect 1234 1903 1261 1906
rect 1314 1903 1356 1906
rect 2538 1903 2565 1906
rect 14 1867 2730 1873
rect 538 1833 549 1836
rect 578 1833 612 1836
rect 642 1833 668 1836
rect 690 1833 708 1836
rect 2266 1833 2301 1836
rect 2402 1833 2444 1836
rect 2458 1833 2484 1836
rect 292 1813 301 1816
rect 396 1813 421 1816
rect 458 1813 484 1816
rect 546 1815 549 1833
rect 586 1823 596 1826
rect 626 1823 652 1826
rect 682 1823 692 1826
rect 716 1823 741 1826
rect 1156 1823 1165 1826
rect 1436 1823 1445 1826
rect 1556 1823 1573 1826
rect 2194 1823 2205 1826
rect 2260 1823 2292 1826
rect 2194 1816 2197 1823
rect 722 1813 748 1816
rect 820 1813 837 1816
rect 866 1813 893 1816
rect 930 1813 948 1816
rect 972 1813 1012 1816
rect 1108 1813 1125 1816
rect 1154 1813 1188 1816
rect 1242 1813 1268 1816
rect 1418 1813 1428 1816
rect 1434 1813 1468 1816
rect 1634 1813 1652 1816
rect 1706 1813 1740 1816
rect 1762 1813 1789 1816
rect 1826 1813 1860 1816
rect 1954 1813 1980 1816
rect 2026 1813 2036 1816
rect 2066 1813 2084 1816
rect 2138 1813 2148 1816
rect 2178 1813 2197 1816
rect 2298 1815 2301 1833
rect 2396 1823 2428 1826
rect 2492 1823 2509 1826
rect 2506 1816 2509 1823
rect 2570 1816 2573 1836
rect 2354 1813 2372 1816
rect 2506 1813 2517 1816
rect 2548 1813 2557 1816
rect 2564 1813 2573 1816
rect 2612 1813 2637 1816
rect 2668 1813 2677 1816
rect 794 1803 812 1806
rect 844 1803 885 1806
rect 890 1805 893 1813
rect 938 1803 956 1806
rect 994 1803 1004 1806
rect 1028 1803 1053 1806
rect 1060 1803 1093 1806
rect 1100 1803 1117 1806
rect 1156 1803 1181 1806
rect 1210 1803 1228 1806
rect 1034 1793 1052 1796
rect 1066 1793 1092 1796
rect 1212 1793 1221 1796
rect 1242 1783 1245 1813
rect 1250 1803 1260 1806
rect 1292 1803 1301 1806
rect 1306 1803 1324 1806
rect 1348 1803 1357 1806
rect 1450 1803 1460 1806
rect 1578 1803 1588 1806
rect 1618 1803 1644 1806
rect 1666 1803 1676 1806
rect 1714 1803 1732 1806
rect 1786 1805 1789 1813
rect 1866 1803 1884 1806
rect 1946 1803 1972 1806
rect 2018 1803 2028 1806
rect 2060 1803 2076 1806
rect 2130 1803 2140 1806
rect 2178 1805 2181 1813
rect 2186 1803 2204 1806
rect 2514 1805 2517 1813
rect 2530 1803 2540 1806
rect 1396 1793 1413 1796
rect 1932 1793 1965 1796
rect 38 1767 2706 1773
rect 762 1736 765 1746
rect 978 1743 988 1746
rect 1002 1743 1028 1746
rect 1082 1743 1100 1746
rect 2578 1743 2588 1746
rect 186 1733 196 1736
rect 226 1733 244 1736
rect 364 1733 373 1736
rect 762 1733 796 1736
rect 882 1733 900 1736
rect 914 1733 932 1736
rect 972 1733 989 1736
rect 996 1733 1029 1736
rect 1108 1733 1133 1736
rect 1138 1733 1148 1736
rect 1186 1733 1196 1736
rect 1258 1733 1284 1736
rect 1338 1733 1364 1736
rect 1490 1733 1516 1736
rect 1570 1733 1588 1736
rect 1610 1733 1628 1736
rect 1716 1733 1724 1736
rect 1898 1733 1908 1736
rect 1938 1733 1972 1736
rect 2196 1733 2213 1736
rect 2468 1733 2493 1736
rect 2554 1733 2564 1736
rect 2596 1733 2637 1736
rect 338 1726 341 1733
rect 546 1726 549 1733
rect 842 1726 860 1727
rect 1138 1726 1141 1733
rect 1186 1726 1189 1733
rect 290 1723 341 1726
rect 362 1723 388 1726
rect 476 1723 485 1726
rect 532 1723 549 1726
rect 572 1723 589 1726
rect 748 1723 765 1726
rect 820 1724 860 1726
rect 820 1723 845 1724
rect 908 1723 917 1726
rect 940 1723 965 1726
rect 1068 1723 1101 1726
rect 1122 1723 1141 1726
rect 1156 1723 1189 1726
rect 1258 1723 1292 1726
rect 1298 1723 1324 1726
rect 1330 1723 1372 1726
rect 1388 1723 1405 1726
rect 586 1716 589 1723
rect 586 1713 613 1716
rect 628 1713 645 1716
rect 676 1713 701 1716
rect 706 1706 709 1715
rect 586 1703 620 1706
rect 658 1703 668 1706
rect 682 1703 709 1706
rect 762 1693 765 1723
rect 842 1713 852 1716
rect 876 1713 885 1716
rect 1332 1713 1341 1716
rect 1402 1706 1405 1723
rect 1410 1713 1420 1716
rect 1426 1706 1429 1725
rect 1474 1716 1477 1733
rect 1484 1723 1501 1726
rect 1506 1723 1524 1726
rect 1444 1713 1477 1716
rect 850 1703 868 1706
rect 1394 1703 1429 1706
rect 1538 1703 1541 1733
rect 2122 1726 2125 1733
rect 2410 1726 2413 1733
rect 1596 1723 1621 1726
rect 1666 1723 1700 1726
rect 1722 1723 1732 1726
rect 1812 1723 1821 1726
rect 1898 1723 1916 1726
rect 2012 1723 2029 1726
rect 2092 1723 2125 1726
rect 2154 1723 2180 1726
rect 2218 1723 2228 1726
rect 2260 1723 2269 1726
rect 2300 1723 2325 1726
rect 2410 1723 2437 1726
rect 2444 1723 2453 1726
rect 2490 1723 2516 1726
rect 2572 1723 2589 1726
rect 2634 1725 2637 1733
rect 2660 1723 2677 1726
rect 2218 1716 2221 1723
rect 1746 1713 1772 1716
rect 1818 1713 1860 1716
rect 1884 1713 1893 1716
rect 1932 1713 1949 1716
rect 2196 1713 2221 1716
rect 1746 1693 1749 1713
rect 1826 1703 1876 1706
rect 2018 1703 2068 1706
rect 2450 1703 2453 1723
rect 14 1667 2730 1673
rect 1418 1653 1437 1656
rect 1434 1636 1437 1653
rect 642 1626 645 1636
rect 714 1633 741 1636
rect 548 1623 557 1626
rect 562 1623 580 1626
rect 610 1623 645 1626
rect 706 1623 732 1626
rect 100 1613 133 1616
rect 156 1613 188 1616
rect 244 1613 260 1616
rect 484 1613 493 1616
rect 530 1613 540 1616
rect 618 1613 644 1616
rect 692 1613 725 1616
rect 738 1615 741 1633
rect 1322 1633 1341 1636
rect 1362 1633 1404 1636
rect 1434 1633 1476 1636
rect 1322 1626 1325 1633
rect 756 1623 781 1626
rect 1284 1623 1325 1626
rect 1362 1623 1388 1626
rect 1418 1623 1460 1626
rect 1484 1623 1501 1626
rect 1564 1623 1573 1626
rect 778 1616 781 1623
rect 1498 1616 1501 1623
rect 778 1613 789 1616
rect 828 1613 845 1616
rect 892 1613 940 1616
rect 970 1613 1012 1616
rect 1036 1613 1084 1616
rect 1228 1613 1269 1616
rect 1498 1613 1509 1616
rect 1578 1613 1604 1616
rect 124 1603 132 1606
rect 276 1603 293 1606
rect 498 1603 508 1606
rect 674 1603 684 1606
rect 786 1605 789 1613
rect 850 1603 876 1606
rect 914 1603 932 1606
rect 962 1603 1020 1606
rect 1114 1603 1140 1606
rect 1162 1603 1172 1606
rect 1506 1605 1509 1613
rect 1610 1606 1613 1625
rect 1764 1623 1781 1626
rect 1820 1623 1853 1626
rect 1898 1623 1917 1626
rect 1948 1623 1965 1626
rect 2130 1623 2149 1626
rect 2180 1623 2197 1626
rect 1898 1616 1901 1623
rect 2130 1616 2133 1623
rect 2402 1616 2405 1626
rect 1658 1613 1708 1616
rect 1746 1613 1756 1616
rect 1770 1613 1804 1616
rect 1834 1613 1860 1616
rect 1892 1613 1901 1616
rect 1906 1613 1932 1616
rect 1970 1613 1996 1616
rect 2082 1613 2108 1616
rect 2122 1613 2133 1616
rect 1538 1603 1548 1606
rect 1570 1603 1595 1606
rect 1610 1603 1644 1606
rect 1690 1603 1700 1606
rect 1724 1603 1741 1606
rect 1762 1603 1796 1606
rect 1826 1603 1868 1606
rect 1884 1603 1893 1606
rect 1906 1603 1924 1606
rect 1948 1603 1973 1606
rect 2020 1603 2037 1606
rect 2122 1605 2125 1613
rect 2234 1606 2237 1614
rect 2242 1613 2276 1616
rect 2314 1613 2356 1616
rect 2370 1613 2405 1616
rect 2444 1613 2485 1616
rect 2522 1613 2548 1616
rect 2612 1613 2637 1616
rect 2138 1603 2156 1606
rect 2234 1603 2268 1606
rect 2300 1603 2341 1606
rect 2370 1605 2373 1613
rect 2378 1603 2412 1606
rect 2450 1603 2484 1606
rect 490 1593 500 1596
rect 828 1593 837 1596
rect 892 1593 925 1596
rect 1036 1593 1053 1596
rect 2202 1593 2220 1596
rect 1050 1583 1053 1593
rect 2074 1583 2093 1586
rect 38 1567 2706 1573
rect 1362 1553 1373 1556
rect 218 1543 228 1546
rect 802 1536 805 1546
rect 810 1543 820 1546
rect 834 1543 860 1546
rect 954 1543 980 1546
rect 994 1543 1029 1546
rect 1026 1536 1029 1543
rect 218 1533 236 1536
rect 466 1533 476 1536
rect 506 1533 548 1536
rect 578 1533 588 1536
rect 642 1533 660 1536
rect 714 1533 724 1536
rect 802 1533 828 1536
rect 858 1533 868 1536
rect 890 1533 916 1536
rect 988 1533 1021 1536
rect 1026 1533 1036 1536
rect 1082 1533 1116 1536
rect 1170 1533 1188 1536
rect 1250 1533 1260 1536
rect 1282 1533 1300 1536
rect 1362 1526 1365 1546
rect 156 1523 181 1526
rect 212 1523 229 1526
rect 244 1523 253 1526
rect 572 1523 589 1526
rect 628 1523 661 1526
rect 700 1523 725 1526
rect 890 1523 924 1526
rect 1002 1523 1044 1526
rect 1074 1523 1124 1526
rect 1162 1523 1196 1526
rect 1242 1523 1268 1526
rect 1308 1523 1349 1526
rect 1356 1523 1365 1526
rect 1370 1516 1373 1553
rect 1874 1543 1900 1546
rect 2418 1536 2421 1556
rect 2482 1543 2492 1546
rect 1506 1526 1509 1534
rect 1530 1533 1540 1536
rect 1570 1533 1588 1536
rect 1602 1533 1636 1536
rect 1650 1533 1676 1536
rect 1706 1533 1724 1536
rect 1738 1533 1772 1536
rect 1786 1533 1804 1536
rect 1362 1513 1380 1516
rect 1404 1513 1429 1516
rect 1458 1506 1461 1525
rect 1498 1523 1509 1526
rect 1548 1523 1565 1526
rect 1498 1516 1501 1523
rect 1476 1513 1501 1516
rect 1602 1515 1605 1533
rect 1842 1526 1845 1534
rect 1868 1533 1901 1536
rect 1908 1533 1917 1536
rect 1922 1533 1940 1536
rect 2034 1533 2044 1536
rect 2066 1533 2092 1536
rect 2314 1526 2317 1534
rect 2322 1533 2348 1536
rect 2418 1533 2428 1536
rect 2460 1533 2469 1536
rect 2500 1533 2525 1536
rect 2546 1533 2564 1536
rect 2588 1533 2637 1536
rect 1644 1523 1677 1526
rect 1684 1523 1717 1526
rect 1732 1523 1773 1526
rect 1780 1523 1805 1526
rect 1812 1523 1845 1526
rect 1948 1523 1957 1526
rect 2010 1523 2036 1526
rect 2132 1523 2149 1526
rect 2260 1523 2285 1526
rect 2314 1523 2349 1526
rect 2404 1523 2421 1526
rect 2514 1523 2540 1526
rect 2572 1523 2581 1526
rect 2634 1525 2637 1533
rect 2660 1523 2669 1526
rect 1740 1513 1749 1516
rect 1868 1513 1893 1516
rect 1956 1513 1965 1516
rect 1970 1513 1980 1516
rect 2146 1513 2156 1516
rect 2180 1513 2213 1516
rect 2316 1513 2333 1516
rect 1418 1503 1461 1506
rect 1962 1503 1996 1506
rect 2138 1503 2172 1506
rect 14 1467 2730 1473
rect 866 1433 901 1436
rect 1330 1433 1357 1436
rect 1386 1433 1428 1436
rect 1938 1433 1964 1436
rect 524 1423 533 1426
rect 724 1423 765 1426
rect 780 1423 789 1426
rect 786 1416 789 1423
rect 108 1413 133 1416
rect 164 1413 205 1416
rect 220 1413 229 1416
rect 394 1413 436 1416
rect 466 1413 509 1416
rect 516 1413 533 1416
rect 596 1413 613 1416
rect 170 1403 212 1406
rect 218 1403 228 1406
rect 276 1403 301 1406
rect 506 1405 509 1413
rect 562 1403 588 1406
rect 602 1403 628 1406
rect 634 1403 637 1414
rect 786 1413 797 1416
rect 860 1413 877 1416
rect 898 1415 901 1433
rect 916 1423 925 1426
rect 1276 1423 1293 1426
rect 650 1403 668 1406
rect 682 1403 700 1406
rect 738 1403 764 1406
rect 794 1405 797 1413
rect 922 1406 925 1423
rect 930 1413 980 1416
rect 1010 1413 1060 1416
rect 1242 1413 1300 1416
rect 1354 1415 1357 1433
rect 1378 1423 1412 1426
rect 1436 1423 1461 1426
rect 1506 1423 1517 1426
rect 1684 1423 1701 1426
rect 1732 1423 1749 1426
rect 1884 1423 1901 1426
rect 1948 1423 1957 1426
rect 1972 1423 1989 1426
rect 2172 1423 2189 1426
rect 1506 1416 1509 1423
rect 1378 1413 1420 1416
rect 1492 1413 1509 1416
rect 1540 1413 1549 1416
rect 1554 1413 1572 1416
rect 1604 1413 1621 1416
rect 1628 1413 1661 1416
rect 1676 1413 1717 1416
rect 1724 1413 1757 1416
rect 1778 1406 1781 1416
rect 1802 1413 1812 1416
rect 1834 1413 1868 1416
rect 1924 1413 1933 1416
rect 2004 1413 2021 1416
rect 2090 1413 2100 1416
rect 2130 1413 2156 1416
rect 2170 1413 2204 1416
rect 2282 1413 2292 1416
rect 2372 1413 2381 1416
rect 2460 1413 2469 1416
rect 2476 1413 2485 1416
rect 810 1403 852 1406
rect 922 1403 972 1406
rect 1132 1403 1173 1406
rect 1188 1403 1205 1406
rect 1498 1403 1516 1406
rect 1610 1403 1619 1406
rect 1642 1403 1668 1406
rect 1706 1403 1716 1406
rect 1746 1403 1764 1406
rect 1770 1403 1804 1406
rect 1828 1403 1845 1406
rect 1850 1403 1860 1406
rect 1884 1403 1893 1406
rect 1986 1403 1996 1406
rect 2058 1403 2092 1406
rect 2172 1403 2189 1406
rect 2252 1403 2284 1406
rect 2378 1405 2381 1413
rect 2522 1406 2525 1414
rect 2548 1413 2557 1416
rect 2412 1403 2421 1406
rect 2492 1403 2525 1406
rect 594 1393 620 1396
rect 1098 1393 1124 1396
rect 2226 1393 2244 1396
rect 2434 1393 2444 1396
rect 38 1367 2706 1373
rect 2090 1336 2093 1346
rect 226 1333 244 1336
rect 258 1333 276 1336
rect 290 1333 309 1336
rect 356 1333 365 1336
rect 428 1333 437 1336
rect 746 1334 764 1336
rect 746 1333 765 1334
rect 842 1333 852 1336
rect 866 1333 884 1336
rect 930 1333 948 1336
rect 954 1333 988 1336
rect 108 1323 125 1326
rect 220 1323 245 1326
rect 290 1325 293 1333
rect 762 1326 765 1333
rect 1034 1326 1037 1334
rect 1050 1333 1068 1336
rect 1090 1333 1108 1336
rect 1426 1333 1452 1336
rect 1466 1333 1492 1336
rect 1610 1326 1613 1334
rect 1682 1326 1685 1334
rect 1698 1333 1740 1336
rect 1764 1333 1773 1336
rect 1794 1326 1797 1334
rect 1818 1333 1852 1336
rect 1876 1333 1893 1336
rect 2012 1333 2029 1336
rect 2034 1333 2044 1336
rect 2090 1333 2116 1336
rect 2156 1333 2165 1336
rect 298 1323 324 1326
rect 364 1323 397 1326
rect 522 1323 532 1326
rect 612 1323 629 1326
rect 714 1323 765 1326
rect 804 1323 829 1326
rect 962 1323 1037 1326
rect 1044 1323 1069 1326
rect 1076 1323 1101 1326
rect 1116 1323 1133 1326
rect 1178 1323 1204 1326
rect 1260 1323 1300 1326
rect 1346 1323 1372 1326
rect 1410 1323 1437 1326
rect 1490 1323 1500 1326
rect 1602 1323 1613 1326
rect 1620 1323 1668 1326
rect 1682 1323 1748 1326
rect 1762 1323 1797 1326
rect 1804 1323 1837 1326
rect 1842 1323 1860 1326
rect 1986 1323 1996 1326
rect 2026 1323 2052 1326
rect 2162 1323 2212 1326
rect 716 1313 725 1316
rect 826 1303 829 1323
rect 1602 1316 1605 1323
rect 2218 1316 2221 1346
rect 2282 1323 2308 1326
rect 2322 1325 2325 1356
rect 2346 1333 2396 1336
rect 2532 1333 2541 1336
rect 2530 1323 2620 1326
rect 1514 1313 1548 1316
rect 1572 1313 1605 1316
rect 1684 1313 1733 1316
rect 1764 1313 1781 1316
rect 1876 1313 1901 1316
rect 2218 1313 2228 1316
rect 2252 1313 2261 1316
rect 1538 1303 1564 1306
rect 2218 1303 2244 1306
rect 14 1267 2730 1273
rect 1338 1226 1341 1246
rect 1354 1233 1404 1236
rect 1682 1233 1724 1236
rect 1874 1233 1893 1236
rect 228 1223 269 1226
rect 562 1223 573 1226
rect 716 1223 741 1226
rect 890 1223 909 1226
rect 948 1223 965 1226
rect 988 1223 1029 1226
rect 1052 1223 1093 1226
rect 1108 1223 1125 1226
rect 1156 1223 1197 1226
rect 1338 1223 1388 1226
rect 1412 1223 1453 1226
rect 1516 1223 1565 1226
rect 562 1216 565 1223
rect 1026 1216 1029 1223
rect 1562 1216 1565 1223
rect 1682 1223 1708 1226
rect 1868 1223 1877 1226
rect 2108 1223 2141 1226
rect 2308 1223 2341 1226
rect 1682 1216 1685 1223
rect 2130 1216 2133 1223
rect 380 1213 389 1216
rect 442 1213 452 1216
rect 532 1213 565 1216
rect 620 1213 685 1216
rect 884 1213 940 1216
rect 954 1213 980 1216
rect 1026 1213 1044 1216
rect 1058 1213 1100 1216
rect 1106 1213 1148 1216
rect 1212 1213 1261 1216
rect 1268 1213 1293 1216
rect 1508 1213 1557 1216
rect 1562 1213 1573 1216
rect 1652 1213 1685 1216
rect 1778 1213 1788 1216
rect 1794 1213 1829 1216
rect 1860 1213 1901 1216
rect 1956 1213 1965 1216
rect 2050 1213 2092 1216
rect 2130 1213 2148 1216
rect 2180 1213 2189 1216
rect 2220 1213 2245 1216
rect 2252 1213 2292 1216
rect 2314 1213 2348 1216
rect 2444 1213 2453 1216
rect 250 1203 284 1206
rect 300 1203 357 1206
rect 458 1203 508 1206
rect 524 1203 549 1206
rect 554 1203 572 1206
rect 612 1203 645 1206
rect 762 1203 780 1206
rect 804 1203 813 1206
rect 842 1203 860 1206
rect 876 1203 893 1206
rect 914 1203 932 1206
rect 954 1203 972 1206
rect 1026 1203 1036 1206
rect 1106 1203 1140 1206
rect 1186 1203 1204 1206
rect 1226 1203 1260 1206
rect 1290 1203 1316 1206
rect 1570 1205 1573 1213
rect 1602 1203 1644 1206
rect 1666 1203 1693 1206
rect 1746 1203 1780 1206
rect 1826 1203 1852 1206
rect 1908 1203 1941 1206
rect 1980 1203 2021 1206
rect 2050 1205 2053 1213
rect 2066 1203 2084 1206
rect 2108 1203 2149 1206
rect 2178 1203 2196 1206
rect 2226 1203 2244 1206
rect 2308 1203 2333 1206
rect 2394 1203 2420 1206
rect 2524 1203 2548 1206
rect 380 1193 405 1196
rect 1026 1183 1029 1203
rect 38 1167 2706 1173
rect 170 1136 173 1145
rect 330 1143 348 1146
rect 1410 1143 1428 1146
rect 82 1133 92 1136
rect 148 1133 173 1136
rect 218 1133 252 1136
rect 276 1133 285 1136
rect 316 1133 325 1136
rect 330 1133 356 1136
rect 482 1133 508 1136
rect 618 1133 628 1136
rect 652 1133 661 1136
rect 682 1133 692 1136
rect 716 1133 725 1136
rect 938 1133 980 1136
rect 1282 1133 1324 1136
rect 1362 1126 1365 1134
rect 1458 1133 1476 1136
rect 1522 1133 1532 1136
rect 1562 1133 1588 1136
rect 1610 1126 1613 1134
rect 1618 1133 1660 1136
rect 1698 1133 1716 1136
rect 1738 1133 1764 1136
rect 1778 1133 1828 1136
rect 1898 1126 1901 1145
rect 1914 1143 1948 1146
rect 2018 1136 2021 1146
rect 2052 1143 2069 1146
rect 2090 1143 2101 1146
rect 1956 1133 1973 1136
rect 1986 1133 2004 1136
rect 2018 1133 2036 1136
rect 2098 1126 2101 1143
rect 2122 1133 2132 1136
rect 2146 1133 2188 1136
rect 2242 1133 2268 1136
rect 2450 1126 2453 1136
rect 2482 1133 2500 1136
rect 2562 1133 2572 1136
rect 2596 1133 2613 1136
rect 2634 1133 2652 1136
rect 66 1123 100 1126
rect 114 1123 124 1126
rect 156 1123 165 1126
rect 372 1123 381 1126
rect 428 1123 452 1126
rect 490 1123 516 1126
rect 522 1123 556 1126
rect 572 1123 589 1126
rect 626 1123 636 1126
rect 714 1123 772 1126
rect 962 1123 988 1126
rect 1026 1123 1036 1126
rect 1050 1123 1100 1126
rect 1170 1123 1220 1126
rect 1226 1123 1276 1126
rect 1314 1123 1365 1126
rect 1372 1123 1381 1126
rect 1444 1123 1477 1126
rect 1490 1123 1540 1126
rect 1610 1123 1629 1126
rect 1668 1123 1693 1126
rect 1706 1123 1724 1126
rect 1746 1123 1772 1126
rect 1826 1123 1836 1126
rect 1860 1123 1901 1126
rect 1916 1123 1933 1126
rect 1978 1123 2012 1126
rect 2098 1123 2109 1126
rect 2140 1123 2180 1126
rect 2292 1123 2317 1126
rect 1314 1116 1317 1123
rect 276 1113 285 1116
rect 316 1113 325 1116
rect 652 1113 661 1116
rect 882 1113 908 1116
rect 932 1113 981 1116
rect 996 1113 1013 1116
rect 1044 1113 1061 1116
rect 1228 1113 1237 1116
rect 1284 1113 1317 1116
rect 1380 1113 1405 1116
rect 1548 1113 1581 1116
rect 1676 1113 1685 1116
rect 834 1103 860 1106
rect 874 1103 924 1106
rect 1706 1103 1709 1123
rect 1978 1083 1981 1123
rect 2124 1113 2133 1116
rect 2148 1113 2165 1116
rect 2314 1113 2324 1116
rect 2330 1106 2333 1125
rect 2354 1123 2380 1126
rect 2402 1113 2420 1116
rect 2426 1106 2429 1125
rect 2450 1123 2468 1126
rect 2530 1123 2540 1126
rect 2602 1123 2628 1126
rect 2660 1123 2669 1126
rect 2444 1113 2453 1116
rect 2298 1103 2333 1106
rect 2394 1103 2429 1106
rect 14 1067 2730 1073
rect 626 1033 652 1036
rect 874 1033 893 1036
rect 2314 1033 2348 1036
rect 2618 1033 2652 1036
rect 260 1023 269 1026
rect 874 1016 877 1033
rect 1252 1023 1285 1026
rect 1548 1023 1565 1026
rect 2122 1023 2140 1026
rect 2164 1023 2181 1026
rect 2178 1016 2181 1023
rect 2322 1023 2341 1026
rect 2356 1023 2365 1026
rect 2612 1023 2629 1026
rect 2322 1016 2325 1023
rect 212 1013 244 1016
rect 316 1013 341 1016
rect 372 1013 397 1016
rect 428 1013 445 1016
rect 506 1013 524 1016
rect 554 1013 564 1016
rect 620 1013 629 1016
rect 762 1013 804 1016
rect 836 1013 877 1016
rect 988 1013 997 1016
rect 1082 1013 1108 1016
rect 1218 1013 1244 1016
rect 1378 1013 1405 1016
rect 1466 1013 1476 1016
rect 1540 1013 1565 1016
rect 1604 1013 1621 1016
rect 1660 1013 1685 1016
rect 1756 1013 1789 1016
rect 1826 1013 1868 1016
rect 2010 1013 2036 1016
rect 2108 1013 2125 1016
rect 2178 1013 2188 1016
rect 2220 1013 2252 1016
rect 2300 1013 2325 1016
rect 2362 1016 2365 1023
rect 2362 1013 2373 1016
rect 2380 1013 2397 1016
rect 2402 1013 2412 1016
rect 2442 1013 2476 1016
rect 2532 1013 2541 1016
rect 2562 1013 2596 1016
rect 394 1006 397 1013
rect 394 1003 412 1006
rect 442 1005 445 1013
rect 1378 1006 1381 1013
rect 468 1003 485 1006
rect 724 1003 741 1006
rect 748 1003 757 1006
rect 778 1003 812 1006
rect 914 1003 957 1006
rect 980 1003 1005 1006
rect 1010 1003 1036 1006
rect 1060 1003 1069 1006
rect 1074 1003 1100 1006
rect 1124 1003 1133 1006
rect 1210 1003 1236 1006
rect 1258 1003 1308 1006
rect 1356 1003 1381 1006
rect 1386 1003 1420 1006
rect 1450 1003 1468 1006
rect 1522 1003 1532 1006
rect 1610 1003 1652 1006
rect 1666 1003 1700 1006
rect 1762 1003 1788 1006
rect 1826 1003 1860 1006
rect 1884 1003 1941 1006
rect 1980 1003 1997 1006
rect 2018 1003 2028 1006
rect 2060 1003 2077 1006
rect 2170 1003 2196 1006
rect 2218 1003 2244 1006
rect 2266 1003 2276 1006
rect 738 995 741 1003
rect 1074 996 1077 1003
rect 1066 993 1077 996
rect 1290 993 1300 996
rect 1338 993 1348 996
rect 1370 993 1412 996
rect 1890 993 1948 996
rect 1962 993 1972 996
rect 1994 986 1997 1003
rect 2108 993 2117 996
rect 2306 993 2309 1013
rect 2370 1005 2373 1013
rect 2442 1003 2461 1006
rect 2506 1003 2524 1006
rect 2548 1003 2557 1006
rect 2562 1003 2588 1006
rect 1994 983 2013 986
rect 38 967 2706 973
rect 282 943 340 946
rect 466 936 469 956
rect 2074 953 2109 956
rect 772 943 781 946
rect 1786 943 1820 946
rect 1938 943 1964 946
rect 2346 943 2364 946
rect 2420 943 2437 946
rect 2626 943 2644 946
rect 348 933 389 936
rect 420 933 469 936
rect 474 926 477 934
rect 586 926 589 934
rect 92 923 109 926
rect 148 923 165 926
rect 244 923 253 926
rect 260 923 285 926
rect 356 923 381 926
rect 404 923 413 926
rect 428 923 477 926
rect 516 923 549 926
rect 586 923 597 926
rect 634 923 685 926
rect 282 913 285 923
rect 594 906 597 923
rect 708 913 741 916
rect 778 913 781 943
rect 2346 936 2349 943
rect 786 933 796 936
rect 826 933 852 936
rect 1010 933 1028 936
rect 1052 933 1061 936
rect 1066 933 1092 936
rect 1170 933 1196 936
rect 1242 933 1284 936
rect 1316 933 1341 936
rect 1346 926 1349 934
rect 1402 933 1420 936
rect 860 923 877 926
rect 916 923 933 926
rect 994 923 1004 926
rect 1066 923 1085 926
rect 1220 923 1229 926
rect 1236 923 1269 926
rect 1282 923 1292 926
rect 1330 923 1349 926
rect 1442 926 1445 934
rect 1450 933 1476 936
rect 1500 933 1517 936
rect 1522 933 1532 936
rect 1610 933 1629 936
rect 1442 923 1477 926
rect 1514 923 1540 926
rect 1610 923 1613 933
rect 1634 926 1637 934
rect 1660 933 1693 936
rect 1930 933 1972 936
rect 1618 923 1637 926
rect 1690 927 1693 933
rect 1690 924 1708 927
rect 2034 926 2037 934
rect 2068 933 2101 936
rect 2172 933 2213 936
rect 2258 933 2276 936
rect 2324 933 2349 936
rect 2378 933 2397 936
rect 2618 933 2652 936
rect 1836 923 1845 926
rect 1852 923 1877 926
rect 1882 923 1900 926
rect 1994 923 2037 926
rect 2124 923 2149 926
rect 2284 923 2301 926
rect 2394 925 2397 933
rect 2420 923 2429 926
rect 2476 923 2485 926
rect 2594 923 2612 926
rect 2660 923 2677 926
rect 868 913 885 916
rect 1052 913 1085 916
rect 1130 913 1140 916
rect 1164 913 1197 916
rect 1596 913 1629 916
rect 1682 913 1700 916
rect 1724 913 1749 916
rect 1780 913 1789 916
rect 2132 913 2141 916
rect 2324 913 2349 916
rect 2538 913 2556 916
rect 594 903 620 906
rect 1698 903 1716 906
rect 1754 903 1772 906
rect 2562 903 2572 906
rect 14 867 2730 873
rect 2258 833 2277 836
rect 2258 826 2261 833
rect 140 823 149 826
rect 220 823 245 826
rect 276 823 285 826
rect 330 823 349 826
rect 748 823 757 826
rect 820 823 845 826
rect 980 823 1005 826
rect 330 816 333 823
rect 1034 816 1037 825
rect 1042 823 1067 826
rect 1092 823 1117 826
rect 1180 823 1197 826
rect 1756 823 1765 826
rect 2140 823 2165 826
rect 2236 823 2261 826
rect 66 813 92 816
rect 114 813 124 816
rect 194 813 204 816
rect 324 813 333 816
rect 338 813 356 816
rect 410 813 420 816
rect 476 813 485 816
rect 532 813 541 816
rect 612 813 629 816
rect 722 813 740 816
rect 762 813 788 816
rect 812 813 852 816
rect 932 813 957 816
rect 994 813 1020 816
rect 1034 813 1053 816
rect 1098 813 1132 816
rect 1228 813 1237 816
rect 1308 813 1349 816
rect 1402 813 1420 816
rect 1482 813 1500 816
rect 1570 813 1621 816
rect 1658 813 1692 816
rect 1706 813 1740 816
rect 338 806 341 813
rect 108 803 116 806
rect 162 803 180 806
rect 186 803 196 806
rect 220 803 229 806
rect 242 803 252 806
rect 276 803 300 806
rect 316 803 341 806
rect 362 803 372 806
rect 386 803 412 806
rect 468 803 493 806
rect 498 803 524 806
rect 666 803 700 806
rect 714 803 732 806
rect 882 803 924 806
rect 938 803 956 806
rect 994 803 1012 806
rect 1180 803 1189 806
rect 1202 803 1220 806
rect 1258 803 1300 806
rect 1314 803 1365 806
rect 1378 803 1428 806
rect 1522 803 1532 806
rect 1786 805 1789 816
rect 1796 813 1821 816
rect 1836 813 1845 816
rect 1874 806 1877 815
rect 1900 813 1909 816
rect 1978 813 1988 816
rect 2002 813 2045 816
rect 2082 813 2124 816
rect 2218 813 2228 816
rect 2274 815 2277 833
rect 2292 823 2317 826
rect 2540 823 2557 826
rect 2314 816 2317 823
rect 2314 813 2325 816
rect 2332 813 2341 816
rect 2346 813 2364 816
rect 2428 813 2445 816
rect 2476 813 2517 816
rect 2538 813 2565 816
rect 2572 813 2613 816
rect 1828 803 1877 806
rect 1948 803 1973 806
rect 2002 805 2005 813
rect 2034 803 2044 806
rect 2090 803 2116 806
rect 2146 803 2164 806
rect 2322 805 2325 813
rect 2338 803 2356 806
rect 2370 803 2412 806
rect 2468 803 2509 806
rect 2562 805 2565 813
rect 2602 803 2620 806
rect 2652 803 2669 806
rect 682 793 692 796
rect 1338 793 1348 796
rect 1922 793 1940 796
rect 38 767 2706 773
rect 146 743 164 746
rect 146 736 149 743
rect 116 733 149 736
rect 258 733 268 736
rect 434 733 452 736
rect 498 733 508 736
rect 642 733 684 736
rect 700 733 725 736
rect 738 733 748 736
rect 772 733 781 736
rect 434 726 437 733
rect 124 723 157 726
rect 250 723 276 726
rect 364 723 389 726
rect 420 723 437 726
rect 468 723 485 726
rect 490 723 500 726
rect 586 723 612 726
rect 628 723 669 726
rect 714 723 756 726
rect 250 713 253 723
rect 786 716 789 756
rect 978 743 988 746
rect 1074 743 1108 746
rect 1666 743 1700 746
rect 2122 743 2132 746
rect 2458 743 2476 746
rect 866 726 869 734
rect 996 733 1052 736
rect 1116 733 1141 736
rect 1162 733 1204 736
rect 1242 733 1284 736
rect 1306 733 1316 736
rect 1418 733 1444 736
rect 1474 733 1492 736
rect 1554 733 1572 736
rect 1604 733 1629 736
rect 1660 733 1693 736
rect 1698 733 1708 736
rect 1740 733 1765 736
rect 1698 726 1701 733
rect 1786 726 1789 734
rect 1820 733 1829 736
rect 1938 733 1956 736
rect 2004 733 2037 736
rect 1938 726 1941 733
rect 2042 726 2045 734
rect 2100 733 2109 736
rect 2114 733 2140 736
rect 2146 733 2156 736
rect 2346 733 2372 736
rect 2410 733 2436 736
rect 2484 733 2516 736
rect 2548 733 2557 736
rect 2634 733 2652 736
rect 2106 726 2109 733
rect 858 723 869 726
rect 876 723 893 726
rect 922 723 956 726
rect 1130 723 1156 726
rect 1162 723 1212 726
rect 1298 723 1324 726
rect 1330 723 1348 726
rect 1474 723 1500 726
rect 1532 723 1573 726
rect 1618 723 1644 726
rect 1658 723 1701 726
rect 1716 723 1725 726
rect 1748 723 1789 726
rect 1876 723 1901 726
rect 1932 723 1941 726
rect 1972 723 1981 726
rect 2018 723 2045 726
rect 2052 723 2069 726
rect 2106 723 2125 726
rect 2340 723 2373 726
rect 2506 723 2524 726
rect 2578 723 2588 726
rect 2612 723 2621 726
rect 858 716 861 723
rect 292 713 301 716
rect 772 713 789 716
rect 836 713 861 716
rect 916 713 949 716
rect 2170 713 2196 716
rect 2220 713 2237 716
rect 2242 706 2245 715
rect 2274 713 2300 716
rect 818 703 828 706
rect 2170 703 2212 706
rect 2226 703 2245 706
rect 2250 703 2260 706
rect 2282 703 2316 706
rect 14 667 2730 673
rect 1282 633 1316 636
rect 348 623 365 626
rect 426 623 444 626
rect 604 623 613 626
rect 1234 623 1252 626
rect 1282 623 1300 626
rect 1492 623 1509 626
rect 2218 623 2229 626
rect 2218 616 2221 623
rect 2274 616 2277 636
rect 124 613 141 616
rect 146 613 172 616
rect 186 613 196 616
rect 202 613 245 616
rect 300 613 333 616
rect 346 613 380 616
rect 386 613 420 616
rect 482 613 516 616
rect 548 613 557 616
rect 602 613 628 616
rect 684 613 709 616
rect 740 613 757 616
rect 802 613 820 616
rect 826 613 860 616
rect 1012 613 1037 616
rect 1068 613 1093 616
rect 1140 613 1149 616
rect 1180 613 1205 616
rect 1220 613 1245 616
rect 1388 613 1428 616
rect 1442 613 1476 616
rect 1546 613 1572 616
rect 1618 613 1644 616
rect 1650 613 1684 616
rect 1756 613 1773 616
rect 1802 613 1837 616
rect 1874 613 1908 616
rect 1996 613 2005 616
rect 2028 613 2045 616
rect 2058 613 2076 616
rect 2130 613 2148 616
rect 2172 613 2189 616
rect 2204 613 2221 616
rect 2252 613 2277 616
rect 116 603 157 606
rect 210 603 244 606
rect 274 603 292 606
rect 330 605 333 613
rect 754 606 757 613
rect 1090 606 1093 613
rect 362 603 372 606
rect 386 603 412 606
rect 490 603 508 606
rect 570 603 580 606
rect 754 603 772 606
rect 802 603 812 606
rect 884 603 924 606
rect 1090 603 1108 606
rect 1122 603 1132 606
rect 1242 603 1245 613
rect 1354 603 1372 606
rect 1442 605 1445 613
rect 1498 603 1532 606
rect 1538 603 1580 606
rect 1596 603 1636 606
rect 1666 603 1676 606
rect 1700 603 1717 606
rect 1722 603 1732 606
rect 1804 603 1821 606
rect 1834 605 1837 613
rect 1882 603 1900 606
rect 1924 603 1948 606
rect 1970 603 1988 606
rect 2218 603 2228 606
rect 2274 605 2277 613
rect 2322 606 2325 616
rect 2338 613 2356 616
rect 2380 613 2397 616
rect 2444 613 2469 616
rect 2500 613 2509 616
rect 2514 613 2532 616
rect 2612 613 2621 616
rect 2298 605 2325 606
rect 2298 603 2324 605
rect 788 593 797 596
rect 38 567 2706 573
rect 434 543 444 546
rect 234 533 252 536
rect 452 533 484 536
rect 522 526 525 534
rect 578 533 604 536
rect 756 533 773 536
rect 66 523 100 526
rect 164 523 181 526
rect 186 523 212 526
rect 316 523 325 526
rect 508 523 525 526
rect 628 523 669 526
rect 706 523 732 526
rect 764 523 773 526
rect 794 523 804 526
rect 842 523 860 526
rect 890 523 916 526
rect 922 523 957 526
rect 1044 523 1053 526
rect 1066 525 1069 546
rect 1410 543 1420 546
rect 2474 543 2524 546
rect 1162 533 1180 536
rect 1194 533 1204 536
rect 1236 533 1245 536
rect 1250 533 1276 536
rect 1282 533 1293 536
rect 1314 533 1324 536
rect 1250 526 1253 533
rect 1194 523 1212 526
rect 1242 523 1253 526
rect 1290 526 1293 533
rect 1362 526 1365 534
rect 1396 533 1428 536
rect 1492 533 1501 536
rect 1506 533 1540 536
rect 1554 533 1564 536
rect 1644 533 1653 536
rect 1778 533 1804 536
rect 1882 533 1908 536
rect 1988 533 2013 536
rect 2074 526 2077 534
rect 2108 533 2117 536
rect 2122 533 2156 536
rect 2306 533 2316 536
rect 2338 533 2380 536
rect 2532 533 2549 536
rect 2578 533 2628 536
rect 1290 523 1308 526
rect 1332 523 1365 526
rect 1522 523 1548 526
rect 1554 523 1572 526
rect 1668 523 1677 526
rect 116 513 125 516
rect 228 513 245 516
rect 636 513 661 516
rect 666 513 676 516
rect 1060 513 1069 516
rect 1090 513 1116 516
rect 658 506 661 513
rect 378 503 412 506
rect 658 503 692 506
rect 1058 503 1076 506
rect 1090 503 1132 506
rect 1194 503 1197 523
rect 1682 513 1700 516
rect 1724 513 1733 516
rect 1738 513 1748 516
rect 1850 513 1853 525
rect 1874 523 1900 526
rect 1994 523 2028 526
rect 2034 523 2077 526
rect 2172 523 2189 526
rect 2282 523 2308 526
rect 2378 523 2388 526
rect 1868 513 1893 516
rect 2220 513 2245 516
rect 2276 513 2285 516
rect 2404 513 2437 516
rect 2450 506 2453 525
rect 2564 523 2636 526
rect 2650 523 2653 534
rect 2572 513 2597 516
rect 2652 513 2661 516
rect 1690 503 1716 506
rect 1834 503 1860 506
rect 2226 503 2268 506
rect 2410 503 2453 506
rect 14 467 2730 473
rect 450 433 492 436
rect 1938 433 1949 436
rect 212 423 237 426
rect 476 423 485 426
rect 642 423 652 426
rect 764 423 781 426
rect 940 423 965 426
rect 1316 423 1333 426
rect 1492 423 1509 426
rect 1738 423 1748 426
rect 1772 423 1797 426
rect 1938 417 1941 433
rect 122 413 140 416
rect 276 413 317 416
rect 338 413 365 416
rect 372 413 381 416
rect 436 413 469 416
rect 548 413 557 416
rect 610 413 628 416
rect 682 413 716 416
rect 730 413 748 416
rect 762 413 796 416
rect 820 413 829 416
rect 834 413 860 416
rect 884 413 917 416
rect 988 413 997 416
rect 1028 413 1053 416
rect 1074 413 1092 416
rect 1156 413 1173 416
rect 1218 413 1244 416
rect 1268 413 1293 416
rect 1346 413 1356 416
rect 1388 413 1405 416
rect 1442 413 1469 416
rect 1490 413 1509 416
rect 1580 413 1589 416
rect 1732 413 1741 416
rect 1778 413 1812 416
rect 1868 413 1893 416
rect 1924 414 1941 417
rect 1978 416 1981 436
rect 2058 433 2100 436
rect 2010 423 2028 426
rect 2066 423 2084 426
rect 2108 423 2117 426
rect 2266 416 2269 436
rect 2554 433 2573 436
rect 2538 423 2564 426
rect 1978 413 1997 416
rect 2146 413 2164 416
rect 2260 413 2269 416
rect 2300 413 2317 416
rect 2388 413 2397 416
rect 2442 413 2452 416
rect 2482 413 2524 416
rect 2570 415 2573 433
rect 2588 423 2621 426
rect 2652 423 2661 426
rect 2626 413 2636 416
rect 116 403 132 406
rect 226 403 252 406
rect 274 403 316 406
rect 338 405 341 413
rect 354 403 364 406
rect 378 403 381 413
rect 682 403 708 406
rect 764 403 773 406
rect 778 403 804 406
rect 914 405 917 413
rect 940 403 957 406
rect 980 403 1013 406
rect 1026 403 1052 406
rect 1066 403 1084 406
rect 1138 403 1148 406
rect 1170 405 1173 413
rect 1204 403 1213 406
rect 1242 403 1252 406
rect 1290 405 1293 413
rect 1362 403 1380 406
rect 1402 403 1412 406
rect 1466 405 1469 413
rect 1506 406 1509 413
rect 1492 403 1501 406
rect 1506 403 1516 406
rect 1602 403 1612 406
rect 1650 403 1660 406
rect 1698 403 1708 406
rect 1786 403 1804 406
rect 1842 403 1860 406
rect 1938 403 1964 406
rect 1994 405 1997 413
rect 2122 403 2132 406
rect 2242 403 2252 406
rect 2282 403 2292 406
rect 2314 405 2317 413
rect 2370 403 2380 406
rect 954 396 957 403
rect 954 393 972 396
rect 986 393 1012 396
rect 2394 395 2397 413
rect 2404 403 2460 406
rect 2506 403 2516 406
rect 2594 403 2628 406
rect 2652 403 2661 406
rect 2476 393 2501 396
rect 2194 383 2221 386
rect 38 367 2706 373
rect 394 343 412 346
rect 890 343 916 346
rect 1026 336 1029 345
rect 1042 343 1061 346
rect 1162 343 1196 346
rect 1690 343 1708 346
rect 2178 343 2204 346
rect 1058 336 1061 343
rect 180 323 205 326
rect 228 323 261 326
rect 298 325 301 336
rect 378 333 420 336
rect 426 333 436 336
rect 450 333 492 336
rect 530 333 548 336
rect 636 333 676 336
rect 682 333 701 336
rect 1018 333 1029 336
rect 1036 333 1053 336
rect 1058 333 1092 336
rect 1106 333 1124 336
rect 314 323 348 326
rect 428 323 477 326
rect 506 323 524 326
rect 538 323 556 326
rect 682 325 685 333
rect 1138 326 1141 334
rect 1204 333 1229 336
rect 1506 333 1540 336
rect 1564 333 1573 336
rect 1674 326 1677 334
rect 1716 333 1748 336
rect 1780 333 1797 336
rect 1834 326 1837 334
rect 1860 333 1869 336
rect 1874 333 1884 336
rect 1954 333 1964 336
rect 2042 327 2045 334
rect 2076 333 2101 336
rect 2130 333 2140 336
rect 2178 333 2212 336
rect 2218 333 2244 336
rect 2268 333 2277 336
rect 2282 333 2292 336
rect 2378 333 2404 336
rect 2474 333 2492 336
rect 2564 333 2612 336
rect 2618 333 2636 336
rect 690 323 724 326
rect 756 323 773 326
rect 804 323 813 326
rect 820 323 853 326
rect 1044 323 1061 326
rect 1100 323 1125 326
rect 1132 323 1141 326
rect 1148 323 1197 326
rect 1266 323 1277 326
rect 1338 323 1348 326
rect 1428 323 1445 326
rect 1492 323 1501 326
rect 1666 323 1677 326
rect 1684 323 1693 326
rect 1724 323 1741 326
rect 1820 323 1837 326
rect 1948 323 1957 326
rect 2036 324 2045 327
rect 2116 323 2141 326
rect 2234 323 2252 326
rect 2266 323 2300 326
rect 538 313 541 323
rect 1274 316 1277 323
rect 1666 316 1669 323
rect 564 313 597 316
rect 834 313 860 316
rect 1156 313 1165 316
rect 1218 313 1236 316
rect 1260 313 1269 316
rect 1274 313 1292 316
rect 1316 313 1333 316
rect 1618 313 1636 316
rect 1660 313 1669 316
rect 1860 313 1877 316
rect 1908 313 1917 316
rect 2268 313 2285 316
rect 2308 313 2341 316
rect 2338 306 2341 313
rect 2354 306 2357 325
rect 2412 323 2429 326
rect 2500 323 2509 326
rect 2514 323 2540 326
rect 2620 323 2629 326
rect 834 303 876 306
rect 938 303 956 306
rect 1274 303 1308 306
rect 1610 303 1652 306
rect 2338 303 2357 306
rect 14 267 2730 273
rect 578 233 597 236
rect 714 233 748 236
rect 578 226 581 233
rect 556 223 581 226
rect 660 223 685 226
rect 196 213 221 216
rect 330 213 380 216
rect 466 206 469 214
rect 500 213 533 216
rect 714 206 717 233
rect 876 223 885 226
rect 1036 223 1053 226
rect 1324 223 1333 226
rect 794 213 804 216
rect 850 213 860 216
rect 978 213 996 216
rect 1010 213 1020 216
rect 978 206 981 213
rect 1106 206 1109 214
rect 1114 213 1156 216
rect 1202 213 1220 216
rect 1226 213 1252 216
rect 1202 206 1205 213
rect 1330 206 1333 223
rect 1372 213 1389 216
rect 1436 213 1469 216
rect 1546 213 1580 216
rect 1594 213 1612 216
rect 1658 213 1668 216
rect 1706 213 1740 216
rect 1756 213 1797 216
rect 1884 213 1901 216
rect 1906 213 1916 216
rect 1940 213 1973 216
rect 2004 213 2013 216
rect 404 203 437 206
rect 442 203 452 206
rect 466 203 492 206
rect 522 203 532 206
rect 618 203 644 206
rect 700 203 717 206
rect 834 203 852 206
rect 890 203 924 206
rect 956 203 981 206
rect 1002 203 1012 206
rect 1036 203 1045 206
rect 1106 203 1148 206
rect 1180 203 1205 206
rect 1234 203 1244 206
rect 1274 203 1300 206
rect 1330 203 1364 206
rect 1404 203 1421 206
rect 1442 203 1468 206
rect 1532 203 1565 206
rect 1684 203 1725 206
rect 1762 203 1796 206
rect 1876 203 1924 206
rect 1946 203 1988 206
rect 2018 196 2021 216
rect 2084 213 2109 216
rect 2196 213 2213 216
rect 2250 213 2292 216
rect 2308 213 2357 216
rect 2500 213 2509 216
rect 2548 213 2589 216
rect 2642 213 2660 216
rect 2642 206 2645 213
rect 2124 203 2181 206
rect 2188 203 2221 206
rect 2252 203 2277 206
rect 2314 203 2356 206
rect 2428 203 2445 206
rect 2450 203 2484 206
rect 2498 203 2540 206
rect 2554 203 2588 206
rect 2620 203 2645 206
rect 316 193 365 196
rect 468 193 477 196
rect 666 193 692 196
rect 1506 193 1524 196
rect 2004 193 2037 196
rect 2394 193 2420 196
rect 38 167 2706 173
rect 538 143 548 146
rect 570 143 580 146
rect 666 143 684 146
rect 834 143 844 146
rect 922 143 940 146
rect 970 143 980 146
rect 1346 143 1372 146
rect 1778 143 1796 146
rect 2218 143 2236 146
rect 2250 143 2268 146
rect 2218 136 2221 143
rect 354 133 364 136
rect 378 133 404 136
rect 514 133 556 136
rect 562 133 588 136
rect 594 133 636 136
rect 666 133 692 136
rect 852 133 884 136
rect 916 133 948 136
rect 988 133 1021 136
rect 1194 133 1228 136
rect 1268 133 1308 136
rect 1340 133 1380 136
rect 1410 133 1420 136
rect 1458 133 1492 136
rect 1516 133 1549 136
rect 1562 133 1580 136
rect 1722 133 1756 136
rect 1770 133 1804 136
rect 276 123 301 126
rect 332 123 349 126
rect 434 123 452 126
rect 564 123 581 126
rect 596 123 637 126
rect 666 116 669 133
rect 764 123 789 126
rect 866 123 892 126
rect 1018 125 1021 133
rect 1546 126 1549 133
rect 1092 123 1117 126
rect 1162 123 1172 126
rect 1236 123 1245 126
rect 1282 123 1316 126
rect 1394 123 1428 126
rect 1500 123 1509 126
rect 1546 123 1572 126
rect 1596 123 1621 126
rect 1772 123 1797 126
rect 1810 125 1813 136
rect 2146 133 2164 136
rect 2188 133 2221 136
rect 2244 133 2261 136
rect 2276 133 2285 136
rect 2290 133 2332 136
rect 2410 133 2420 136
rect 2626 133 2644 136
rect 1924 123 1949 126
rect 2138 123 2172 126
rect 2298 123 2340 126
rect 2370 123 2412 126
rect 2436 123 2461 126
rect 660 113 669 116
rect 2090 113 2108 116
rect 2132 113 2157 116
rect 2098 103 2124 106
rect 14 67 2730 73
rect 38 37 2706 57
rect 14 13 2730 33
<< metal2 >>
rect 14 13 34 2527
rect 38 37 58 2503
rect 810 2453 853 2456
rect 82 2413 85 2436
rect 90 2413 109 2416
rect 90 2406 93 2413
rect 74 2403 93 2406
rect 90 2393 109 2396
rect 114 2316 117 2406
rect 146 2333 149 2406
rect 162 2403 165 2436
rect 170 2393 173 2416
rect 210 2413 213 2446
rect 234 2443 285 2446
rect 234 2423 237 2443
rect 242 2413 245 2436
rect 250 2433 269 2436
rect 194 2336 197 2406
rect 250 2366 253 2433
rect 170 2333 197 2336
rect 242 2363 253 2366
rect 122 2323 141 2326
rect 106 2313 117 2316
rect 122 2313 133 2316
rect 74 2213 77 2226
rect 90 2213 93 2256
rect 106 2213 109 2313
rect 114 2213 117 2226
rect 122 2206 125 2313
rect 138 2306 141 2323
rect 186 2313 189 2326
rect 138 2303 149 2306
rect 146 2236 149 2303
rect 138 2233 149 2236
rect 138 2213 141 2233
rect 178 2213 181 2226
rect 82 2193 85 2206
rect 106 2196 109 2206
rect 114 2203 125 2206
rect 130 2196 133 2206
rect 106 2193 133 2196
rect 82 2126 85 2136
rect 106 2133 109 2193
rect 74 2106 77 2126
rect 70 2103 77 2106
rect 82 2123 109 2126
rect 70 2026 73 2103
rect 70 2023 77 2026
rect 74 1983 77 2023
rect 82 2013 85 2123
rect 106 2113 117 2116
rect 106 1966 109 2026
rect 138 2006 141 2136
rect 170 2133 173 2206
rect 186 2203 189 2216
rect 194 2203 197 2326
rect 242 2323 245 2363
rect 258 2356 261 2426
rect 266 2423 269 2433
rect 250 2353 261 2356
rect 202 2193 205 2216
rect 218 2213 221 2236
rect 210 2156 213 2206
rect 226 2203 229 2246
rect 234 2233 237 2256
rect 242 2213 245 2226
rect 250 2213 253 2353
rect 266 2243 269 2416
rect 282 2413 285 2443
rect 290 2406 293 2446
rect 298 2413 301 2426
rect 306 2413 309 2436
rect 394 2433 421 2436
rect 394 2413 397 2433
rect 290 2403 309 2406
rect 418 2363 421 2433
rect 442 2346 445 2416
rect 522 2413 525 2436
rect 434 2343 445 2346
rect 298 2316 301 2336
rect 274 2313 301 2316
rect 322 2306 325 2326
rect 322 2303 333 2306
rect 282 2233 293 2236
rect 322 2233 325 2303
rect 338 2296 341 2336
rect 354 2333 389 2336
rect 346 2316 349 2326
rect 354 2323 357 2333
rect 362 2323 373 2326
rect 362 2316 365 2323
rect 346 2313 365 2316
rect 370 2303 373 2316
rect 338 2293 349 2296
rect 266 2206 269 2226
rect 290 2223 293 2233
rect 266 2203 277 2206
rect 194 2153 213 2156
rect 194 2133 197 2153
rect 202 2143 213 2146
rect 218 2136 221 2156
rect 162 2096 165 2126
rect 178 2103 181 2126
rect 194 2096 197 2126
rect 202 2116 205 2136
rect 210 2133 221 2136
rect 226 2123 229 2196
rect 282 2176 285 2216
rect 314 2213 317 2226
rect 330 2213 333 2226
rect 338 2213 341 2226
rect 346 2216 349 2293
rect 370 2223 373 2256
rect 346 2213 373 2216
rect 378 2213 381 2236
rect 386 2216 389 2333
rect 394 2316 397 2336
rect 434 2333 437 2343
rect 410 2323 437 2326
rect 394 2313 429 2316
rect 394 2226 397 2256
rect 394 2223 413 2226
rect 386 2213 397 2216
rect 370 2206 373 2213
rect 354 2196 357 2206
rect 370 2203 381 2206
rect 394 2196 397 2213
rect 354 2193 397 2196
rect 242 2173 285 2176
rect 202 2113 213 2116
rect 162 2093 197 2096
rect 162 2043 205 2046
rect 154 2023 157 2036
rect 162 2013 165 2043
rect 178 2013 189 2016
rect 194 2013 197 2036
rect 202 2013 205 2043
rect 138 2003 149 2006
rect 82 1963 109 1966
rect 74 1883 77 1926
rect 82 1923 85 1963
rect 146 1933 149 1946
rect 66 1873 93 1876
rect 66 1856 69 1873
rect 66 1853 77 1856
rect 74 1786 77 1853
rect 66 1783 77 1786
rect 66 1576 69 1783
rect 98 1766 101 1916
rect 146 1913 149 1926
rect 162 1896 165 2006
rect 186 1986 189 2006
rect 202 1993 205 2006
rect 210 1986 213 2113
rect 234 2093 237 2126
rect 242 2116 245 2173
rect 258 2133 269 2136
rect 274 2116 277 2136
rect 282 2123 285 2166
rect 290 2133 293 2146
rect 298 2116 301 2126
rect 242 2113 249 2116
rect 246 2056 249 2113
rect 266 2103 269 2116
rect 274 2113 301 2116
rect 298 2086 301 2113
rect 306 2093 309 2136
rect 362 2133 373 2136
rect 386 2133 389 2156
rect 338 2123 365 2126
rect 314 2086 317 2106
rect 330 2103 333 2116
rect 346 2113 357 2116
rect 346 2093 349 2106
rect 298 2083 317 2086
rect 246 2053 253 2056
rect 226 2013 229 2046
rect 250 2036 253 2053
rect 250 2033 285 2036
rect 186 1983 213 1986
rect 218 1983 221 2006
rect 186 1976 189 1983
rect 178 1973 189 1976
rect 178 1933 181 1973
rect 186 1933 189 1956
rect 170 1903 173 1926
rect 178 1923 189 1926
rect 202 1913 205 1926
rect 162 1893 189 1896
rect 82 1763 101 1766
rect 74 1733 77 1756
rect 82 1723 85 1763
rect 98 1636 101 1716
rect 74 1633 101 1636
rect 74 1603 77 1633
rect 122 1586 125 1796
rect 162 1743 165 1756
rect 138 1703 141 1716
rect 170 1646 173 1736
rect 178 1723 181 1746
rect 186 1736 189 1893
rect 186 1733 197 1736
rect 186 1713 189 1726
rect 170 1643 181 1646
rect 130 1613 133 1626
rect 130 1593 133 1606
rect 178 1603 181 1643
rect 194 1603 197 1733
rect 202 1693 205 1726
rect 202 1613 205 1636
rect 210 1603 213 1983
rect 218 1933 221 1946
rect 226 1933 229 1956
rect 218 1896 221 1916
rect 234 1913 245 1916
rect 218 1893 229 1896
rect 226 1776 229 1893
rect 250 1836 253 2033
rect 266 2006 269 2016
rect 258 2003 269 2006
rect 282 2006 285 2033
rect 290 2013 293 2046
rect 298 2023 301 2083
rect 346 2013 349 2026
rect 362 2013 365 2123
rect 370 2116 373 2133
rect 370 2113 381 2116
rect 378 2056 381 2113
rect 370 2053 381 2056
rect 282 2003 293 2006
rect 258 1993 261 2003
rect 266 1953 269 1996
rect 274 1983 277 1996
rect 346 1966 349 2006
rect 354 1983 357 2006
rect 346 1963 365 1966
rect 282 1943 301 1946
rect 282 1933 285 1943
rect 266 1923 285 1926
rect 282 1903 285 1916
rect 242 1833 253 1836
rect 242 1786 245 1833
rect 290 1823 293 1936
rect 298 1926 301 1943
rect 298 1923 305 1926
rect 302 1836 305 1923
rect 338 1876 341 1936
rect 362 1923 365 1963
rect 370 1903 373 2053
rect 410 2036 413 2223
rect 418 2123 421 2206
rect 434 2193 437 2323
rect 442 2306 445 2336
rect 458 2323 461 2336
rect 498 2333 501 2346
rect 522 2333 525 2386
rect 442 2303 453 2306
rect 450 2236 453 2303
rect 442 2233 453 2236
rect 442 2213 445 2233
rect 482 2226 485 2326
rect 506 2243 509 2326
rect 522 2226 525 2326
rect 538 2316 541 2406
rect 586 2376 589 2416
rect 634 2413 645 2416
rect 626 2376 629 2406
rect 586 2373 629 2376
rect 534 2313 541 2316
rect 534 2236 537 2313
rect 570 2306 573 2366
rect 594 2323 597 2346
rect 482 2223 525 2226
rect 530 2233 537 2236
rect 546 2303 573 2306
rect 482 2213 485 2223
rect 490 2213 501 2216
rect 442 2133 445 2206
rect 450 2126 453 2206
rect 482 2203 493 2206
rect 514 2193 517 2216
rect 530 2176 533 2233
rect 490 2173 533 2176
rect 466 2133 469 2166
rect 442 2123 453 2126
rect 418 2113 437 2116
rect 418 2103 421 2113
rect 426 2046 429 2106
rect 442 2093 445 2123
rect 474 2073 477 2116
rect 490 2096 493 2173
rect 546 2166 549 2303
rect 634 2276 637 2406
rect 626 2273 637 2276
rect 570 2213 573 2226
rect 626 2206 629 2273
rect 642 2223 645 2413
rect 650 2373 653 2436
rect 666 2393 669 2406
rect 666 2333 669 2366
rect 650 2296 653 2326
rect 698 2323 701 2386
rect 714 2376 717 2416
rect 746 2383 749 2416
rect 754 2376 757 2406
rect 762 2393 765 2406
rect 714 2373 757 2376
rect 762 2333 765 2376
rect 778 2326 781 2416
rect 810 2413 813 2453
rect 850 2413 853 2453
rect 978 2453 1021 2456
rect 930 2413 941 2416
rect 978 2413 981 2453
rect 1018 2413 1021 2453
rect 2050 2453 2093 2456
rect 786 2353 789 2406
rect 826 2393 829 2406
rect 794 2346 797 2376
rect 786 2343 821 2346
rect 650 2293 661 2296
rect 658 2236 661 2293
rect 746 2236 749 2326
rect 770 2303 773 2326
rect 778 2323 805 2326
rect 650 2233 661 2236
rect 730 2233 749 2236
rect 650 2213 653 2233
rect 658 2213 693 2216
rect 626 2203 637 2206
rect 634 2166 637 2203
rect 530 2163 589 2166
rect 486 2093 493 2096
rect 426 2043 437 2046
rect 394 2033 413 2036
rect 378 1896 381 1976
rect 394 1966 397 2033
rect 410 1973 413 2006
rect 434 1983 437 2043
rect 486 2026 489 2093
rect 482 2023 489 2026
rect 394 1963 413 1966
rect 298 1833 305 1836
rect 314 1873 341 1876
rect 370 1893 381 1896
rect 298 1813 301 1833
rect 242 1783 253 1786
rect 218 1773 229 1776
rect 218 1743 221 1773
rect 250 1756 253 1783
rect 266 1776 269 1806
rect 314 1776 317 1873
rect 266 1773 317 1776
rect 218 1703 221 1726
rect 218 1613 221 1626
rect 114 1583 125 1586
rect 66 1573 85 1576
rect 82 1466 85 1573
rect 114 1566 117 1583
rect 66 1463 85 1466
rect 106 1563 117 1566
rect 178 1563 197 1566
rect 106 1466 109 1563
rect 106 1463 113 1466
rect 66 363 69 1463
rect 82 1386 85 1406
rect 74 1383 85 1386
rect 74 1116 77 1383
rect 82 1316 85 1376
rect 110 1366 113 1463
rect 130 1426 133 1536
rect 178 1523 181 1563
rect 194 1536 197 1563
rect 218 1546 221 1606
rect 210 1543 221 1546
rect 194 1533 221 1536
rect 194 1476 197 1526
rect 226 1523 229 1756
rect 242 1753 253 1756
rect 306 1756 309 1773
rect 306 1753 317 1756
rect 242 1666 245 1753
rect 290 1733 293 1746
rect 274 1713 277 1726
rect 290 1666 293 1726
rect 314 1666 317 1753
rect 346 1736 349 1836
rect 370 1803 373 1893
rect 402 1876 405 1936
rect 398 1873 405 1876
rect 398 1756 401 1873
rect 410 1766 413 1963
rect 418 1933 429 1936
rect 418 1883 421 1933
rect 434 1873 437 1926
rect 450 1923 453 2016
rect 482 1973 485 2023
rect 418 1853 461 1856
rect 418 1813 421 1853
rect 450 1813 453 1826
rect 458 1813 461 1853
rect 466 1796 469 1946
rect 490 1923 493 2016
rect 450 1793 469 1796
rect 474 1793 477 1876
rect 410 1763 437 1766
rect 242 1663 293 1666
rect 306 1663 317 1666
rect 338 1733 349 1736
rect 234 1516 237 1606
rect 250 1603 253 1663
rect 274 1623 277 1636
rect 266 1533 269 1586
rect 122 1423 133 1426
rect 186 1473 197 1476
rect 206 1513 237 1516
rect 122 1386 125 1423
rect 130 1393 133 1416
rect 186 1406 189 1473
rect 206 1466 209 1513
rect 202 1463 209 1466
rect 202 1413 205 1463
rect 170 1393 173 1406
rect 186 1403 205 1406
rect 122 1383 133 1386
rect 130 1376 133 1383
rect 130 1373 141 1376
rect 110 1363 117 1366
rect 114 1346 117 1363
rect 90 1343 117 1346
rect 90 1333 93 1343
rect 82 1313 89 1316
rect 86 1196 89 1313
rect 98 1236 101 1336
rect 114 1276 117 1343
rect 138 1333 141 1373
rect 170 1336 173 1366
rect 170 1333 181 1336
rect 122 1286 125 1326
rect 162 1286 165 1326
rect 122 1283 165 1286
rect 178 1276 181 1333
rect 114 1273 133 1276
rect 98 1233 125 1236
rect 114 1213 117 1226
rect 122 1216 125 1233
rect 130 1226 133 1273
rect 162 1273 181 1276
rect 162 1236 165 1273
rect 162 1233 181 1236
rect 130 1223 149 1226
rect 122 1213 133 1216
rect 106 1203 117 1206
rect 130 1203 133 1213
rect 86 1193 109 1196
rect 82 1133 85 1156
rect 106 1126 109 1193
rect 114 1133 117 1203
rect 106 1123 117 1126
rect 74 1113 85 1116
rect 82 1036 85 1113
rect 74 1033 85 1036
rect 74 376 77 1033
rect 106 1016 109 1123
rect 114 1103 117 1116
rect 130 1113 133 1136
rect 138 1103 141 1126
rect 98 1013 109 1016
rect 98 956 101 1013
rect 98 953 109 956
rect 106 936 109 953
rect 82 813 85 936
rect 94 933 109 936
rect 122 933 125 1016
rect 94 846 97 933
rect 106 913 109 926
rect 90 843 97 846
rect 82 793 85 806
rect 90 613 93 843
rect 98 823 109 826
rect 98 743 101 823
rect 114 813 117 846
rect 138 803 141 816
rect 146 786 149 1223
rect 178 1166 181 1233
rect 202 1213 205 1403
rect 210 1386 213 1426
rect 218 1403 221 1506
rect 250 1453 253 1526
rect 290 1523 293 1606
rect 306 1583 309 1663
rect 330 1593 333 1616
rect 338 1536 341 1733
rect 346 1723 365 1726
rect 362 1693 365 1716
rect 370 1656 373 1736
rect 378 1733 381 1756
rect 398 1753 405 1756
rect 370 1653 377 1656
rect 362 1556 365 1576
rect 374 1566 377 1653
rect 386 1583 389 1616
rect 402 1613 405 1753
rect 426 1736 429 1756
rect 418 1733 429 1736
rect 418 1666 421 1733
rect 434 1676 437 1763
rect 434 1673 441 1676
rect 418 1663 429 1666
rect 426 1613 429 1663
rect 438 1606 441 1673
rect 402 1573 405 1606
rect 434 1603 441 1606
rect 418 1566 421 1596
rect 374 1563 397 1566
rect 362 1553 373 1556
rect 334 1533 341 1536
rect 370 1533 373 1553
rect 334 1486 337 1533
rect 346 1503 349 1526
rect 394 1523 397 1563
rect 414 1563 421 1566
rect 434 1566 437 1603
rect 450 1573 453 1793
rect 482 1723 485 1826
rect 490 1823 493 1836
rect 498 1806 501 2086
rect 522 2016 525 2116
rect 494 1803 501 1806
rect 506 2013 525 2016
rect 494 1716 497 1803
rect 506 1766 509 2013
rect 530 2006 533 2163
rect 586 2133 589 2163
rect 626 2163 637 2166
rect 538 2086 541 2126
rect 538 2083 557 2086
rect 514 1993 517 2006
rect 522 2003 533 2006
rect 522 1976 525 2003
rect 530 1983 533 1996
rect 514 1973 525 1976
rect 514 1943 517 1973
rect 538 1933 541 2066
rect 554 2013 557 2083
rect 562 2013 565 2076
rect 570 1966 573 2126
rect 610 2123 613 2136
rect 626 2086 629 2163
rect 626 2083 637 2086
rect 634 2063 637 2083
rect 658 2073 661 2213
rect 682 2203 717 2206
rect 674 2193 685 2196
rect 666 2056 669 2126
rect 650 2053 669 2056
rect 610 2006 613 2016
rect 578 2003 613 2006
rect 610 1966 613 2003
rect 570 1963 589 1966
rect 562 1933 565 1946
rect 530 1923 549 1926
rect 586 1923 589 1963
rect 602 1963 613 1966
rect 626 1966 629 2016
rect 634 1993 637 2026
rect 626 1963 633 1966
rect 514 1796 517 1906
rect 530 1846 533 1923
rect 602 1886 605 1963
rect 602 1883 613 1886
rect 522 1843 533 1846
rect 522 1803 525 1843
rect 530 1813 533 1836
rect 538 1833 541 1846
rect 538 1803 541 1826
rect 514 1793 525 1796
rect 506 1763 517 1766
rect 474 1713 497 1716
rect 474 1576 477 1713
rect 514 1623 517 1763
rect 490 1613 501 1616
rect 490 1596 493 1606
rect 458 1573 477 1576
rect 482 1593 493 1596
rect 434 1563 441 1566
rect 414 1506 417 1563
rect 410 1503 417 1506
rect 334 1483 341 1486
rect 226 1433 261 1436
rect 226 1413 229 1433
rect 258 1413 261 1433
rect 338 1426 341 1483
rect 306 1423 341 1426
rect 298 1393 301 1406
rect 306 1403 309 1423
rect 314 1413 325 1416
rect 322 1386 325 1406
rect 330 1393 333 1416
rect 338 1403 341 1423
rect 370 1413 373 1456
rect 410 1436 413 1503
rect 438 1486 441 1563
rect 434 1483 441 1486
rect 410 1433 417 1436
rect 386 1403 389 1416
rect 210 1383 217 1386
rect 322 1383 333 1386
rect 214 1316 217 1383
rect 226 1333 229 1346
rect 242 1316 245 1326
rect 250 1323 253 1336
rect 258 1316 261 1336
rect 214 1313 221 1316
rect 242 1313 261 1316
rect 266 1316 269 1326
rect 290 1323 293 1346
rect 298 1316 301 1326
rect 266 1313 301 1316
rect 218 1246 221 1313
rect 210 1243 221 1246
rect 202 1186 205 1206
rect 210 1196 213 1243
rect 226 1203 229 1226
rect 210 1193 237 1196
rect 202 1183 221 1186
rect 162 1163 181 1166
rect 162 1106 165 1163
rect 170 1143 197 1146
rect 202 1143 205 1176
rect 178 1133 205 1136
rect 210 1133 213 1156
rect 218 1133 221 1183
rect 202 1126 205 1133
rect 194 1113 197 1126
rect 202 1123 221 1126
rect 162 1103 173 1106
rect 170 976 173 1103
rect 218 1093 221 1123
rect 234 1086 237 1193
rect 250 1153 253 1206
rect 258 1106 261 1266
rect 306 1256 309 1336
rect 314 1333 325 1336
rect 330 1316 333 1383
rect 298 1253 309 1256
rect 266 1223 293 1226
rect 162 973 173 976
rect 194 1083 237 1086
rect 250 1103 261 1106
rect 162 936 165 973
rect 154 933 165 936
rect 154 896 157 933
rect 162 913 165 926
rect 154 893 165 896
rect 162 826 165 893
rect 142 783 149 786
rect 154 823 165 826
rect 98 713 101 736
rect 142 726 145 783
rect 106 723 117 726
rect 130 676 133 726
rect 142 723 149 726
rect 154 723 157 823
rect 178 813 189 816
rect 162 793 165 806
rect 170 783 173 796
rect 178 776 181 813
rect 186 793 189 806
rect 170 773 181 776
rect 162 743 165 756
rect 170 733 173 773
rect 178 763 181 773
rect 146 706 149 723
rect 186 713 189 726
rect 146 703 157 706
rect 130 673 141 676
rect 98 603 101 626
rect 114 623 133 626
rect 114 616 117 623
rect 106 613 117 616
rect 130 606 133 623
rect 138 613 141 673
rect 154 636 157 703
rect 154 633 173 636
rect 146 613 149 626
rect 122 603 133 606
rect 90 533 93 546
rect 90 403 93 526
rect 114 523 117 536
rect 98 413 101 426
rect 114 423 117 516
rect 122 513 125 603
rect 154 583 157 606
rect 162 603 165 626
rect 146 543 149 556
rect 154 533 157 546
rect 170 513 173 633
rect 178 543 181 626
rect 186 613 189 626
rect 186 583 189 606
rect 178 503 181 526
rect 186 486 189 526
rect 178 483 189 486
rect 178 426 181 483
rect 178 423 189 426
rect 74 373 101 376
rect 98 293 101 373
rect 122 323 125 416
rect 186 403 189 423
rect 194 353 197 1083
rect 250 1036 253 1103
rect 226 1016 229 1036
rect 250 1033 261 1036
rect 218 1013 229 1016
rect 258 1016 261 1033
rect 266 1023 269 1186
rect 274 1023 277 1216
rect 290 1213 293 1223
rect 282 1133 285 1146
rect 282 1103 285 1116
rect 290 1033 293 1206
rect 298 1123 301 1253
rect 314 1246 317 1316
rect 306 1243 317 1246
rect 326 1313 333 1316
rect 306 1123 309 1243
rect 326 1236 329 1313
rect 318 1233 329 1236
rect 318 1176 321 1233
rect 338 1203 341 1386
rect 394 1363 397 1416
rect 414 1356 417 1433
rect 434 1413 437 1483
rect 450 1413 453 1536
rect 458 1413 461 1573
rect 466 1413 469 1536
rect 482 1523 485 1593
rect 498 1586 501 1606
rect 490 1583 501 1586
rect 490 1543 493 1583
rect 498 1523 501 1536
rect 506 1533 509 1586
rect 506 1506 509 1526
rect 498 1503 509 1506
rect 474 1466 477 1486
rect 474 1463 485 1466
rect 482 1406 485 1463
rect 498 1436 501 1503
rect 498 1433 509 1436
rect 506 1413 509 1433
rect 426 1403 445 1406
rect 442 1393 445 1403
rect 450 1373 453 1406
rect 474 1403 485 1406
rect 346 1343 349 1356
rect 386 1353 417 1356
rect 314 1173 321 1176
rect 314 1046 317 1173
rect 322 1133 325 1156
rect 330 1143 333 1166
rect 322 1103 325 1116
rect 314 1043 321 1046
rect 258 1013 273 1016
rect 202 923 205 1006
rect 218 926 221 1013
rect 234 953 237 1006
rect 258 936 261 1006
rect 234 933 261 936
rect 270 936 273 1013
rect 290 1003 293 1016
rect 282 943 285 956
rect 270 933 277 936
rect 218 923 229 926
rect 226 856 229 923
rect 250 856 253 926
rect 226 853 237 856
rect 250 853 261 856
rect 226 803 229 846
rect 234 816 237 853
rect 242 823 245 836
rect 234 813 245 816
rect 226 743 229 766
rect 202 723 205 736
rect 210 733 237 736
rect 210 723 229 726
rect 202 523 205 616
rect 210 523 213 723
rect 234 706 237 733
rect 226 703 237 706
rect 226 606 229 703
rect 242 613 245 813
rect 258 733 261 853
rect 266 733 269 916
rect 250 696 253 716
rect 274 703 277 933
rect 282 823 285 916
rect 282 783 285 806
rect 290 766 293 996
rect 318 976 321 1043
rect 314 973 321 976
rect 314 956 317 973
rect 306 953 317 956
rect 306 906 309 953
rect 306 903 317 906
rect 314 883 317 903
rect 322 876 325 946
rect 330 943 333 1136
rect 338 1013 341 1176
rect 346 1133 349 1246
rect 354 1213 357 1236
rect 354 1146 357 1206
rect 362 1203 365 1336
rect 386 1313 389 1353
rect 394 1343 429 1346
rect 394 1333 397 1343
rect 394 1303 397 1326
rect 402 1286 405 1326
rect 410 1303 413 1336
rect 426 1326 429 1343
rect 434 1343 469 1346
rect 434 1333 437 1343
rect 442 1326 445 1336
rect 402 1283 413 1286
rect 402 1226 405 1283
rect 418 1253 421 1326
rect 426 1323 445 1326
rect 442 1246 445 1316
rect 370 1223 405 1226
rect 426 1243 445 1246
rect 354 1143 365 1146
rect 354 1056 357 1126
rect 370 1086 373 1223
rect 378 1193 381 1216
rect 378 1133 381 1186
rect 386 1173 389 1216
rect 410 1203 413 1216
rect 378 1116 381 1126
rect 386 1123 389 1146
rect 378 1113 397 1116
rect 378 1103 381 1113
rect 370 1083 381 1086
rect 354 1053 365 1056
rect 362 976 365 1053
rect 354 973 365 976
rect 354 886 357 973
rect 378 956 381 1083
rect 402 1043 405 1196
rect 418 1143 421 1216
rect 426 1206 429 1243
rect 434 1213 437 1236
rect 442 1213 445 1243
rect 450 1206 453 1326
rect 466 1323 469 1343
rect 426 1203 433 1206
rect 442 1203 453 1206
rect 418 1016 421 1136
rect 430 1086 433 1203
rect 458 1193 461 1306
rect 474 1263 477 1403
rect 482 1313 485 1336
rect 442 1096 445 1166
rect 450 1103 453 1126
rect 442 1093 449 1096
rect 430 1083 437 1086
rect 370 953 381 956
rect 370 936 373 953
rect 314 873 325 876
rect 346 883 357 886
rect 366 933 373 936
rect 282 763 293 766
rect 250 693 261 696
rect 258 646 261 693
rect 250 643 261 646
rect 250 613 253 643
rect 282 636 285 763
rect 290 733 293 756
rect 298 713 301 846
rect 306 813 309 836
rect 314 796 317 873
rect 346 823 349 883
rect 366 866 369 933
rect 366 863 373 866
rect 362 823 365 846
rect 310 793 317 796
rect 310 696 313 793
rect 306 693 313 696
rect 282 633 293 636
rect 266 616 269 626
rect 258 613 269 616
rect 226 603 237 606
rect 234 566 237 603
rect 218 563 237 566
rect 218 516 221 563
rect 210 513 221 516
rect 210 446 213 513
rect 202 443 213 446
rect 202 323 205 443
rect 210 403 213 426
rect 226 403 229 556
rect 258 546 261 613
rect 266 583 269 606
rect 274 573 277 606
rect 290 576 293 633
rect 282 573 293 576
rect 306 576 309 693
rect 306 573 317 576
rect 234 533 237 546
rect 242 543 269 546
rect 242 513 245 543
rect 258 446 261 526
rect 266 513 269 543
rect 258 443 269 446
rect 234 423 261 426
rect 242 413 253 416
rect 258 413 261 423
rect 218 333 253 336
rect 170 153 173 296
rect 218 213 221 236
rect 250 213 253 333
rect 258 323 261 406
rect 266 403 269 443
rect 274 403 277 506
rect 282 413 285 573
rect 298 543 301 556
rect 290 506 293 526
rect 290 503 297 506
rect 294 396 297 503
rect 266 333 269 396
rect 290 393 297 396
rect 290 373 293 393
rect 274 353 301 356
rect 274 323 277 353
rect 282 333 285 346
rect 290 306 293 336
rect 298 333 301 353
rect 282 303 293 306
rect 282 236 285 303
rect 282 233 293 236
rect 290 213 293 233
rect 306 206 309 536
rect 314 503 317 573
rect 322 556 325 816
rect 362 806 365 816
rect 346 803 365 806
rect 338 733 341 776
rect 362 623 365 636
rect 330 613 341 616
rect 346 596 349 616
rect 362 603 365 616
rect 338 593 349 596
rect 322 553 333 556
rect 322 523 325 546
rect 330 496 333 553
rect 338 533 341 593
rect 362 533 365 556
rect 346 523 357 526
rect 314 493 333 496
rect 314 413 317 493
rect 322 383 325 416
rect 338 413 341 426
rect 354 403 357 446
rect 362 413 365 516
rect 370 406 373 863
rect 378 856 381 936
rect 386 893 389 936
rect 394 903 397 936
rect 378 853 389 856
rect 378 763 381 816
rect 386 783 389 853
rect 402 766 405 1016
rect 418 1013 429 1016
rect 434 996 437 1083
rect 446 1036 449 1093
rect 446 1033 453 1036
rect 450 1013 453 1033
rect 410 936 413 946
rect 426 943 429 996
rect 434 993 445 996
rect 442 946 445 993
rect 434 943 445 946
rect 410 933 429 936
rect 410 906 413 926
rect 426 916 429 933
rect 434 923 437 943
rect 458 926 461 1156
rect 466 1123 469 1146
rect 474 1123 477 1136
rect 482 1133 485 1186
rect 490 1133 493 1326
rect 498 1323 509 1326
rect 514 1303 517 1556
rect 522 1393 525 1793
rect 530 1613 533 1796
rect 538 1703 541 1726
rect 530 1423 533 1606
rect 530 1403 533 1416
rect 538 1366 541 1526
rect 546 1506 549 1856
rect 554 1823 557 1836
rect 562 1823 565 1866
rect 570 1816 573 1846
rect 594 1843 605 1846
rect 554 1813 573 1816
rect 554 1723 557 1813
rect 554 1603 557 1626
rect 562 1623 565 1806
rect 578 1796 581 1836
rect 574 1793 581 1796
rect 586 1796 589 1826
rect 602 1813 605 1843
rect 586 1793 597 1796
rect 610 1793 613 1883
rect 630 1876 633 1963
rect 630 1873 637 1876
rect 574 1736 577 1793
rect 594 1746 597 1793
rect 618 1763 621 1826
rect 626 1756 629 1836
rect 586 1743 597 1746
rect 610 1753 629 1756
rect 574 1733 581 1736
rect 578 1716 581 1733
rect 586 1723 589 1743
rect 610 1723 613 1753
rect 578 1713 597 1716
rect 570 1703 589 1706
rect 586 1616 589 1703
rect 594 1623 597 1713
rect 610 1646 613 1716
rect 610 1643 621 1646
rect 602 1623 605 1636
rect 610 1616 613 1626
rect 578 1526 581 1616
rect 586 1613 613 1616
rect 618 1613 621 1643
rect 626 1596 629 1636
rect 622 1593 629 1596
rect 602 1533 605 1576
rect 610 1526 613 1546
rect 622 1536 625 1593
rect 554 1523 581 1526
rect 546 1503 557 1506
rect 554 1446 557 1503
rect 546 1443 557 1446
rect 546 1413 549 1443
rect 530 1363 541 1366
rect 522 1333 525 1346
rect 498 1196 501 1216
rect 506 1213 517 1216
rect 522 1213 525 1326
rect 498 1193 525 1196
rect 466 953 469 1026
rect 458 923 465 926
rect 426 913 453 916
rect 410 903 445 906
rect 434 816 437 886
rect 410 803 413 816
rect 418 813 437 816
rect 402 763 409 766
rect 386 723 389 736
rect 406 686 409 763
rect 386 616 389 686
rect 402 683 409 686
rect 402 633 405 683
rect 418 636 421 813
rect 426 803 437 806
rect 442 803 445 903
rect 450 786 453 913
rect 462 806 465 923
rect 474 873 477 1046
rect 482 1003 485 1126
rect 490 1093 493 1126
rect 498 1053 501 1136
rect 506 1026 509 1136
rect 514 1106 517 1176
rect 522 1123 525 1193
rect 530 1153 533 1363
rect 538 1333 541 1356
rect 554 1333 557 1406
rect 546 1313 549 1326
rect 514 1103 525 1106
rect 522 1036 525 1103
rect 490 1023 509 1026
rect 514 1033 525 1036
rect 482 883 485 926
rect 490 906 493 1023
rect 514 1016 517 1033
rect 506 1013 517 1016
rect 538 1013 541 1256
rect 562 1243 565 1406
rect 578 1393 581 1456
rect 578 1346 581 1376
rect 586 1353 589 1526
rect 594 1523 613 1526
rect 618 1533 625 1536
rect 618 1506 621 1533
rect 610 1503 621 1506
rect 610 1456 613 1503
rect 610 1453 621 1456
rect 570 1306 573 1346
rect 578 1343 589 1346
rect 586 1326 589 1343
rect 594 1333 597 1396
rect 602 1333 605 1406
rect 610 1386 613 1416
rect 618 1393 621 1453
rect 634 1413 637 1873
rect 642 1853 645 2026
rect 650 1903 653 2053
rect 658 2003 661 2046
rect 674 2013 677 2166
rect 682 2006 685 2193
rect 706 2133 709 2146
rect 690 2113 693 2126
rect 714 2103 717 2126
rect 722 2096 725 2216
rect 730 2163 733 2233
rect 706 2093 725 2096
rect 666 2003 685 2006
rect 658 1933 661 1976
rect 666 1936 669 1996
rect 674 1943 677 2003
rect 690 1993 693 2016
rect 698 1943 701 2076
rect 706 2013 709 2093
rect 730 2043 733 2126
rect 666 1933 677 1936
rect 658 1853 661 1926
rect 666 1893 669 1926
rect 642 1813 645 1836
rect 650 1746 653 1826
rect 658 1813 661 1846
rect 674 1836 677 1933
rect 682 1853 693 1856
rect 666 1833 677 1836
rect 650 1743 661 1746
rect 658 1723 661 1743
rect 642 1703 645 1716
rect 650 1646 653 1716
rect 658 1703 661 1716
rect 642 1643 653 1646
rect 642 1633 645 1643
rect 650 1623 653 1636
rect 658 1603 661 1626
rect 642 1533 645 1576
rect 666 1536 669 1833
rect 674 1706 677 1826
rect 682 1823 685 1836
rect 690 1803 693 1853
rect 698 1813 701 1846
rect 706 1776 709 1976
rect 714 1943 717 2006
rect 714 1813 717 1926
rect 722 1813 725 1936
rect 730 1916 733 2016
rect 738 1973 741 2226
rect 778 2213 781 2323
rect 810 2306 813 2336
rect 802 2303 813 2306
rect 802 2236 805 2303
rect 786 2233 805 2236
rect 746 2203 765 2206
rect 746 2003 749 2136
rect 754 2106 757 2136
rect 786 2133 789 2233
rect 818 2226 821 2343
rect 834 2293 837 2346
rect 850 2323 853 2336
rect 866 2333 869 2356
rect 898 2323 901 2336
rect 906 2323 909 2346
rect 914 2333 925 2336
rect 930 2326 933 2413
rect 946 2386 949 2406
rect 994 2393 997 2406
rect 946 2383 989 2386
rect 914 2323 933 2326
rect 890 2313 901 2316
rect 802 2213 805 2226
rect 810 2223 821 2226
rect 810 2213 837 2216
rect 810 2206 813 2213
rect 794 2203 813 2206
rect 762 2123 781 2126
rect 754 2103 765 2106
rect 778 2103 781 2116
rect 762 2036 765 2103
rect 754 2033 765 2036
rect 754 2013 757 2033
rect 770 2013 789 2016
rect 738 1933 741 1966
rect 730 1913 737 1916
rect 734 1846 737 1913
rect 746 1906 749 1996
rect 754 1923 757 2006
rect 794 1996 797 2136
rect 826 2133 829 2146
rect 834 2133 853 2136
rect 834 2126 837 2133
rect 810 2123 837 2126
rect 826 2093 829 2116
rect 826 2013 829 2036
rect 842 2013 845 2126
rect 850 2123 853 2133
rect 858 2123 861 2136
rect 866 2106 869 2206
rect 874 2156 877 2226
rect 906 2223 909 2256
rect 882 2176 885 2206
rect 890 2193 893 2216
rect 914 2196 917 2323
rect 922 2296 925 2316
rect 922 2293 933 2296
rect 930 2246 933 2293
rect 946 2246 949 2326
rect 922 2243 933 2246
rect 942 2243 949 2246
rect 962 2243 965 2336
rect 970 2323 973 2336
rect 986 2333 989 2383
rect 1090 2376 1093 2416
rect 1154 2413 1157 2426
rect 1210 2406 1213 2416
rect 1218 2413 1221 2426
rect 1106 2393 1109 2406
rect 1090 2373 1137 2376
rect 1002 2323 1005 2346
rect 1090 2343 1125 2346
rect 978 2313 989 2316
rect 922 2203 925 2243
rect 930 2213 933 2226
rect 914 2193 925 2196
rect 882 2173 893 2176
rect 874 2153 881 2156
rect 858 2103 869 2106
rect 858 2036 861 2103
rect 878 2096 881 2153
rect 874 2093 881 2096
rect 858 2033 869 2036
rect 770 1993 797 1996
rect 818 1993 821 2006
rect 770 1936 773 1993
rect 770 1933 781 1936
rect 834 1933 837 2006
rect 858 1933 861 1956
rect 746 1903 757 1906
rect 730 1843 737 1846
rect 690 1773 709 1776
rect 674 1703 685 1706
rect 674 1543 677 1606
rect 682 1536 685 1616
rect 650 1533 669 1536
rect 674 1533 685 1536
rect 690 1536 693 1773
rect 698 1713 701 1726
rect 698 1583 701 1626
rect 706 1543 709 1766
rect 730 1743 733 1843
rect 754 1836 757 1903
rect 778 1876 781 1933
rect 746 1833 757 1836
rect 770 1873 781 1876
rect 738 1803 741 1826
rect 714 1703 717 1726
rect 730 1713 733 1736
rect 722 1696 725 1706
rect 738 1703 741 1736
rect 746 1696 749 1833
rect 770 1826 773 1873
rect 770 1823 781 1826
rect 722 1693 749 1696
rect 722 1673 725 1693
rect 754 1686 757 1816
rect 762 1703 765 1806
rect 778 1803 781 1823
rect 738 1683 757 1686
rect 690 1533 701 1536
rect 650 1516 653 1533
rect 646 1513 653 1516
rect 646 1466 649 1513
rect 658 1473 661 1526
rect 666 1523 693 1526
rect 698 1506 701 1533
rect 690 1503 701 1506
rect 646 1463 653 1466
rect 634 1386 637 1406
rect 650 1393 653 1463
rect 690 1436 693 1503
rect 690 1433 701 1436
rect 674 1413 685 1416
rect 610 1383 637 1386
rect 586 1323 605 1326
rect 602 1306 605 1323
rect 570 1303 581 1306
rect 578 1256 581 1303
rect 570 1253 581 1256
rect 594 1303 605 1306
rect 570 1236 573 1253
rect 594 1246 597 1303
rect 594 1243 605 1246
rect 562 1233 573 1236
rect 546 1153 549 1206
rect 554 1183 557 1206
rect 562 1173 565 1233
rect 570 1223 589 1226
rect 570 1213 581 1216
rect 586 1206 589 1223
rect 546 1136 549 1146
rect 546 1133 565 1136
rect 546 1013 557 1016
rect 506 946 509 1013
rect 514 1003 525 1006
rect 530 996 533 1006
rect 546 1003 549 1013
rect 530 993 541 996
rect 554 993 557 1006
rect 506 943 533 946
rect 498 923 501 936
rect 506 933 517 936
rect 498 913 509 916
rect 490 903 509 906
rect 462 803 477 806
rect 482 803 485 816
rect 458 793 469 796
rect 414 633 421 636
rect 434 783 469 786
rect 378 613 389 616
rect 378 503 381 613
rect 386 503 389 606
rect 362 403 373 406
rect 314 303 317 366
rect 314 213 317 236
rect 298 203 309 206
rect 330 193 333 356
rect 338 343 349 346
rect 338 333 341 343
rect 346 333 357 336
rect 362 313 365 403
rect 378 396 381 406
rect 370 393 381 396
rect 394 396 397 576
rect 414 556 417 633
rect 426 573 429 626
rect 414 553 421 556
rect 418 536 421 553
rect 434 543 437 783
rect 466 743 469 783
rect 474 726 477 803
rect 442 713 445 726
rect 466 723 477 726
rect 482 723 485 786
rect 490 723 493 806
rect 498 733 501 806
rect 466 656 469 723
rect 506 716 509 903
rect 514 793 517 806
rect 522 746 525 876
rect 530 776 533 943
rect 538 813 541 993
rect 562 933 565 1116
rect 570 1106 573 1206
rect 578 1203 589 1206
rect 594 1203 597 1216
rect 578 1186 581 1203
rect 602 1193 605 1243
rect 610 1216 613 1383
rect 642 1333 645 1386
rect 626 1306 629 1326
rect 622 1303 629 1306
rect 622 1236 625 1303
rect 642 1286 645 1326
rect 650 1323 653 1346
rect 666 1326 669 1336
rect 658 1323 669 1326
rect 658 1313 661 1323
rect 666 1296 669 1316
rect 662 1293 669 1296
rect 642 1283 653 1286
rect 622 1233 629 1236
rect 610 1213 621 1216
rect 578 1183 589 1186
rect 578 1116 581 1136
rect 586 1123 589 1183
rect 578 1113 589 1116
rect 570 1103 581 1106
rect 546 873 549 926
rect 554 876 557 926
rect 570 923 573 936
rect 578 886 581 1103
rect 586 1093 589 1113
rect 594 1003 597 1186
rect 586 893 589 916
rect 594 906 597 956
rect 602 913 605 1136
rect 610 953 613 1206
rect 618 1156 621 1206
rect 626 1163 629 1233
rect 634 1196 637 1276
rect 650 1226 653 1283
rect 642 1223 653 1226
rect 662 1226 665 1293
rect 662 1223 669 1226
rect 674 1223 677 1413
rect 682 1333 685 1406
rect 698 1366 701 1433
rect 706 1413 709 1496
rect 714 1453 717 1636
rect 722 1613 725 1626
rect 722 1523 725 1576
rect 738 1556 741 1683
rect 746 1633 749 1676
rect 738 1553 749 1556
rect 730 1513 733 1526
rect 738 1496 741 1546
rect 730 1493 741 1496
rect 730 1426 733 1493
rect 730 1423 741 1426
rect 722 1383 725 1406
rect 738 1393 741 1423
rect 698 1363 733 1366
rect 690 1323 693 1336
rect 714 1333 717 1346
rect 698 1323 717 1326
rect 642 1203 645 1223
rect 650 1203 661 1206
rect 634 1193 653 1196
rect 658 1193 661 1203
rect 642 1166 645 1186
rect 638 1163 645 1166
rect 618 1153 629 1156
rect 594 903 601 906
rect 578 883 589 886
rect 554 873 565 876
rect 562 823 565 873
rect 538 783 541 806
rect 546 786 549 816
rect 554 803 565 806
rect 546 783 553 786
rect 586 783 589 883
rect 598 846 601 903
rect 598 843 605 846
rect 594 813 597 826
rect 530 773 537 776
rect 490 713 509 716
rect 514 743 525 746
rect 466 653 477 656
rect 458 623 461 636
rect 450 546 453 616
rect 466 613 469 626
rect 442 543 453 546
rect 402 493 405 526
rect 402 413 405 426
rect 410 403 413 536
rect 418 533 437 536
rect 418 443 421 516
rect 394 393 413 396
rect 418 393 421 416
rect 426 403 429 506
rect 434 476 437 533
rect 442 493 445 543
rect 434 473 441 476
rect 370 333 373 393
rect 410 386 413 393
rect 378 333 381 346
rect 394 343 397 386
rect 410 383 429 386
rect 426 293 429 383
rect 438 296 441 473
rect 450 433 453 536
rect 458 483 461 526
rect 466 476 469 576
rect 474 533 477 653
rect 482 603 485 616
rect 490 603 493 713
rect 514 573 517 743
rect 522 723 525 736
rect 534 716 537 773
rect 550 726 553 783
rect 562 743 565 766
rect 550 723 557 726
rect 534 713 541 716
rect 530 613 533 646
rect 538 606 541 713
rect 554 636 557 723
rect 522 526 525 606
rect 490 523 525 526
rect 530 603 541 606
rect 546 633 557 636
rect 490 493 493 523
rect 530 496 533 603
rect 538 533 541 546
rect 458 473 469 476
rect 458 346 461 473
rect 514 456 517 476
rect 510 453 517 456
rect 466 443 501 446
rect 466 413 469 443
rect 482 423 485 436
rect 498 423 501 443
rect 482 363 485 416
rect 510 366 513 453
rect 522 403 525 496
rect 530 493 541 496
rect 530 413 533 426
rect 510 363 517 366
rect 458 343 465 346
rect 482 343 509 346
rect 434 293 441 296
rect 250 133 253 156
rect 298 113 301 126
rect 346 123 349 146
rect 354 133 357 206
rect 370 203 373 226
rect 394 213 405 216
rect 434 213 437 293
rect 442 213 445 256
rect 362 146 365 196
rect 378 146 381 156
rect 362 143 381 146
rect 370 133 381 136
rect 370 126 373 133
rect 386 126 389 206
rect 394 143 397 176
rect 354 123 373 126
rect 378 113 381 126
rect 386 123 413 126
rect 434 123 437 206
rect 442 143 445 206
rect 450 203 453 336
rect 462 246 465 343
rect 458 243 465 246
rect 458 153 461 243
rect 466 213 469 226
rect 474 193 477 326
rect 498 323 501 336
rect 506 323 509 343
rect 514 333 517 363
rect 498 176 501 306
rect 522 203 525 376
rect 538 373 541 493
rect 546 446 549 633
rect 554 533 557 616
rect 562 596 565 606
rect 570 603 573 736
rect 602 726 605 843
rect 610 736 613 946
rect 618 746 621 1136
rect 626 1073 629 1153
rect 626 1033 629 1056
rect 638 1046 641 1163
rect 638 1043 645 1046
rect 626 1003 629 1016
rect 634 943 637 1026
rect 642 1013 645 1043
rect 626 903 629 916
rect 634 883 637 926
rect 626 813 629 826
rect 634 813 637 836
rect 650 813 653 1193
rect 658 1133 661 1146
rect 666 1126 669 1223
rect 658 1123 669 1126
rect 658 1103 661 1123
rect 658 993 661 1026
rect 666 933 669 946
rect 674 916 677 1216
rect 682 1196 685 1216
rect 690 1203 693 1316
rect 698 1213 701 1236
rect 682 1193 693 1196
rect 682 1083 685 1136
rect 690 1066 693 1193
rect 714 1183 717 1206
rect 722 1146 725 1356
rect 730 1306 733 1363
rect 746 1333 749 1553
rect 754 1543 757 1666
rect 762 1533 765 1696
rect 770 1623 773 1796
rect 770 1523 773 1586
rect 778 1553 781 1746
rect 786 1706 789 1866
rect 802 1826 805 1926
rect 810 1906 813 1926
rect 834 1913 837 1926
rect 866 1916 869 2033
rect 874 1936 877 2093
rect 890 2076 893 2173
rect 882 2073 893 2076
rect 882 2043 885 2073
rect 906 2063 909 2116
rect 914 2066 917 2136
rect 922 2123 925 2193
rect 930 2093 933 2206
rect 942 2156 945 2243
rect 954 2213 965 2216
rect 942 2153 949 2156
rect 938 2123 941 2136
rect 946 2133 949 2153
rect 954 2076 957 2213
rect 962 2193 965 2206
rect 986 2156 989 2313
rect 1018 2263 1021 2336
rect 1034 2333 1045 2336
rect 1058 2296 1061 2316
rect 1050 2293 1061 2296
rect 994 2203 997 2226
rect 982 2153 989 2156
rect 970 2113 973 2126
rect 982 2086 985 2153
rect 994 2133 997 2146
rect 1002 2133 1005 2206
rect 1026 2186 1029 2226
rect 1034 2203 1037 2246
rect 1050 2236 1053 2293
rect 1050 2233 1061 2236
rect 1058 2213 1061 2233
rect 1018 2183 1029 2186
rect 994 2093 997 2126
rect 982 2083 989 2086
rect 954 2073 965 2076
rect 914 2063 925 2066
rect 890 2053 917 2056
rect 890 2013 893 2053
rect 898 2016 901 2046
rect 906 2023 909 2036
rect 898 2013 909 2016
rect 914 2013 917 2053
rect 882 2005 893 2008
rect 890 1993 893 2005
rect 906 2003 909 2013
rect 922 1996 925 2063
rect 930 2003 933 2016
rect 906 1993 925 1996
rect 874 1933 893 1936
rect 810 1903 821 1906
rect 842 1903 845 1916
rect 862 1913 869 1916
rect 818 1836 821 1903
rect 818 1833 825 1836
rect 802 1823 813 1826
rect 794 1803 797 1816
rect 810 1733 813 1823
rect 822 1746 825 1833
rect 834 1813 837 1836
rect 822 1743 829 1746
rect 786 1703 793 1706
rect 790 1636 793 1703
rect 802 1663 805 1726
rect 810 1723 821 1726
rect 786 1633 793 1636
rect 786 1586 789 1633
rect 794 1603 797 1616
rect 786 1583 793 1586
rect 790 1526 793 1583
rect 802 1543 805 1616
rect 810 1583 813 1706
rect 762 1423 773 1426
rect 754 1326 757 1386
rect 754 1323 765 1326
rect 770 1323 773 1416
rect 730 1303 741 1306
rect 738 1246 741 1303
rect 730 1243 741 1246
rect 730 1153 733 1243
rect 722 1143 733 1146
rect 698 1123 717 1126
rect 686 1063 693 1066
rect 706 1113 717 1116
rect 686 956 689 1063
rect 698 1003 701 1056
rect 706 1023 709 1113
rect 722 1023 725 1136
rect 730 1016 733 1143
rect 706 993 709 1016
rect 722 1013 733 1016
rect 686 953 693 956
rect 690 936 693 953
rect 682 933 693 936
rect 698 926 701 966
rect 706 933 709 946
rect 666 913 677 916
rect 666 846 669 913
rect 666 843 677 846
rect 626 796 629 806
rect 634 803 645 806
rect 658 803 661 826
rect 666 796 669 806
rect 626 793 669 796
rect 650 773 661 776
rect 658 756 661 773
rect 654 753 661 756
rect 618 743 645 746
rect 610 733 637 736
rect 578 703 581 726
rect 586 636 589 726
rect 602 723 629 726
rect 578 633 589 636
rect 562 593 569 596
rect 566 466 569 593
rect 578 546 581 633
rect 586 613 589 626
rect 594 613 605 616
rect 578 543 589 546
rect 594 543 597 613
rect 602 563 605 606
rect 586 536 589 543
rect 610 536 613 626
rect 618 603 621 676
rect 566 463 573 466
rect 546 443 565 446
rect 570 426 573 463
rect 578 433 581 536
rect 586 533 593 536
rect 590 456 593 533
rect 602 533 613 536
rect 590 453 597 456
rect 554 383 557 416
rect 562 413 565 426
rect 570 423 581 426
rect 586 423 589 436
rect 570 366 573 416
rect 578 406 581 423
rect 578 403 585 406
rect 562 363 573 366
rect 530 213 533 336
rect 538 296 541 316
rect 538 293 549 296
rect 546 236 549 293
rect 562 276 565 363
rect 582 356 585 403
rect 578 353 585 356
rect 562 273 573 276
rect 570 253 573 273
rect 538 233 549 236
rect 538 183 541 233
rect 554 176 557 206
rect 442 123 445 136
rect 474 116 477 136
rect 482 123 485 146
rect 490 133 493 176
rect 498 173 525 176
rect 498 123 501 173
rect 506 133 509 166
rect 514 116 517 136
rect 474 113 517 116
rect 522 103 525 173
rect 538 143 541 176
rect 554 173 573 176
rect 554 163 565 166
rect 562 133 565 163
rect 570 143 573 173
rect 578 123 581 353
rect 594 313 597 453
rect 602 413 605 533
rect 610 506 613 526
rect 618 513 621 536
rect 626 506 629 723
rect 634 513 637 733
rect 642 713 645 743
rect 654 656 657 753
rect 654 653 661 656
rect 666 653 669 776
rect 674 723 677 843
rect 682 793 685 926
rect 690 923 701 926
rect 706 873 709 916
rect 722 866 725 1013
rect 738 996 741 1226
rect 746 1173 749 1206
rect 734 993 741 996
rect 734 936 737 993
rect 746 953 749 1156
rect 754 1116 757 1216
rect 762 1203 765 1323
rect 778 1306 781 1526
rect 790 1523 797 1526
rect 786 1423 789 1436
rect 794 1373 797 1523
rect 810 1436 813 1546
rect 818 1486 821 1676
rect 826 1493 829 1743
rect 834 1646 837 1796
rect 842 1693 845 1806
rect 850 1773 853 1846
rect 862 1826 865 1913
rect 858 1823 865 1826
rect 858 1786 861 1823
rect 866 1803 869 1816
rect 858 1783 865 1786
rect 850 1673 853 1746
rect 862 1646 865 1783
rect 834 1643 853 1646
rect 834 1593 837 1606
rect 834 1543 837 1586
rect 834 1513 837 1526
rect 842 1496 845 1616
rect 850 1603 853 1643
rect 858 1643 865 1646
rect 858 1596 861 1643
rect 866 1613 869 1626
rect 838 1493 845 1496
rect 850 1593 861 1596
rect 818 1483 829 1486
rect 802 1433 813 1436
rect 802 1383 805 1433
rect 810 1403 813 1426
rect 826 1423 829 1483
rect 838 1406 841 1493
rect 850 1426 853 1593
rect 858 1483 861 1536
rect 858 1433 869 1436
rect 850 1423 869 1426
rect 826 1403 841 1406
rect 786 1323 789 1336
rect 794 1333 797 1346
rect 826 1336 829 1403
rect 842 1383 845 1396
rect 842 1343 845 1366
rect 826 1333 837 1336
rect 834 1316 837 1333
rect 786 1313 837 1316
rect 774 1303 781 1306
rect 826 1303 837 1306
rect 762 1133 765 1166
rect 774 1146 777 1303
rect 770 1143 777 1146
rect 786 1146 789 1266
rect 802 1193 805 1226
rect 810 1203 813 1236
rect 802 1166 805 1186
rect 802 1163 809 1166
rect 786 1143 797 1146
rect 754 1113 761 1116
rect 758 1036 761 1113
rect 754 1033 761 1036
rect 754 1013 757 1033
rect 734 933 741 936
rect 754 933 757 1006
rect 738 913 741 933
rect 746 903 749 926
rect 714 863 725 866
rect 706 773 709 816
rect 714 763 717 863
rect 754 823 757 836
rect 690 733 717 736
rect 690 723 693 733
rect 642 576 645 616
rect 658 603 661 653
rect 690 583 693 666
rect 706 663 709 726
rect 714 723 717 733
rect 722 673 725 816
rect 762 813 765 1016
rect 770 936 773 1143
rect 778 1133 789 1136
rect 786 1053 789 1126
rect 778 973 781 1006
rect 770 933 781 936
rect 786 933 789 1026
rect 778 926 781 933
rect 770 796 773 926
rect 778 923 789 926
rect 778 863 781 916
rect 762 793 773 796
rect 738 713 741 736
rect 762 726 765 793
rect 778 746 781 806
rect 786 753 789 923
rect 794 906 797 1143
rect 806 986 809 1163
rect 818 1036 821 1126
rect 826 1113 829 1303
rect 842 1203 845 1336
rect 850 1263 853 1356
rect 858 1323 861 1406
rect 866 1333 869 1423
rect 874 1263 877 1916
rect 882 1903 885 1926
rect 882 1803 885 1826
rect 882 1723 885 1736
rect 882 1703 885 1716
rect 890 1636 893 1933
rect 898 1833 901 1946
rect 906 1906 909 1993
rect 922 1926 925 1976
rect 914 1923 925 1926
rect 906 1903 913 1906
rect 910 1846 913 1903
rect 938 1896 941 2066
rect 946 2013 949 2026
rect 946 1993 949 2006
rect 954 1983 957 2006
rect 946 1923 949 1956
rect 938 1893 945 1896
rect 906 1843 913 1846
rect 906 1826 909 1843
rect 906 1823 925 1826
rect 898 1756 901 1816
rect 906 1813 917 1816
rect 906 1783 909 1806
rect 922 1803 925 1823
rect 930 1793 933 1866
rect 942 1826 945 1893
rect 938 1823 945 1826
rect 930 1756 933 1776
rect 898 1753 933 1756
rect 906 1733 917 1736
rect 882 1633 893 1636
rect 882 1363 885 1633
rect 890 1533 893 1616
rect 914 1546 917 1726
rect 930 1616 933 1753
rect 938 1713 941 1823
rect 946 1626 949 1736
rect 954 1716 957 1836
rect 962 1793 965 2073
rect 986 1873 989 2083
rect 1010 2073 1013 2126
rect 1018 2013 1021 2183
rect 1042 2156 1045 2206
rect 1026 2153 1045 2156
rect 1026 2053 1029 2153
rect 1042 2133 1061 2136
rect 1066 2133 1069 2336
rect 1090 2323 1093 2343
rect 1106 2326 1109 2336
rect 1098 2323 1109 2326
rect 1098 2316 1101 2323
rect 1074 2313 1101 2316
rect 1106 2273 1109 2316
rect 1074 2153 1077 2216
rect 1074 2133 1077 2146
rect 1058 2126 1061 2133
rect 1058 2123 1069 2126
rect 1066 2113 1085 2116
rect 1002 1976 1005 2006
rect 1010 1993 1013 2006
rect 1026 1983 1029 2006
rect 1034 1993 1037 2016
rect 1050 2013 1053 2046
rect 1002 1973 1021 1976
rect 1002 1923 1005 1966
rect 970 1783 973 1796
rect 962 1743 981 1746
rect 978 1733 981 1743
rect 986 1733 989 1826
rect 1002 1816 1005 1916
rect 1010 1903 1013 1926
rect 1018 1913 1021 1973
rect 1042 1946 1045 2006
rect 1034 1943 1045 1946
rect 1034 1926 1037 1943
rect 1030 1923 1037 1926
rect 1030 1846 1033 1923
rect 1030 1843 1037 1846
rect 1042 1843 1045 1936
rect 1050 1873 1053 1926
rect 1058 1866 1061 2016
rect 1082 2013 1085 2113
rect 1090 2083 1093 2206
rect 1114 2143 1117 2226
rect 1122 2203 1125 2343
rect 1134 2296 1137 2373
rect 1194 2366 1197 2406
rect 1210 2403 1229 2406
rect 1146 2306 1149 2336
rect 1154 2323 1157 2366
rect 1186 2363 1197 2366
rect 1186 2333 1189 2363
rect 1170 2313 1173 2326
rect 1202 2323 1205 2346
rect 1210 2323 1213 2336
rect 1234 2333 1237 2366
rect 1234 2306 1237 2326
rect 1146 2303 1157 2306
rect 1134 2293 1141 2296
rect 1130 2213 1133 2226
rect 1130 2183 1133 2206
rect 1130 2106 1133 2136
rect 1122 2103 1133 2106
rect 1122 2036 1125 2103
rect 1122 2033 1133 2036
rect 1130 2013 1133 2033
rect 1138 2013 1141 2293
rect 1154 2216 1157 2303
rect 1226 2303 1237 2306
rect 1146 2136 1149 2216
rect 1154 2213 1165 2216
rect 1162 2203 1165 2213
rect 1170 2176 1173 2226
rect 1186 2223 1221 2226
rect 1178 2193 1181 2216
rect 1162 2173 1173 2176
rect 1146 2133 1157 2136
rect 1146 2033 1149 2126
rect 1090 1956 1093 2006
rect 1074 1953 1093 1956
rect 1066 1923 1069 1936
rect 1050 1863 1061 1866
rect 1018 1823 1029 1826
rect 1002 1813 1009 1816
rect 962 1723 981 1726
rect 954 1713 973 1716
rect 970 1696 973 1713
rect 946 1623 957 1626
rect 930 1613 941 1616
rect 922 1593 933 1596
rect 906 1543 917 1546
rect 890 1493 893 1526
rect 906 1446 909 1543
rect 914 1516 917 1536
rect 930 1533 933 1593
rect 914 1513 925 1516
rect 898 1443 909 1446
rect 890 1373 893 1426
rect 890 1313 893 1346
rect 850 1213 853 1236
rect 818 1033 829 1036
rect 802 983 809 986
rect 802 963 805 983
rect 818 936 821 1016
rect 826 1003 829 1033
rect 810 933 821 936
rect 810 926 813 933
rect 802 923 813 926
rect 794 903 805 906
rect 818 903 821 926
rect 802 826 805 903
rect 826 876 829 936
rect 794 823 805 826
rect 818 873 829 876
rect 818 826 821 873
rect 818 823 829 826
rect 778 743 789 746
rect 746 723 765 726
rect 746 656 749 723
rect 706 653 749 656
rect 706 613 709 653
rect 722 613 765 616
rect 642 573 649 576
rect 646 506 649 573
rect 674 533 709 536
rect 674 526 677 533
rect 666 523 677 526
rect 658 513 669 516
rect 610 503 629 506
rect 642 503 649 506
rect 642 423 645 503
rect 610 376 613 416
rect 658 413 661 456
rect 666 436 669 506
rect 682 453 685 526
rect 706 523 709 533
rect 690 513 701 516
rect 666 433 685 436
rect 674 406 677 426
rect 682 413 685 433
rect 618 403 677 406
rect 682 376 685 406
rect 602 373 613 376
rect 602 333 605 373
rect 610 333 621 336
rect 610 273 613 326
rect 626 323 629 376
rect 666 373 685 376
rect 666 343 669 373
rect 682 353 685 373
rect 690 306 693 326
rect 682 303 693 306
rect 586 223 589 236
rect 594 226 597 236
rect 602 233 605 266
rect 682 246 685 303
rect 682 243 693 246
rect 594 223 613 226
rect 594 206 597 216
rect 618 206 621 236
rect 594 203 621 206
rect 650 196 653 216
rect 642 193 653 196
rect 666 193 669 226
rect 682 203 685 226
rect 594 133 597 186
rect 634 116 637 126
rect 642 123 645 193
rect 690 183 693 243
rect 658 123 661 136
rect 666 116 669 176
rect 698 123 701 376
rect 714 333 717 386
rect 706 213 709 286
rect 722 216 725 613
rect 738 533 741 606
rect 746 473 749 526
rect 730 403 733 416
rect 738 403 741 436
rect 738 333 741 356
rect 730 223 733 236
rect 738 226 741 316
rect 746 253 749 456
rect 762 413 765 586
rect 770 533 773 676
rect 778 623 781 736
rect 770 513 773 526
rect 778 423 781 616
rect 786 613 789 743
rect 794 663 797 823
rect 826 806 829 823
rect 834 813 837 1106
rect 842 1003 845 1116
rect 850 1113 853 1126
rect 850 986 853 1076
rect 846 983 853 986
rect 846 846 849 983
rect 846 843 853 846
rect 802 803 829 806
rect 802 726 805 803
rect 802 723 821 726
rect 794 556 797 656
rect 802 613 805 716
rect 810 683 813 716
rect 818 686 821 706
rect 818 683 829 686
rect 810 606 813 666
rect 826 636 829 683
rect 842 643 845 826
rect 850 716 853 843
rect 858 836 861 1206
rect 866 1173 869 1216
rect 890 1186 893 1226
rect 898 1206 901 1443
rect 922 1436 925 1513
rect 906 1336 909 1436
rect 918 1433 925 1436
rect 918 1346 921 1433
rect 938 1426 941 1613
rect 954 1563 957 1606
rect 962 1603 965 1696
rect 970 1693 981 1696
rect 978 1646 981 1693
rect 994 1653 997 1806
rect 1006 1756 1009 1813
rect 1034 1806 1037 1843
rect 1018 1803 1037 1806
rect 1050 1803 1053 1863
rect 1066 1813 1069 1846
rect 1006 1753 1013 1756
rect 1002 1733 1005 1746
rect 970 1643 981 1646
rect 970 1613 973 1643
rect 1002 1606 1005 1726
rect 1010 1633 1013 1753
rect 1018 1716 1021 1803
rect 1026 1733 1029 1786
rect 1034 1753 1037 1796
rect 1034 1733 1045 1736
rect 1018 1713 1029 1716
rect 994 1603 1005 1606
rect 946 1513 949 1536
rect 954 1516 957 1546
rect 994 1543 997 1556
rect 1010 1526 1013 1606
rect 1026 1566 1029 1713
rect 1042 1596 1045 1733
rect 1050 1723 1053 1766
rect 1058 1706 1061 1736
rect 1050 1703 1061 1706
rect 1066 1693 1069 1796
rect 1074 1673 1077 1953
rect 1082 1913 1085 1946
rect 1082 1756 1085 1876
rect 1090 1803 1093 1906
rect 1098 1843 1101 1936
rect 1082 1753 1093 1756
rect 1082 1733 1085 1746
rect 1090 1666 1093 1753
rect 1098 1716 1101 1726
rect 1106 1723 1109 1926
rect 1114 1803 1117 2006
rect 1122 1913 1125 1946
rect 1154 1936 1157 2133
rect 1162 2063 1165 2173
rect 1162 2003 1165 2016
rect 1130 1876 1133 1926
rect 1138 1923 1141 1936
rect 1146 1933 1157 1936
rect 1122 1873 1133 1876
rect 1122 1813 1125 1873
rect 1138 1813 1141 1826
rect 1130 1803 1141 1806
rect 1114 1716 1117 1726
rect 1122 1723 1125 1736
rect 1130 1733 1133 1756
rect 1138 1733 1141 1746
rect 1098 1713 1117 1716
rect 1086 1663 1093 1666
rect 1018 1563 1029 1566
rect 1038 1593 1045 1596
rect 1018 1533 1021 1563
rect 1038 1546 1041 1593
rect 1026 1543 1041 1546
rect 954 1513 965 1516
rect 962 1426 965 1513
rect 994 1486 997 1526
rect 938 1423 945 1426
rect 930 1383 933 1416
rect 942 1376 945 1423
rect 938 1373 945 1376
rect 954 1423 965 1426
rect 986 1483 997 1486
rect 986 1426 989 1483
rect 1002 1453 1005 1526
rect 1010 1523 1017 1526
rect 1014 1466 1017 1523
rect 1014 1463 1021 1466
rect 986 1423 1005 1426
rect 938 1353 941 1373
rect 918 1343 925 1346
rect 906 1333 917 1336
rect 906 1223 909 1326
rect 914 1213 917 1333
rect 922 1286 925 1343
rect 930 1306 933 1336
rect 938 1333 941 1346
rect 946 1326 949 1346
rect 954 1333 957 1423
rect 946 1323 957 1326
rect 962 1323 965 1336
rect 930 1303 941 1306
rect 922 1283 929 1286
rect 926 1206 929 1283
rect 898 1203 905 1206
rect 882 1183 893 1186
rect 882 1136 885 1183
rect 866 1113 869 1136
rect 882 1133 893 1136
rect 874 1063 877 1106
rect 882 1103 885 1116
rect 866 896 869 1056
rect 882 1026 885 1086
rect 890 1053 893 1133
rect 902 1066 905 1203
rect 914 1113 917 1206
rect 922 1203 929 1206
rect 898 1063 905 1066
rect 898 1043 901 1063
rect 874 1023 885 1026
rect 890 1026 893 1036
rect 898 1033 917 1036
rect 890 1023 909 1026
rect 874 1006 877 1023
rect 874 1003 881 1006
rect 890 1003 893 1016
rect 914 1003 917 1033
rect 878 946 881 1003
rect 890 983 909 986
rect 878 943 885 946
rect 874 906 877 926
rect 882 913 885 943
rect 890 933 893 983
rect 898 926 901 976
rect 906 966 909 983
rect 906 963 913 966
rect 890 923 901 926
rect 910 916 913 963
rect 906 913 913 916
rect 874 903 893 906
rect 866 893 877 896
rect 858 833 869 836
rect 858 803 861 833
rect 866 783 869 816
rect 850 713 869 716
rect 818 633 829 636
rect 818 613 821 633
rect 786 553 797 556
rect 786 446 789 553
rect 794 533 797 546
rect 794 463 797 526
rect 786 443 793 446
rect 770 403 773 416
rect 770 306 773 366
rect 762 303 773 306
rect 762 246 765 303
rect 762 243 773 246
rect 738 223 757 226
rect 722 213 741 216
rect 738 203 741 213
rect 770 173 773 243
rect 778 233 781 406
rect 790 356 793 443
rect 802 403 805 606
rect 810 603 821 606
rect 810 396 813 536
rect 818 473 821 603
rect 826 533 829 616
rect 850 603 853 686
rect 866 616 869 713
rect 874 706 877 893
rect 890 836 893 903
rect 882 833 893 836
rect 882 813 885 833
rect 882 783 885 806
rect 890 723 893 796
rect 898 733 901 756
rect 906 723 909 913
rect 922 823 925 1203
rect 938 1186 941 1303
rect 954 1213 957 1236
rect 930 1183 941 1186
rect 930 1116 933 1183
rect 938 1133 941 1166
rect 930 1113 937 1116
rect 934 1006 937 1113
rect 930 1003 937 1006
rect 930 983 933 1003
rect 930 933 933 946
rect 930 903 933 926
rect 938 923 941 936
rect 946 906 949 1126
rect 954 1113 957 1206
rect 962 1143 965 1226
rect 970 1206 973 1406
rect 986 1396 989 1406
rect 978 1393 989 1396
rect 994 1376 997 1416
rect 986 1373 997 1376
rect 986 1306 989 1373
rect 1002 1313 1005 1423
rect 1010 1413 1013 1446
rect 986 1303 997 1306
rect 970 1203 981 1206
rect 978 1136 981 1203
rect 970 1133 981 1136
rect 962 1076 965 1126
rect 970 1096 973 1133
rect 994 1123 997 1303
rect 1018 1226 1021 1463
rect 1026 1383 1029 1543
rect 1050 1533 1053 1586
rect 1058 1493 1061 1526
rect 1034 1366 1037 1476
rect 1066 1436 1069 1536
rect 1074 1513 1077 1606
rect 1086 1586 1089 1663
rect 1098 1623 1101 1706
rect 1098 1586 1101 1606
rect 1114 1603 1117 1696
rect 1130 1646 1133 1726
rect 1146 1703 1149 1933
rect 1154 1913 1157 1926
rect 1162 1916 1165 1946
rect 1170 1926 1173 2126
rect 1178 2106 1181 2136
rect 1186 2123 1189 2223
rect 1194 2173 1197 2206
rect 1226 2203 1229 2303
rect 1242 2256 1245 2416
rect 1266 2346 1269 2406
rect 1274 2373 1277 2416
rect 1266 2343 1293 2346
rect 1298 2343 1301 2426
rect 1330 2423 1349 2426
rect 1330 2413 1333 2423
rect 1346 2416 1349 2423
rect 1330 2353 1333 2406
rect 1338 2363 1341 2416
rect 1346 2413 1357 2416
rect 1354 2373 1357 2406
rect 1266 2323 1269 2336
rect 1282 2326 1285 2336
rect 1274 2323 1285 2326
rect 1290 2326 1293 2343
rect 1290 2323 1301 2326
rect 1274 2316 1277 2323
rect 1250 2313 1277 2316
rect 1282 2273 1285 2316
rect 1298 2266 1301 2323
rect 1290 2263 1301 2266
rect 1242 2253 1253 2256
rect 1234 2183 1237 2206
rect 1250 2186 1253 2253
rect 1266 2213 1285 2216
rect 1242 2183 1253 2186
rect 1194 2136 1197 2146
rect 1194 2133 1213 2136
rect 1234 2133 1237 2146
rect 1194 2123 1205 2126
rect 1210 2116 1213 2133
rect 1202 2113 1213 2116
rect 1178 2103 1185 2106
rect 1182 2026 1185 2103
rect 1182 2023 1189 2026
rect 1178 1996 1181 2016
rect 1186 2003 1189 2023
rect 1194 2013 1197 2066
rect 1202 2003 1205 2113
rect 1210 2013 1213 2046
rect 1178 1993 1217 1996
rect 1170 1923 1181 1926
rect 1162 1913 1173 1916
rect 1154 1813 1157 1866
rect 1162 1753 1165 1826
rect 1170 1746 1173 1846
rect 1178 1803 1181 1923
rect 1194 1803 1197 1956
rect 1202 1923 1205 1966
rect 1214 1936 1217 1993
rect 1214 1933 1221 1936
rect 1202 1913 1213 1916
rect 1218 1913 1221 1933
rect 1226 1903 1229 2006
rect 1234 1983 1237 2126
rect 1242 2106 1245 2183
rect 1250 2123 1253 2136
rect 1258 2133 1261 2166
rect 1266 2133 1269 2146
rect 1258 2123 1269 2126
rect 1242 2103 1253 2106
rect 1250 2046 1253 2103
rect 1242 2043 1253 2046
rect 1242 2013 1245 2043
rect 1274 2026 1277 2213
rect 1290 2203 1293 2263
rect 1314 2226 1317 2336
rect 1322 2323 1325 2346
rect 1362 2333 1365 2426
rect 1394 2403 1397 2416
rect 1402 2403 1405 2446
rect 1410 2346 1413 2416
rect 1442 2393 1445 2406
rect 1466 2403 1469 2416
rect 1522 2413 1525 2446
rect 1554 2413 1589 2416
rect 1370 2343 1413 2346
rect 1370 2326 1373 2343
rect 1362 2323 1373 2326
rect 1378 2323 1381 2336
rect 1394 2333 1405 2336
rect 1386 2323 1405 2326
rect 1338 2273 1341 2316
rect 1298 2186 1301 2226
rect 1314 2223 1325 2226
rect 1322 2216 1325 2223
rect 1322 2213 1333 2216
rect 1306 2193 1309 2206
rect 1330 2203 1333 2213
rect 1298 2183 1317 2186
rect 1298 2093 1301 2126
rect 1314 2123 1317 2183
rect 1322 2133 1325 2186
rect 1338 2133 1341 2226
rect 1362 2216 1365 2323
rect 1386 2303 1389 2323
rect 1362 2213 1373 2216
rect 1258 2023 1277 2026
rect 1242 1976 1245 1996
rect 1242 1973 1249 1976
rect 1234 1913 1237 1956
rect 1210 1813 1213 1826
rect 1234 1813 1237 1906
rect 1246 1876 1249 1973
rect 1242 1873 1249 1876
rect 1242 1853 1245 1873
rect 1202 1803 1213 1806
rect 1162 1743 1173 1746
rect 1162 1733 1165 1743
rect 1122 1643 1133 1646
rect 1086 1583 1093 1586
rect 1098 1583 1105 1586
rect 1058 1433 1069 1436
rect 1030 1363 1037 1366
rect 1030 1256 1033 1363
rect 1030 1253 1037 1256
rect 1034 1233 1037 1253
rect 1002 1206 1005 1226
rect 1018 1223 1037 1226
rect 1002 1203 1013 1206
rect 1010 1136 1013 1203
rect 1002 1133 1013 1136
rect 1026 1133 1029 1186
rect 978 1106 981 1116
rect 978 1103 997 1106
rect 970 1093 989 1096
rect 954 1073 965 1076
rect 954 1013 957 1073
rect 962 1016 965 1026
rect 962 1013 973 1016
rect 978 1006 981 1046
rect 954 933 957 1006
rect 962 953 965 1006
rect 974 1003 981 1006
rect 942 903 949 906
rect 954 903 957 916
rect 942 826 945 903
rect 954 836 957 886
rect 962 843 965 946
rect 954 833 965 836
rect 942 823 949 826
rect 938 793 941 806
rect 914 713 917 776
rect 946 726 949 823
rect 954 796 957 816
rect 962 813 965 833
rect 974 826 977 1003
rect 970 823 977 826
rect 954 793 965 796
rect 970 753 973 823
rect 978 743 981 806
rect 986 773 989 1093
rect 994 1013 997 1103
rect 1002 1083 1005 1133
rect 1010 1103 1013 1116
rect 1002 983 1005 1006
rect 994 933 997 956
rect 1010 936 1013 1006
rect 1002 933 1013 936
rect 994 906 997 926
rect 994 903 1005 906
rect 1002 846 1005 903
rect 994 843 1005 846
rect 994 813 997 843
rect 1002 813 1005 826
rect 994 763 997 806
rect 874 703 893 706
rect 866 613 877 616
rect 866 546 869 606
rect 882 603 885 626
rect 890 603 893 703
rect 922 686 925 726
rect 906 683 925 686
rect 938 723 949 726
rect 1002 723 1005 796
rect 1018 776 1021 1116
rect 1026 1003 1029 1126
rect 1034 926 1037 1223
rect 1042 1013 1045 1406
rect 1050 1403 1053 1426
rect 1058 1413 1061 1433
rect 1074 1426 1077 1436
rect 1066 1423 1077 1426
rect 1082 1423 1085 1566
rect 1090 1533 1093 1583
rect 1050 1333 1053 1356
rect 1066 1336 1069 1423
rect 1074 1413 1085 1416
rect 1090 1406 1093 1516
rect 1102 1496 1105 1583
rect 1082 1403 1093 1406
rect 1098 1493 1105 1496
rect 1098 1403 1101 1493
rect 1082 1393 1085 1403
rect 1058 1333 1069 1336
rect 1058 1306 1061 1333
rect 1050 1303 1061 1306
rect 1066 1306 1069 1326
rect 1066 1303 1073 1306
rect 1050 1183 1053 1303
rect 1058 1213 1061 1296
rect 1070 1196 1073 1303
rect 1066 1193 1073 1196
rect 1066 1173 1069 1193
rect 1050 1063 1053 1126
rect 1058 1083 1061 1116
rect 1026 923 1037 926
rect 1042 906 1045 1006
rect 1034 903 1045 906
rect 1034 846 1037 903
rect 1034 843 1045 846
rect 1034 803 1037 816
rect 1018 773 1025 776
rect 858 543 869 546
rect 810 393 821 396
rect 826 383 829 416
rect 834 413 837 486
rect 842 463 845 526
rect 850 513 853 536
rect 858 493 861 543
rect 866 416 869 536
rect 882 533 885 566
rect 874 473 877 526
rect 890 523 893 546
rect 866 413 885 416
rect 786 353 793 356
rect 786 163 789 353
rect 794 306 797 336
rect 810 333 837 336
rect 810 323 813 333
rect 826 313 829 326
rect 834 313 837 333
rect 850 306 853 356
rect 866 323 869 406
rect 882 393 885 413
rect 794 303 829 306
rect 826 286 829 303
rect 818 283 829 286
rect 818 236 821 283
rect 794 213 797 236
rect 818 233 829 236
rect 826 213 829 233
rect 834 216 837 306
rect 850 303 861 306
rect 858 236 861 303
rect 882 296 885 316
rect 874 293 885 296
rect 874 246 877 293
rect 890 286 893 346
rect 906 323 909 683
rect 938 623 941 723
rect 946 713 965 716
rect 962 643 965 713
rect 1010 646 1013 766
rect 1022 696 1025 773
rect 1018 693 1025 696
rect 1018 673 1021 693
rect 1034 673 1037 796
rect 1042 733 1045 843
rect 1050 813 1053 1036
rect 1058 973 1061 1026
rect 1066 1003 1069 1136
rect 1058 893 1061 936
rect 1066 933 1069 996
rect 1058 766 1061 866
rect 1066 793 1069 926
rect 1074 846 1077 1106
rect 1082 923 1085 1356
rect 1090 1333 1093 1366
rect 1098 1323 1101 1396
rect 1090 1223 1093 1256
rect 1106 1223 1109 1446
rect 1114 1313 1117 1526
rect 1122 1433 1125 1643
rect 1122 1313 1125 1396
rect 1130 1353 1133 1636
rect 1146 1533 1149 1616
rect 1162 1603 1165 1646
rect 1178 1626 1181 1756
rect 1202 1746 1205 1803
rect 1218 1793 1221 1806
rect 1250 1803 1253 1826
rect 1258 1786 1261 2023
rect 1266 2013 1277 2016
rect 1282 2003 1285 2046
rect 1330 2043 1333 2126
rect 1346 2116 1349 2196
rect 1354 2193 1357 2206
rect 1342 2113 1349 2116
rect 1322 2013 1325 2036
rect 1342 2016 1345 2113
rect 1354 2103 1357 2166
rect 1370 2146 1373 2213
rect 1386 2196 1389 2296
rect 1394 2203 1397 2323
rect 1402 2293 1405 2316
rect 1418 2276 1421 2356
rect 1442 2333 1445 2346
rect 1418 2273 1425 2276
rect 1386 2193 1397 2196
rect 1362 2143 1373 2146
rect 1362 2123 1365 2143
rect 1386 2133 1389 2156
rect 1394 2116 1397 2193
rect 1402 2173 1405 2216
rect 1410 2166 1413 2266
rect 1422 2226 1425 2273
rect 1370 2113 1381 2116
rect 1390 2113 1397 2116
rect 1402 2163 1413 2166
rect 1418 2223 1425 2226
rect 1370 2106 1373 2113
rect 1362 2103 1373 2106
rect 1330 2013 1345 2016
rect 1330 2006 1333 2013
rect 1354 2006 1357 2056
rect 1322 2003 1333 2006
rect 1282 1973 1285 1996
rect 1290 1936 1293 1946
rect 1282 1906 1285 1936
rect 1290 1933 1301 1936
rect 1290 1913 1293 1926
rect 1266 1903 1285 1906
rect 1298 1876 1301 1933
rect 1306 1923 1309 1996
rect 1314 1903 1317 1926
rect 1294 1873 1301 1876
rect 1294 1826 1297 1873
rect 1294 1823 1301 1826
rect 1274 1813 1285 1816
rect 1266 1803 1277 1806
rect 1298 1803 1301 1823
rect 1306 1803 1309 1866
rect 1242 1773 1245 1786
rect 1258 1783 1285 1786
rect 1186 1743 1205 1746
rect 1226 1763 1261 1766
rect 1186 1723 1189 1743
rect 1226 1736 1229 1763
rect 1194 1733 1229 1736
rect 1170 1623 1181 1626
rect 1170 1596 1173 1623
rect 1162 1593 1173 1596
rect 1138 1496 1141 1526
rect 1138 1493 1149 1496
rect 1138 1423 1141 1493
rect 1154 1436 1157 1536
rect 1162 1523 1165 1593
rect 1170 1533 1173 1566
rect 1178 1546 1181 1616
rect 1202 1593 1205 1726
rect 1210 1723 1221 1726
rect 1226 1646 1229 1733
rect 1234 1723 1237 1756
rect 1250 1733 1253 1756
rect 1258 1733 1261 1763
rect 1226 1643 1237 1646
rect 1234 1623 1237 1643
rect 1218 1556 1221 1606
rect 1218 1553 1229 1556
rect 1178 1543 1221 1546
rect 1178 1526 1181 1543
rect 1194 1533 1205 1536
rect 1218 1533 1221 1543
rect 1178 1523 1185 1526
rect 1150 1433 1157 1436
rect 1138 1363 1141 1416
rect 1150 1356 1153 1433
rect 1138 1353 1153 1356
rect 1098 1213 1109 1216
rect 1114 1213 1117 1246
rect 1090 1163 1093 1206
rect 1090 1053 1093 1136
rect 1098 1046 1101 1186
rect 1106 1113 1109 1206
rect 1122 1203 1125 1226
rect 1130 1173 1133 1326
rect 1138 1286 1141 1353
rect 1162 1336 1165 1426
rect 1170 1403 1173 1486
rect 1182 1416 1185 1523
rect 1178 1413 1185 1416
rect 1194 1416 1197 1526
rect 1210 1493 1213 1526
rect 1226 1426 1229 1553
rect 1242 1523 1245 1706
rect 1250 1653 1253 1726
rect 1258 1713 1261 1726
rect 1258 1636 1261 1706
rect 1254 1633 1261 1636
rect 1254 1556 1257 1633
rect 1266 1613 1269 1736
rect 1282 1716 1285 1783
rect 1298 1723 1301 1796
rect 1278 1713 1285 1716
rect 1278 1646 1281 1713
rect 1274 1643 1281 1646
rect 1274 1613 1277 1643
rect 1254 1553 1261 1556
rect 1250 1506 1253 1536
rect 1242 1503 1253 1506
rect 1242 1436 1245 1503
rect 1242 1433 1253 1436
rect 1210 1423 1229 1426
rect 1194 1413 1205 1416
rect 1178 1336 1181 1413
rect 1146 1333 1173 1336
rect 1178 1333 1189 1336
rect 1194 1333 1197 1396
rect 1146 1306 1149 1333
rect 1154 1323 1181 1326
rect 1178 1306 1181 1323
rect 1146 1303 1157 1306
rect 1138 1283 1145 1286
rect 1142 1226 1145 1283
rect 1138 1223 1145 1226
rect 1130 1136 1133 1156
rect 1122 1133 1133 1136
rect 1090 1043 1101 1046
rect 1122 1046 1125 1133
rect 1122 1043 1133 1046
rect 1082 856 1085 916
rect 1090 883 1093 1043
rect 1122 1003 1125 1026
rect 1130 1003 1133 1043
rect 1098 923 1101 976
rect 1114 933 1117 956
rect 1114 856 1117 916
rect 1082 853 1117 856
rect 1074 843 1093 846
rect 1050 763 1061 766
rect 1050 746 1053 763
rect 1074 756 1077 816
rect 1082 813 1085 836
rect 1090 766 1093 843
rect 1098 813 1101 853
rect 1122 846 1125 996
rect 1138 973 1141 1223
rect 1154 1206 1157 1303
rect 1146 1203 1157 1206
rect 1170 1303 1181 1306
rect 1146 1183 1149 1203
rect 1170 1196 1173 1303
rect 1186 1203 1189 1333
rect 1170 1193 1181 1196
rect 1178 1136 1181 1193
rect 1194 1183 1197 1226
rect 1202 1146 1205 1406
rect 1210 1363 1213 1423
rect 1218 1413 1245 1416
rect 1234 1356 1237 1406
rect 1226 1353 1237 1356
rect 1210 1313 1213 1326
rect 1226 1246 1229 1353
rect 1250 1346 1253 1433
rect 1258 1423 1261 1553
rect 1266 1493 1269 1606
rect 1282 1586 1285 1626
rect 1290 1596 1293 1696
rect 1298 1613 1301 1716
rect 1314 1703 1317 1736
rect 1322 1686 1325 2003
rect 1338 1993 1341 2006
rect 1346 2003 1357 2006
rect 1338 1913 1341 1926
rect 1346 1923 1349 2003
rect 1330 1813 1333 1826
rect 1338 1733 1341 1886
rect 1346 1783 1349 1826
rect 1354 1803 1357 1986
rect 1314 1683 1325 1686
rect 1314 1606 1317 1683
rect 1314 1603 1325 1606
rect 1290 1593 1297 1596
rect 1274 1583 1285 1586
rect 1274 1443 1277 1583
rect 1210 1243 1229 1246
rect 1238 1343 1253 1346
rect 1210 1203 1213 1243
rect 1218 1193 1221 1226
rect 1226 1153 1229 1236
rect 1198 1143 1205 1146
rect 1146 1043 1149 1136
rect 1178 1133 1189 1136
rect 1130 933 1141 936
rect 1130 876 1133 933
rect 1146 893 1149 926
rect 1154 903 1157 1126
rect 1162 1113 1165 1126
rect 1170 1103 1173 1126
rect 1186 1076 1189 1133
rect 1178 1073 1189 1076
rect 1178 1056 1181 1073
rect 1162 1053 1189 1056
rect 1162 1013 1165 1053
rect 1186 1013 1189 1053
rect 1198 1016 1201 1143
rect 1238 1136 1241 1343
rect 1258 1336 1261 1406
rect 1250 1333 1261 1336
rect 1266 1313 1269 1326
rect 1194 1013 1201 1016
rect 1162 916 1165 946
rect 1170 933 1173 966
rect 1162 913 1169 916
rect 1130 873 1141 876
rect 1106 843 1125 846
rect 1090 763 1097 766
rect 1074 753 1085 756
rect 1050 743 1069 746
rect 1042 703 1045 726
rect 1066 666 1069 726
rect 1034 663 1069 666
rect 1010 643 1017 646
rect 978 633 989 636
rect 930 596 933 616
rect 922 593 933 596
rect 922 546 925 593
rect 938 583 941 606
rect 922 543 933 546
rect 922 513 925 526
rect 930 463 933 543
rect 938 496 941 566
rect 946 516 949 616
rect 954 523 957 606
rect 986 603 989 633
rect 1014 596 1017 643
rect 1010 593 1017 596
rect 946 513 957 516
rect 938 493 949 496
rect 922 353 925 416
rect 914 343 933 346
rect 890 283 901 286
rect 874 243 885 246
rect 850 233 861 236
rect 834 213 845 216
rect 850 213 853 233
rect 882 223 885 243
rect 898 226 901 283
rect 890 223 901 226
rect 914 223 917 343
rect 922 306 925 336
rect 930 323 933 343
rect 938 313 941 336
rect 922 303 941 306
rect 946 303 949 493
rect 954 473 957 513
rect 962 433 965 536
rect 970 463 973 556
rect 810 203 821 206
rect 834 203 837 213
rect 738 123 741 136
rect 634 113 669 116
rect 786 113 789 126
rect 818 123 821 203
rect 826 173 829 196
rect 834 143 837 196
rect 874 193 877 206
rect 890 203 893 223
rect 930 203 933 266
rect 946 213 949 236
rect 858 123 861 166
rect 866 123 869 146
rect 898 133 901 176
rect 922 143 925 196
rect 938 163 941 206
rect 906 103 909 126
rect 954 123 957 326
rect 962 313 965 426
rect 978 403 981 536
rect 994 533 997 546
rect 1010 526 1013 593
rect 986 473 989 526
rect 1002 523 1013 526
rect 1026 526 1029 656
rect 1034 613 1037 663
rect 1066 626 1069 646
rect 1058 623 1069 626
rect 1058 566 1061 623
rect 1074 593 1077 746
rect 1082 613 1085 753
rect 1094 686 1097 763
rect 1090 683 1097 686
rect 1090 603 1093 683
rect 1106 676 1109 843
rect 1114 803 1117 826
rect 1138 816 1141 873
rect 1130 813 1141 816
rect 1122 776 1125 806
rect 1130 783 1133 813
rect 1154 803 1157 886
rect 1166 836 1169 913
rect 1162 833 1169 836
rect 1162 813 1165 833
rect 1138 793 1165 796
rect 1138 776 1141 793
rect 1122 773 1141 776
rect 1106 673 1113 676
rect 1058 563 1069 566
rect 1066 546 1069 563
rect 1066 543 1077 546
rect 1034 533 1085 536
rect 1026 523 1037 526
rect 1002 446 1005 523
rect 994 443 1005 446
rect 970 393 989 396
rect 994 373 997 443
rect 1010 403 1013 416
rect 1018 403 1021 426
rect 1026 396 1029 406
rect 1010 393 1029 396
rect 1034 386 1037 523
rect 1050 473 1053 526
rect 1066 513 1077 516
rect 1082 513 1085 533
rect 1090 513 1093 576
rect 1098 563 1101 666
rect 1110 626 1113 673
rect 1106 623 1113 626
rect 1106 523 1109 623
rect 1122 613 1125 773
rect 1138 733 1141 746
rect 1146 733 1149 786
rect 1162 733 1165 793
rect 1130 663 1133 726
rect 1154 723 1165 726
rect 1154 706 1157 723
rect 1146 703 1157 706
rect 1146 636 1149 703
rect 1146 633 1157 636
rect 1162 633 1165 716
rect 1114 603 1125 606
rect 1114 513 1117 603
rect 1146 596 1149 616
rect 1122 593 1149 596
rect 1122 523 1125 546
rect 1058 503 1093 506
rect 1018 383 1037 386
rect 1050 386 1053 416
rect 1058 413 1061 503
rect 1066 403 1069 416
rect 1074 413 1077 446
rect 1050 383 1061 386
rect 994 336 997 356
rect 986 333 997 336
rect 1002 333 1013 336
rect 986 226 989 333
rect 986 223 997 226
rect 994 206 997 223
rect 1010 213 1013 326
rect 1018 323 1021 383
rect 1042 336 1045 346
rect 1034 333 1045 336
rect 1018 283 1021 316
rect 1034 276 1037 333
rect 1026 273 1037 276
rect 986 193 989 206
rect 994 203 1005 206
rect 970 143 973 176
rect 994 123 997 166
rect 1026 133 1029 273
rect 1050 223 1053 336
rect 1058 323 1061 383
rect 1098 346 1101 406
rect 1106 363 1109 466
rect 1114 403 1117 476
rect 1130 443 1133 476
rect 1138 403 1141 516
rect 1082 343 1101 346
rect 1082 213 1085 336
rect 1106 213 1109 356
rect 1122 323 1133 326
rect 1138 303 1141 326
rect 1146 286 1149 593
rect 1138 283 1149 286
rect 1114 213 1117 266
rect 1138 206 1141 283
rect 1042 193 1045 206
rect 1090 176 1093 206
rect 1106 193 1109 206
rect 1138 203 1149 206
rect 1146 183 1149 203
rect 1090 173 1149 176
rect 1154 173 1157 633
rect 1170 603 1173 746
rect 1170 543 1173 566
rect 1162 516 1165 536
rect 1162 513 1169 516
rect 1166 406 1169 513
rect 1178 463 1181 1006
rect 1194 926 1197 1013
rect 1202 993 1205 1006
rect 1210 1003 1213 1136
rect 1234 1133 1241 1136
rect 1226 1103 1229 1126
rect 1234 1113 1237 1133
rect 1218 1013 1221 1026
rect 1250 1016 1253 1276
rect 1258 1213 1261 1246
rect 1274 1223 1277 1366
rect 1282 1206 1285 1536
rect 1294 1436 1297 1593
rect 1306 1506 1309 1586
rect 1314 1513 1317 1536
rect 1306 1503 1317 1506
rect 1294 1433 1309 1436
rect 1290 1423 1301 1426
rect 1306 1416 1309 1433
rect 1290 1413 1309 1416
rect 1290 1343 1293 1413
rect 1314 1406 1317 1503
rect 1298 1403 1317 1406
rect 1290 1293 1293 1326
rect 1290 1213 1293 1276
rect 1266 1203 1285 1206
rect 1266 1133 1269 1203
rect 1282 1126 1285 1176
rect 1290 1163 1293 1206
rect 1282 1123 1293 1126
rect 1282 1093 1285 1116
rect 1282 1023 1285 1066
rect 1242 1013 1253 1016
rect 1242 956 1245 1013
rect 1242 953 1253 956
rect 1186 923 1197 926
rect 1202 923 1205 936
rect 1210 933 1229 936
rect 1234 933 1245 936
rect 1186 883 1189 923
rect 1210 916 1213 933
rect 1234 926 1237 933
rect 1226 923 1237 926
rect 1194 913 1213 916
rect 1186 803 1189 816
rect 1186 623 1189 756
rect 1194 733 1197 826
rect 1202 803 1205 816
rect 1210 736 1213 856
rect 1250 853 1253 953
rect 1258 906 1261 1006
rect 1290 993 1293 1123
rect 1298 996 1301 1403
rect 1306 1266 1309 1316
rect 1314 1283 1317 1336
rect 1322 1333 1325 1603
rect 1330 1433 1333 1726
rect 1354 1723 1357 1796
rect 1362 1746 1365 2103
rect 1370 2076 1373 2096
rect 1370 2073 1381 2076
rect 1378 2026 1381 2073
rect 1390 2036 1393 2113
rect 1390 2033 1397 2036
rect 1370 2023 1381 2026
rect 1370 1913 1373 2023
rect 1394 2013 1397 2033
rect 1402 2013 1405 2163
rect 1410 2113 1413 2126
rect 1418 2036 1421 2223
rect 1426 2123 1429 2206
rect 1418 2033 1425 2036
rect 1378 2003 1397 2006
rect 1378 1993 1381 2003
rect 1410 1943 1413 2026
rect 1422 1956 1425 2033
rect 1434 2013 1437 2326
rect 1442 2313 1445 2326
rect 1482 2303 1485 2316
rect 1498 2266 1501 2336
rect 1506 2293 1509 2326
rect 1498 2263 1505 2266
rect 1458 2213 1469 2216
rect 1442 2123 1445 2176
rect 1450 2116 1453 2206
rect 1458 2193 1461 2206
rect 1474 2133 1477 2246
rect 1482 2213 1485 2226
rect 1490 2213 1493 2256
rect 1502 2206 1505 2263
rect 1498 2203 1505 2206
rect 1498 2183 1501 2203
rect 1514 2193 1517 2336
rect 1522 2223 1525 2326
rect 1530 2313 1533 2326
rect 1546 2296 1549 2336
rect 1538 2293 1549 2296
rect 1538 2226 1541 2293
rect 1538 2223 1549 2226
rect 1546 2176 1549 2223
rect 1522 2173 1549 2176
rect 1482 2133 1493 2136
rect 1450 2113 1461 2116
rect 1458 2056 1461 2113
rect 1450 2053 1461 2056
rect 1450 2033 1453 2053
rect 1418 1953 1425 1956
rect 1370 1813 1373 1876
rect 1378 1803 1381 1936
rect 1394 1836 1397 1926
rect 1402 1903 1405 1916
rect 1410 1913 1413 1926
rect 1386 1833 1397 1836
rect 1362 1743 1373 1746
rect 1338 1633 1341 1716
rect 1338 1613 1341 1626
rect 1330 1396 1333 1426
rect 1338 1406 1341 1556
rect 1346 1546 1349 1646
rect 1354 1623 1357 1696
rect 1362 1633 1365 1736
rect 1362 1553 1365 1626
rect 1346 1543 1365 1546
rect 1346 1533 1365 1536
rect 1346 1503 1349 1526
rect 1346 1423 1349 1466
rect 1362 1433 1365 1533
rect 1370 1503 1373 1743
rect 1378 1733 1381 1786
rect 1386 1733 1389 1833
rect 1394 1813 1397 1826
rect 1418 1813 1421 1953
rect 1426 1913 1429 1936
rect 1434 1903 1437 1946
rect 1394 1716 1397 1786
rect 1402 1776 1405 1796
rect 1410 1783 1413 1796
rect 1402 1773 1413 1776
rect 1386 1713 1397 1716
rect 1362 1423 1373 1426
rect 1378 1423 1381 1646
rect 1386 1433 1389 1713
rect 1394 1613 1397 1706
rect 1402 1663 1405 1716
rect 1410 1713 1413 1773
rect 1418 1726 1421 1806
rect 1426 1766 1429 1896
rect 1434 1773 1437 1816
rect 1442 1813 1445 1996
rect 1450 1803 1453 2016
rect 1450 1776 1453 1796
rect 1446 1773 1453 1776
rect 1426 1763 1437 1766
rect 1418 1723 1429 1726
rect 1402 1653 1421 1656
rect 1402 1606 1405 1653
rect 1394 1603 1405 1606
rect 1394 1503 1397 1603
rect 1354 1413 1381 1416
rect 1338 1403 1357 1406
rect 1330 1393 1341 1396
rect 1306 1263 1313 1266
rect 1310 1196 1313 1263
rect 1330 1236 1333 1326
rect 1338 1283 1341 1393
rect 1346 1293 1349 1326
rect 1354 1286 1357 1403
rect 1362 1326 1365 1346
rect 1362 1323 1373 1326
rect 1346 1283 1357 1286
rect 1338 1243 1341 1276
rect 1330 1233 1341 1236
rect 1306 1193 1313 1196
rect 1306 1006 1309 1193
rect 1314 1013 1317 1176
rect 1322 1106 1325 1216
rect 1330 1123 1333 1226
rect 1322 1103 1329 1106
rect 1326 1036 1329 1103
rect 1322 1033 1329 1036
rect 1306 1003 1317 1006
rect 1298 993 1309 996
rect 1266 923 1269 946
rect 1274 933 1301 936
rect 1258 903 1265 906
rect 1262 836 1265 903
rect 1262 833 1269 836
rect 1250 823 1261 826
rect 1202 733 1213 736
rect 1218 733 1221 746
rect 1234 733 1237 816
rect 1242 753 1245 806
rect 1202 656 1205 733
rect 1194 653 1205 656
rect 1194 543 1197 653
rect 1186 493 1189 526
rect 1194 513 1197 536
rect 1194 463 1197 506
rect 1178 413 1181 446
rect 1166 403 1177 406
rect 1162 343 1165 356
rect 1174 316 1177 403
rect 1186 323 1189 406
rect 1194 343 1197 416
rect 1202 333 1205 636
rect 1210 593 1213 606
rect 1218 576 1221 696
rect 1226 596 1229 726
rect 1242 703 1245 736
rect 1250 636 1253 816
rect 1258 753 1261 806
rect 1266 763 1269 833
rect 1274 743 1277 933
rect 1282 863 1285 926
rect 1306 923 1309 993
rect 1290 796 1293 826
rect 1306 816 1309 846
rect 1314 823 1317 1003
rect 1306 813 1317 816
rect 1298 803 1309 806
rect 1314 803 1317 813
rect 1290 793 1301 796
rect 1242 633 1253 636
rect 1234 613 1237 626
rect 1242 616 1245 633
rect 1242 613 1253 616
rect 1258 613 1261 666
rect 1282 656 1285 766
rect 1290 723 1293 746
rect 1282 653 1293 656
rect 1298 653 1301 793
rect 1322 786 1325 1033
rect 1338 1016 1341 1233
rect 1346 1216 1349 1283
rect 1354 1233 1357 1266
rect 1370 1226 1373 1323
rect 1386 1256 1389 1356
rect 1394 1343 1397 1436
rect 1362 1223 1373 1226
rect 1382 1253 1389 1256
rect 1402 1253 1405 1596
rect 1410 1333 1413 1626
rect 1418 1503 1421 1646
rect 1426 1596 1429 1723
rect 1434 1613 1437 1763
rect 1446 1686 1449 1773
rect 1446 1683 1453 1686
rect 1426 1593 1433 1596
rect 1430 1526 1433 1593
rect 1430 1523 1437 1526
rect 1346 1213 1353 1216
rect 1318 783 1325 786
rect 1330 1013 1341 1016
rect 1266 633 1285 636
rect 1226 593 1233 596
rect 1210 573 1221 576
rect 1210 443 1213 573
rect 1218 533 1221 566
rect 1230 536 1233 593
rect 1230 533 1237 536
rect 1242 533 1245 606
rect 1218 523 1229 526
rect 1234 496 1237 533
rect 1242 513 1245 526
rect 1234 493 1241 496
rect 1210 403 1213 426
rect 1218 413 1221 486
rect 1226 396 1229 476
rect 1238 426 1241 493
rect 1210 393 1229 396
rect 1234 423 1241 426
rect 1162 283 1165 316
rect 1174 313 1181 316
rect 1178 246 1181 313
rect 1194 263 1197 326
rect 1178 243 1189 246
rect 1170 213 1173 236
rect 1042 143 1045 156
rect 1042 113 1045 126
rect 1066 123 1069 136
rect 1114 113 1117 126
rect 1146 123 1149 173
rect 1162 163 1165 206
rect 1186 176 1189 243
rect 1210 223 1213 393
rect 1226 323 1229 336
rect 1218 303 1221 316
rect 1226 213 1229 266
rect 1234 233 1237 423
rect 1250 406 1253 613
rect 1266 556 1269 633
rect 1274 593 1277 626
rect 1282 603 1285 626
rect 1266 553 1277 556
rect 1258 453 1261 546
rect 1266 523 1269 546
rect 1274 536 1277 553
rect 1274 533 1285 536
rect 1290 526 1293 653
rect 1306 643 1309 736
rect 1318 716 1321 783
rect 1330 723 1333 1013
rect 1350 1006 1353 1213
rect 1362 1013 1365 1223
rect 1382 1206 1385 1253
rect 1378 1203 1385 1206
rect 1378 1146 1381 1203
rect 1378 1143 1389 1146
rect 1338 993 1341 1006
rect 1346 1003 1353 1006
rect 1338 933 1341 946
rect 1346 926 1349 1003
rect 1370 993 1373 1006
rect 1342 923 1349 926
rect 1342 836 1345 923
rect 1338 833 1345 836
rect 1338 783 1341 833
rect 1346 776 1349 816
rect 1354 813 1357 986
rect 1378 953 1381 1126
rect 1386 1123 1389 1143
rect 1362 913 1365 926
rect 1378 916 1381 946
rect 1374 913 1381 916
rect 1374 856 1377 913
rect 1362 813 1365 856
rect 1370 853 1377 856
rect 1338 773 1349 776
rect 1318 713 1325 716
rect 1314 636 1317 666
rect 1306 633 1317 636
rect 1322 636 1325 713
rect 1322 633 1333 636
rect 1306 613 1309 633
rect 1314 623 1325 626
rect 1282 523 1293 526
rect 1282 426 1285 523
rect 1298 506 1301 536
rect 1314 533 1317 623
rect 1330 606 1333 633
rect 1326 603 1333 606
rect 1326 526 1329 603
rect 1322 523 1329 526
rect 1298 503 1309 506
rect 1306 436 1309 503
rect 1306 433 1317 436
rect 1242 403 1253 406
rect 1258 423 1285 426
rect 1242 326 1245 403
rect 1258 383 1261 423
rect 1266 393 1269 416
rect 1282 413 1301 416
rect 1266 326 1269 346
rect 1242 323 1269 326
rect 1250 293 1253 306
rect 1266 223 1269 316
rect 1274 303 1277 326
rect 1282 296 1285 413
rect 1314 403 1317 433
rect 1322 396 1325 523
rect 1314 393 1325 396
rect 1298 323 1309 326
rect 1314 303 1317 393
rect 1330 313 1333 426
rect 1338 393 1341 773
rect 1362 753 1365 806
rect 1346 733 1357 736
rect 1346 716 1349 733
rect 1346 713 1353 716
rect 1350 626 1353 713
rect 1362 653 1365 736
rect 1346 623 1353 626
rect 1370 626 1373 853
rect 1378 803 1381 816
rect 1386 763 1389 1006
rect 1394 746 1397 1246
rect 1402 1113 1405 1186
rect 1410 1163 1413 1326
rect 1418 1293 1421 1496
rect 1426 1463 1429 1516
rect 1426 1333 1429 1446
rect 1418 1223 1421 1246
rect 1402 946 1405 1016
rect 1410 993 1413 1146
rect 1402 943 1413 946
rect 1402 823 1405 936
rect 1410 863 1413 943
rect 1378 743 1397 746
rect 1378 643 1381 743
rect 1386 713 1389 736
rect 1402 726 1405 816
rect 1410 733 1413 846
rect 1418 826 1421 1156
rect 1426 1113 1429 1326
rect 1434 1323 1437 1523
rect 1434 1223 1437 1296
rect 1426 1013 1429 1076
rect 1426 913 1429 926
rect 1434 843 1437 1136
rect 1442 1043 1445 1666
rect 1450 1593 1453 1683
rect 1450 1513 1453 1536
rect 1450 1363 1453 1456
rect 1458 1443 1461 2016
rect 1466 1983 1469 2026
rect 1474 1993 1477 2006
rect 1466 1923 1469 1976
rect 1474 1923 1477 1936
rect 1482 1916 1485 2126
rect 1490 2113 1493 2126
rect 1514 2103 1517 2136
rect 1490 2043 1517 2046
rect 1490 2003 1493 2043
rect 1498 2013 1501 2026
rect 1506 2003 1509 2036
rect 1514 2003 1517 2043
rect 1490 1923 1493 1966
rect 1474 1913 1485 1916
rect 1474 1846 1477 1913
rect 1466 1843 1477 1846
rect 1466 1716 1469 1843
rect 1482 1813 1485 1826
rect 1474 1783 1477 1806
rect 1490 1803 1493 1906
rect 1498 1763 1501 1926
rect 1474 1733 1501 1736
rect 1466 1713 1493 1716
rect 1466 1693 1469 1713
rect 1466 1613 1469 1626
rect 1474 1606 1477 1636
rect 1470 1603 1477 1606
rect 1470 1536 1473 1603
rect 1466 1533 1473 1536
rect 1466 1503 1469 1533
rect 1474 1476 1477 1516
rect 1466 1473 1477 1476
rect 1458 1396 1461 1426
rect 1466 1403 1469 1473
rect 1474 1443 1477 1473
rect 1474 1413 1477 1426
rect 1458 1393 1469 1396
rect 1466 1333 1469 1393
rect 1450 1223 1453 1266
rect 1458 1133 1461 1326
rect 1466 1283 1469 1316
rect 1474 1226 1477 1346
rect 1466 1223 1477 1226
rect 1466 1133 1469 1223
rect 1474 1203 1477 1216
rect 1482 1176 1485 1676
rect 1490 1183 1493 1706
rect 1498 1673 1501 1726
rect 1506 1663 1509 1946
rect 1514 1913 1517 1936
rect 1506 1613 1509 1646
rect 1514 1616 1517 1906
rect 1522 1696 1525 2173
rect 1538 2136 1541 2166
rect 1530 2133 1541 2136
rect 1530 1916 1533 2133
rect 1538 2123 1549 2126
rect 1538 1933 1541 1996
rect 1530 1913 1537 1916
rect 1546 1913 1549 2123
rect 1554 2103 1557 2413
rect 1562 2286 1565 2406
rect 1570 2373 1573 2406
rect 1586 2336 1589 2396
rect 1610 2376 1613 2416
rect 1626 2393 1629 2436
rect 1674 2403 1677 2416
rect 1610 2373 1629 2376
rect 1706 2373 1709 2416
rect 1582 2333 1589 2336
rect 1602 2333 1605 2346
rect 1570 2303 1573 2326
rect 1562 2283 1569 2286
rect 1566 2186 1569 2283
rect 1582 2266 1585 2333
rect 1594 2293 1597 2326
rect 1610 2276 1613 2336
rect 1626 2333 1629 2373
rect 1666 2333 1669 2346
rect 1650 2313 1653 2326
rect 1610 2273 1621 2276
rect 1582 2263 1589 2266
rect 1586 2243 1589 2263
rect 1578 2223 1597 2226
rect 1578 2213 1581 2223
rect 1594 2216 1597 2223
rect 1586 2203 1589 2216
rect 1594 2213 1605 2216
rect 1566 2183 1573 2186
rect 1570 2116 1573 2183
rect 1610 2156 1613 2226
rect 1618 2203 1621 2273
rect 1642 2203 1645 2216
rect 1610 2153 1621 2156
rect 1562 2113 1573 2116
rect 1594 2113 1597 2136
rect 1562 2063 1565 2113
rect 1570 2013 1573 2096
rect 1578 2023 1581 2036
rect 1586 1993 1589 2086
rect 1602 2036 1605 2136
rect 1610 2123 1613 2146
rect 1618 2123 1621 2153
rect 1610 2096 1613 2116
rect 1610 2093 1617 2096
rect 1594 2033 1605 2036
rect 1614 2026 1617 2093
rect 1610 2023 1617 2026
rect 1534 1846 1537 1913
rect 1530 1843 1537 1846
rect 1530 1803 1533 1843
rect 1538 1746 1541 1826
rect 1530 1743 1541 1746
rect 1530 1716 1533 1743
rect 1546 1723 1549 1856
rect 1554 1803 1557 1936
rect 1530 1713 1549 1716
rect 1554 1713 1557 1736
rect 1522 1693 1529 1696
rect 1526 1626 1529 1693
rect 1538 1643 1541 1706
rect 1526 1623 1533 1626
rect 1514 1613 1525 1616
rect 1498 1513 1501 1596
rect 1530 1556 1533 1623
rect 1522 1553 1533 1556
rect 1498 1403 1501 1466
rect 1506 1396 1509 1546
rect 1522 1533 1525 1553
rect 1530 1533 1533 1546
rect 1514 1493 1517 1526
rect 1538 1503 1541 1606
rect 1546 1496 1549 1713
rect 1554 1613 1557 1696
rect 1554 1513 1557 1576
rect 1562 1523 1565 1926
rect 1570 1903 1573 1986
rect 1586 1943 1589 1956
rect 1610 1933 1613 2023
rect 1578 1913 1581 1926
rect 1602 1873 1613 1876
rect 1570 1863 1597 1866
rect 1570 1823 1573 1863
rect 1570 1733 1573 1816
rect 1578 1813 1581 1856
rect 1586 1806 1589 1826
rect 1594 1813 1597 1863
rect 1578 1803 1589 1806
rect 1594 1803 1605 1806
rect 1570 1623 1573 1646
rect 1578 1613 1581 1803
rect 1586 1686 1589 1736
rect 1610 1733 1613 1873
rect 1618 1863 1621 1926
rect 1618 1803 1621 1856
rect 1618 1723 1621 1736
rect 1602 1703 1605 1716
rect 1626 1693 1629 2186
rect 1634 2093 1637 2126
rect 1634 1833 1637 1936
rect 1642 1886 1645 2166
rect 1658 2116 1661 2326
rect 1674 2296 1677 2326
rect 1682 2313 1685 2336
rect 1722 2333 1725 2416
rect 1730 2356 1733 2386
rect 1738 2366 1741 2406
rect 1754 2403 1757 2416
rect 1738 2363 1757 2366
rect 1730 2353 1741 2356
rect 1730 2316 1733 2346
rect 1722 2313 1733 2316
rect 1674 2293 1685 2296
rect 1666 2123 1669 2136
rect 1650 2113 1661 2116
rect 1650 2053 1653 2113
rect 1666 2106 1669 2116
rect 1658 2103 1669 2106
rect 1658 2073 1661 2103
rect 1674 2096 1677 2293
rect 1722 2246 1725 2313
rect 1738 2306 1741 2353
rect 1746 2323 1749 2346
rect 1754 2333 1757 2363
rect 1762 2353 1765 2396
rect 1786 2386 1789 2426
rect 1874 2423 1917 2426
rect 1786 2383 1793 2386
rect 1762 2343 1773 2346
rect 1778 2333 1781 2366
rect 1770 2323 1781 2326
rect 1738 2303 1749 2306
rect 1722 2243 1733 2246
rect 1682 2223 1701 2226
rect 1698 2206 1701 2223
rect 1706 2223 1725 2226
rect 1706 2213 1709 2223
rect 1698 2203 1709 2206
rect 1722 2203 1725 2223
rect 1682 2113 1685 2136
rect 1690 2113 1693 2146
rect 1658 1983 1661 2016
rect 1666 1993 1669 2096
rect 1674 2093 1681 2096
rect 1678 2016 1681 2093
rect 1674 2013 1681 2016
rect 1674 1996 1677 2013
rect 1674 1993 1685 1996
rect 1674 1973 1677 1993
rect 1650 1923 1661 1926
rect 1674 1923 1677 1956
rect 1690 1933 1693 2096
rect 1698 2083 1701 2203
rect 1706 2166 1709 2186
rect 1706 2163 1717 2166
rect 1714 2076 1717 2163
rect 1698 2073 1717 2076
rect 1642 1883 1653 1886
rect 1634 1773 1637 1816
rect 1642 1766 1645 1876
rect 1634 1763 1645 1766
rect 1586 1683 1597 1686
rect 1594 1606 1597 1683
rect 1570 1553 1573 1606
rect 1586 1603 1597 1606
rect 1586 1566 1589 1603
rect 1610 1573 1613 1606
rect 1586 1563 1605 1566
rect 1570 1496 1573 1536
rect 1538 1493 1549 1496
rect 1554 1493 1573 1496
rect 1514 1406 1517 1426
rect 1522 1413 1525 1446
rect 1530 1406 1533 1436
rect 1514 1403 1533 1406
rect 1502 1393 1509 1396
rect 1502 1246 1505 1393
rect 1530 1386 1533 1403
rect 1526 1383 1533 1386
rect 1514 1313 1517 1366
rect 1526 1296 1529 1383
rect 1538 1303 1541 1493
rect 1546 1323 1549 1416
rect 1554 1403 1557 1493
rect 1562 1363 1565 1466
rect 1570 1343 1573 1456
rect 1578 1443 1581 1546
rect 1554 1323 1565 1326
rect 1526 1293 1533 1296
rect 1498 1243 1505 1246
rect 1498 1203 1501 1243
rect 1474 1123 1477 1176
rect 1482 1173 1501 1176
rect 1482 1103 1485 1166
rect 1490 1096 1493 1126
rect 1450 1003 1453 1096
rect 1466 1093 1493 1096
rect 1466 1036 1469 1093
rect 1458 1033 1469 1036
rect 1442 903 1445 916
rect 1450 843 1453 936
rect 1418 823 1429 826
rect 1418 813 1437 816
rect 1418 756 1421 813
rect 1442 803 1445 836
rect 1426 763 1429 796
rect 1418 753 1429 756
rect 1394 693 1397 726
rect 1402 723 1413 726
rect 1410 713 1413 723
rect 1418 706 1421 736
rect 1402 656 1405 706
rect 1386 653 1405 656
rect 1370 623 1377 626
rect 1346 523 1349 623
rect 1354 563 1357 606
rect 1346 413 1349 436
rect 1346 356 1349 406
rect 1354 396 1357 546
rect 1362 483 1365 616
rect 1374 556 1377 623
rect 1386 613 1389 653
rect 1386 583 1389 596
rect 1370 553 1377 556
rect 1370 523 1373 553
rect 1378 493 1381 536
rect 1362 403 1365 456
rect 1370 416 1373 436
rect 1370 413 1377 416
rect 1354 393 1365 396
rect 1346 353 1357 356
rect 1338 333 1341 346
rect 1274 293 1285 296
rect 1210 193 1213 206
rect 1234 203 1237 216
rect 1258 203 1269 206
rect 1274 203 1277 293
rect 1338 216 1341 326
rect 1354 313 1357 353
rect 1306 213 1341 216
rect 1178 173 1189 176
rect 1178 133 1181 173
rect 1194 143 1197 156
rect 1186 133 1197 136
rect 1162 76 1165 126
rect 1186 76 1189 133
rect 1194 113 1197 126
rect 1218 123 1221 146
rect 1242 123 1245 166
rect 1258 143 1261 203
rect 1322 193 1325 206
rect 1362 196 1365 393
rect 1374 326 1377 413
rect 1386 403 1389 526
rect 1394 383 1397 646
rect 1402 496 1405 653
rect 1410 703 1421 706
rect 1410 613 1413 703
rect 1410 513 1413 546
rect 1402 493 1409 496
rect 1406 436 1409 493
rect 1418 443 1421 646
rect 1406 433 1421 436
rect 1402 413 1405 426
rect 1418 413 1421 433
rect 1386 333 1389 346
rect 1402 333 1405 406
rect 1426 396 1429 753
rect 1434 433 1437 736
rect 1442 623 1445 776
rect 1450 723 1453 816
rect 1442 473 1445 586
rect 1450 466 1453 616
rect 1458 483 1461 1033
rect 1482 1023 1485 1046
rect 1498 1033 1501 1173
rect 1506 1063 1509 1226
rect 1466 723 1469 1016
rect 1474 916 1477 926
rect 1482 923 1485 996
rect 1506 983 1509 1046
rect 1514 996 1517 1216
rect 1522 1153 1525 1226
rect 1522 1003 1525 1136
rect 1530 1073 1533 1293
rect 1514 993 1533 996
rect 1514 933 1517 946
rect 1522 933 1525 986
rect 1474 913 1501 916
rect 1514 913 1517 926
rect 1530 896 1533 993
rect 1522 893 1533 896
rect 1474 736 1477 866
rect 1482 813 1485 846
rect 1522 826 1525 893
rect 1538 833 1541 1186
rect 1546 1103 1549 1316
rect 1570 1306 1573 1336
rect 1566 1303 1573 1306
rect 1554 1213 1557 1226
rect 1566 1216 1569 1303
rect 1562 1213 1569 1216
rect 1578 1213 1581 1286
rect 1562 1133 1565 1213
rect 1586 1206 1589 1536
rect 1602 1533 1605 1563
rect 1610 1526 1613 1556
rect 1618 1533 1621 1666
rect 1594 1513 1597 1526
rect 1602 1523 1613 1526
rect 1594 1403 1597 1426
rect 1602 1396 1605 1523
rect 1610 1403 1613 1426
rect 1602 1393 1613 1396
rect 1594 1223 1597 1266
rect 1610 1263 1613 1393
rect 1618 1383 1621 1466
rect 1618 1283 1621 1326
rect 1626 1266 1629 1616
rect 1634 1543 1637 1763
rect 1642 1733 1645 1746
rect 1650 1726 1653 1883
rect 1642 1723 1653 1726
rect 1642 1553 1645 1723
rect 1650 1646 1653 1716
rect 1658 1653 1661 1923
rect 1666 1813 1669 1826
rect 1682 1813 1685 1916
rect 1698 1893 1701 2073
rect 1730 2036 1733 2243
rect 1746 2236 1749 2303
rect 1742 2233 1749 2236
rect 1742 2156 1745 2233
rect 1754 2173 1757 2216
rect 1742 2153 1749 2156
rect 1746 2046 1749 2153
rect 1762 2073 1765 2216
rect 1770 2203 1773 2323
rect 1790 2316 1793 2383
rect 1786 2313 1793 2316
rect 1778 2143 1781 2216
rect 1786 2126 1789 2313
rect 1802 2296 1805 2346
rect 1798 2293 1805 2296
rect 1798 2216 1801 2293
rect 1798 2213 1805 2216
rect 1794 2173 1797 2196
rect 1802 2133 1805 2213
rect 1770 2103 1773 2126
rect 1786 2123 1805 2126
rect 1778 2113 1789 2116
rect 1802 2083 1805 2123
rect 1810 2066 1813 2406
rect 1818 2346 1821 2416
rect 1826 2403 1837 2406
rect 1826 2373 1829 2396
rect 1818 2343 1829 2346
rect 1818 2243 1821 2336
rect 1826 2306 1829 2343
rect 1834 2326 1837 2403
rect 1842 2353 1845 2416
rect 1850 2383 1853 2416
rect 1858 2403 1861 2416
rect 1874 2403 1877 2423
rect 1890 2386 1893 2406
rect 1898 2403 1901 2416
rect 1906 2403 1909 2416
rect 1914 2403 1917 2423
rect 1930 2403 1973 2406
rect 1930 2393 1933 2403
rect 1946 2386 1949 2396
rect 1890 2383 1949 2386
rect 1858 2333 1901 2336
rect 1834 2323 1885 2326
rect 1850 2313 1877 2316
rect 1882 2313 1885 2323
rect 1826 2303 1837 2306
rect 1818 2143 1821 2206
rect 1826 2136 1829 2256
rect 1822 2133 1829 2136
rect 1834 2136 1837 2303
rect 1842 2213 1845 2246
rect 1874 2183 1877 2313
rect 1882 2223 1885 2236
rect 1874 2146 1877 2156
rect 1858 2143 1877 2146
rect 1834 2133 1853 2136
rect 1858 2133 1861 2143
rect 1822 2076 1825 2133
rect 1850 2126 1853 2133
rect 1806 2063 1813 2066
rect 1818 2073 1825 2076
rect 1706 2033 1733 2036
rect 1738 2043 1749 2046
rect 1706 2006 1709 2033
rect 1738 2026 1741 2043
rect 1762 2036 1765 2056
rect 1762 2033 1769 2036
rect 1714 2013 1717 2026
rect 1722 2023 1741 2026
rect 1722 2013 1725 2023
rect 1706 2003 1733 2006
rect 1666 1793 1669 1806
rect 1690 1776 1693 1856
rect 1698 1796 1701 1816
rect 1706 1813 1709 1866
rect 1714 1803 1717 1836
rect 1698 1793 1705 1796
rect 1682 1773 1693 1776
rect 1682 1756 1685 1773
rect 1678 1753 1685 1756
rect 1666 1683 1669 1726
rect 1678 1666 1681 1753
rect 1666 1646 1669 1666
rect 1678 1663 1685 1666
rect 1650 1643 1661 1646
rect 1666 1643 1673 1646
rect 1650 1613 1653 1626
rect 1658 1623 1661 1643
rect 1658 1603 1661 1616
rect 1670 1596 1673 1643
rect 1666 1593 1673 1596
rect 1666 1536 1669 1593
rect 1634 1533 1653 1536
rect 1662 1533 1669 1536
rect 1650 1493 1653 1516
rect 1622 1263 1629 1266
rect 1578 1203 1589 1206
rect 1554 1096 1557 1126
rect 1578 1113 1581 1203
rect 1546 1093 1557 1096
rect 1546 863 1549 1093
rect 1490 803 1493 826
rect 1522 823 1533 826
rect 1474 733 1485 736
rect 1466 616 1469 686
rect 1474 663 1477 726
rect 1482 696 1485 733
rect 1498 716 1501 796
rect 1522 793 1525 806
rect 1506 733 1509 746
rect 1522 726 1525 776
rect 1514 723 1525 726
rect 1498 713 1525 716
rect 1482 693 1493 696
rect 1490 636 1493 693
rect 1482 633 1493 636
rect 1466 613 1477 616
rect 1466 593 1469 606
rect 1474 583 1477 613
rect 1482 543 1485 633
rect 1490 603 1493 616
rect 1498 596 1501 606
rect 1490 593 1501 596
rect 1474 533 1485 536
rect 1498 533 1501 546
rect 1466 513 1469 526
rect 1474 523 1485 526
rect 1474 496 1477 523
rect 1470 493 1477 496
rect 1450 463 1457 466
rect 1422 393 1429 396
rect 1374 323 1381 326
rect 1378 246 1381 323
rect 1378 243 1389 246
rect 1386 213 1389 243
rect 1354 193 1389 196
rect 1394 193 1397 326
rect 1410 283 1413 326
rect 1422 226 1425 393
rect 1410 213 1413 226
rect 1422 223 1429 226
rect 1274 123 1277 186
rect 1282 123 1285 146
rect 1346 143 1349 166
rect 1322 123 1325 136
rect 1330 93 1333 126
rect 1386 123 1389 193
rect 1394 123 1397 146
rect 1410 133 1413 206
rect 1418 196 1421 206
rect 1426 203 1429 223
rect 1434 203 1437 416
rect 1442 413 1445 426
rect 1454 406 1457 463
rect 1470 436 1473 493
rect 1466 433 1473 436
rect 1454 403 1461 406
rect 1442 296 1445 326
rect 1458 323 1461 403
rect 1466 316 1469 433
rect 1474 413 1477 426
rect 1482 393 1485 496
rect 1450 303 1453 316
rect 1458 313 1469 316
rect 1474 333 1485 336
rect 1474 313 1477 333
rect 1442 293 1449 296
rect 1446 226 1449 293
rect 1446 223 1453 226
rect 1442 196 1445 206
rect 1418 193 1445 196
rect 1434 133 1437 146
rect 1442 93 1445 186
rect 1450 133 1453 223
rect 1458 133 1461 313
rect 1490 306 1493 526
rect 1498 403 1501 526
rect 1506 513 1509 626
rect 1506 423 1509 446
rect 1466 303 1493 306
rect 1466 283 1469 303
rect 1466 213 1469 226
rect 1474 213 1477 266
rect 1482 193 1485 206
rect 1490 203 1493 216
rect 1498 203 1501 326
rect 1506 243 1509 336
rect 1514 293 1517 706
rect 1522 593 1525 713
rect 1522 423 1525 526
rect 1522 393 1525 416
rect 1530 316 1533 823
rect 1538 693 1541 816
rect 1546 783 1549 826
rect 1554 773 1557 1086
rect 1562 1023 1565 1056
rect 1538 613 1541 686
rect 1546 613 1549 766
rect 1554 703 1557 736
rect 1562 686 1565 1016
rect 1570 906 1573 936
rect 1578 923 1581 976
rect 1570 903 1577 906
rect 1574 836 1577 903
rect 1570 833 1577 836
rect 1586 836 1589 1136
rect 1594 1123 1597 1206
rect 1602 1203 1605 1236
rect 1622 1196 1625 1263
rect 1606 1193 1625 1196
rect 1606 1136 1609 1193
rect 1602 1133 1609 1136
rect 1602 1053 1605 1133
rect 1610 1083 1613 1116
rect 1618 1093 1621 1136
rect 1610 1023 1613 1066
rect 1626 1026 1629 1126
rect 1634 1123 1637 1426
rect 1634 1083 1637 1106
rect 1626 1023 1633 1026
rect 1594 1003 1613 1006
rect 1594 933 1597 986
rect 1618 936 1621 1016
rect 1630 956 1633 1023
rect 1642 1003 1645 1486
rect 1662 1436 1665 1533
rect 1662 1433 1669 1436
rect 1650 1206 1653 1406
rect 1658 1346 1661 1416
rect 1666 1353 1669 1433
rect 1658 1343 1669 1346
rect 1658 1223 1661 1336
rect 1666 1213 1669 1343
rect 1674 1333 1677 1526
rect 1650 1203 1657 1206
rect 1654 986 1657 1203
rect 1666 1023 1669 1206
rect 1650 983 1657 986
rect 1650 963 1653 983
rect 1602 933 1621 936
rect 1626 953 1633 956
rect 1626 933 1629 953
rect 1586 833 1593 836
rect 1570 813 1573 833
rect 1570 793 1573 806
rect 1578 786 1581 816
rect 1570 783 1581 786
rect 1570 733 1573 783
rect 1590 756 1593 833
rect 1590 753 1597 756
rect 1570 703 1573 726
rect 1538 486 1541 606
rect 1554 533 1557 686
rect 1562 683 1569 686
rect 1566 536 1569 683
rect 1578 643 1581 726
rect 1586 683 1589 736
rect 1594 733 1597 753
rect 1594 713 1597 726
rect 1602 696 1605 933
rect 1598 693 1605 696
rect 1598 636 1601 693
rect 1578 633 1601 636
rect 1578 566 1581 633
rect 1586 613 1597 616
rect 1594 573 1597 606
rect 1602 603 1605 616
rect 1610 586 1613 926
rect 1618 723 1621 926
rect 1634 923 1645 926
rect 1626 913 1661 916
rect 1642 833 1645 856
rect 1626 783 1629 826
rect 1650 823 1653 836
rect 1634 806 1637 816
rect 1658 813 1661 913
rect 1666 806 1669 1006
rect 1634 803 1669 806
rect 1674 796 1677 1306
rect 1682 1233 1685 1663
rect 1690 1603 1693 1736
rect 1702 1706 1705 1793
rect 1702 1703 1709 1706
rect 1698 1646 1701 1696
rect 1706 1663 1709 1703
rect 1698 1643 1705 1646
rect 1702 1596 1705 1643
rect 1714 1626 1717 1796
rect 1722 1693 1725 1946
rect 1730 1676 1733 1976
rect 1738 1906 1741 2016
rect 1746 1983 1749 2006
rect 1754 1923 1757 2026
rect 1766 1916 1769 2033
rect 1794 2026 1797 2036
rect 1762 1913 1769 1916
rect 1778 2023 1797 2026
rect 1738 1903 1749 1906
rect 1746 1846 1749 1903
rect 1762 1853 1765 1913
rect 1722 1673 1733 1676
rect 1738 1843 1749 1846
rect 1722 1653 1725 1673
rect 1738 1666 1741 1843
rect 1746 1823 1765 1826
rect 1746 1803 1749 1823
rect 1754 1793 1757 1816
rect 1762 1813 1765 1823
rect 1730 1663 1741 1666
rect 1714 1623 1725 1626
rect 1698 1593 1705 1596
rect 1690 1316 1693 1516
rect 1698 1356 1701 1593
rect 1730 1583 1733 1663
rect 1738 1603 1741 1656
rect 1746 1613 1749 1716
rect 1770 1683 1773 1746
rect 1778 1723 1781 2023
rect 1806 2006 1809 2063
rect 1818 2013 1821 2073
rect 1826 2033 1829 2056
rect 1834 2016 1837 2126
rect 1842 2033 1845 2126
rect 1850 2123 1893 2126
rect 1898 2123 1901 2333
rect 1938 2323 1941 2356
rect 1946 2333 1949 2366
rect 1970 2333 1973 2403
rect 1978 2396 1981 2416
rect 2002 2413 2029 2416
rect 1978 2393 1989 2396
rect 1986 2336 1989 2393
rect 2018 2346 2021 2406
rect 1978 2333 1989 2336
rect 2002 2343 2021 2346
rect 1858 2023 1861 2066
rect 1830 2013 1837 2016
rect 1786 2003 1809 2006
rect 1786 1923 1789 2003
rect 1794 1933 1797 1956
rect 1794 1923 1805 1926
rect 1794 1813 1797 1856
rect 1802 1803 1805 1916
rect 1810 1813 1813 1996
rect 1818 1943 1821 1956
rect 1830 1936 1833 2013
rect 1818 1916 1821 1936
rect 1830 1933 1837 1936
rect 1818 1913 1825 1916
rect 1822 1836 1825 1913
rect 1818 1833 1825 1836
rect 1818 1816 1821 1833
rect 1818 1813 1829 1816
rect 1794 1733 1805 1736
rect 1794 1713 1797 1733
rect 1818 1723 1821 1806
rect 1818 1706 1821 1716
rect 1754 1643 1773 1646
rect 1746 1576 1749 1606
rect 1738 1573 1749 1576
rect 1706 1403 1709 1536
rect 1714 1523 1717 1546
rect 1738 1536 1741 1573
rect 1722 1533 1741 1536
rect 1746 1513 1749 1536
rect 1754 1506 1757 1616
rect 1714 1413 1717 1436
rect 1698 1353 1709 1356
rect 1698 1333 1701 1346
rect 1690 1313 1697 1316
rect 1694 1256 1697 1313
rect 1690 1253 1697 1256
rect 1690 1203 1693 1253
rect 1706 1236 1709 1353
rect 1722 1326 1725 1426
rect 1738 1376 1741 1506
rect 1746 1503 1757 1506
rect 1746 1423 1749 1503
rect 1754 1413 1757 1466
rect 1746 1383 1749 1406
rect 1762 1403 1765 1606
rect 1770 1546 1773 1643
rect 1778 1623 1781 1676
rect 1786 1613 1789 1706
rect 1802 1703 1821 1706
rect 1826 1703 1829 1736
rect 1802 1686 1805 1703
rect 1834 1696 1837 1933
rect 1842 1896 1845 1996
rect 1866 1953 1869 2026
rect 1874 2013 1877 2026
rect 1890 2016 1893 2046
rect 1898 2023 1901 2036
rect 1906 2023 1909 2136
rect 1914 2116 1917 2226
rect 1938 2223 1941 2236
rect 1946 2206 1949 2226
rect 1954 2213 1957 2326
rect 1978 2303 1981 2333
rect 2002 2326 2005 2343
rect 1998 2323 2005 2326
rect 1978 2233 1981 2246
rect 1970 2223 1981 2226
rect 1986 2223 1989 2316
rect 1998 2236 2001 2323
rect 1998 2233 2005 2236
rect 1978 2216 1981 2223
rect 1962 2213 1973 2216
rect 1978 2213 1997 2216
rect 1922 2203 1949 2206
rect 1970 2173 1973 2213
rect 2002 2186 2005 2233
rect 2010 2196 2013 2336
rect 2026 2333 2029 2413
rect 2034 2393 2037 2426
rect 2050 2413 2053 2453
rect 2042 2333 2045 2356
rect 2018 2283 2021 2326
rect 2034 2293 2037 2326
rect 2066 2316 2069 2436
rect 2090 2413 2093 2453
rect 2402 2453 2445 2456
rect 2146 2336 2149 2416
rect 2154 2413 2197 2416
rect 2154 2343 2157 2413
rect 2178 2383 2181 2396
rect 2202 2393 2205 2416
rect 2210 2396 2213 2406
rect 2218 2403 2221 2416
rect 2234 2403 2237 2446
rect 2242 2403 2245 2416
rect 2250 2396 2253 2406
rect 2266 2403 2269 2416
rect 2210 2393 2253 2396
rect 2266 2386 2269 2396
rect 2306 2393 2309 2446
rect 2266 2383 2277 2386
rect 2090 2333 2149 2336
rect 2058 2313 2069 2316
rect 2082 2316 2085 2326
rect 2082 2313 2093 2316
rect 2106 2313 2109 2326
rect 2058 2236 2061 2313
rect 2058 2233 2069 2236
rect 2034 2203 2037 2226
rect 2010 2193 2037 2196
rect 2002 2183 2029 2186
rect 1970 2163 2021 2166
rect 1930 2123 1933 2136
rect 1970 2133 1973 2163
rect 1914 2113 1957 2116
rect 1882 1936 1885 2016
rect 1890 2013 1901 2016
rect 1874 1933 1885 1936
rect 1850 1913 1853 1926
rect 1842 1893 1853 1896
rect 1850 1826 1853 1893
rect 1874 1836 1877 1933
rect 1890 1876 1893 1936
rect 1898 1913 1901 2013
rect 1906 1983 1909 2016
rect 1914 1943 1917 2086
rect 1930 2036 1933 2056
rect 1930 2033 1937 2036
rect 1922 1973 1925 2016
rect 1934 1976 1937 2033
rect 1930 1973 1937 1976
rect 1946 1973 1949 2006
rect 1962 2003 1965 2046
rect 1970 1986 1973 2076
rect 1978 2063 1981 2136
rect 1986 2123 1989 2156
rect 2002 2133 2005 2146
rect 2018 2143 2021 2163
rect 2026 2133 2029 2183
rect 2018 2046 2021 2126
rect 2034 2116 2037 2176
rect 2010 2043 2021 2046
rect 2030 2113 2037 2116
rect 2030 2046 2033 2113
rect 2030 2043 2037 2046
rect 1978 2003 1981 2026
rect 1930 1933 1933 1973
rect 1914 1886 1917 1926
rect 1954 1886 1957 1926
rect 1914 1883 1957 1886
rect 1962 1876 1965 1986
rect 1970 1983 1977 1986
rect 1890 1873 1941 1876
rect 1874 1833 1885 1836
rect 1798 1683 1805 1686
rect 1810 1693 1837 1696
rect 1842 1823 1853 1826
rect 1770 1543 1781 1546
rect 1770 1483 1773 1536
rect 1770 1413 1773 1426
rect 1778 1413 1781 1543
rect 1786 1526 1789 1576
rect 1798 1556 1801 1683
rect 1798 1553 1805 1556
rect 1802 1533 1805 1553
rect 1786 1523 1797 1526
rect 1770 1396 1773 1406
rect 1754 1393 1773 1396
rect 1738 1373 1749 1376
rect 1718 1323 1725 1326
rect 1718 1246 1721 1323
rect 1718 1243 1725 1246
rect 1698 1233 1709 1236
rect 1698 1196 1701 1233
rect 1682 1193 1701 1196
rect 1706 1193 1709 1226
rect 1714 1213 1717 1226
rect 1682 1113 1685 1193
rect 1682 1013 1685 1106
rect 1690 1076 1693 1126
rect 1698 1093 1701 1136
rect 1722 1126 1725 1243
rect 1730 1223 1733 1316
rect 1738 1253 1741 1356
rect 1746 1203 1749 1373
rect 1754 1323 1765 1326
rect 1770 1323 1773 1336
rect 1778 1313 1781 1406
rect 1786 1353 1789 1516
rect 1794 1336 1797 1523
rect 1802 1493 1805 1526
rect 1802 1413 1805 1456
rect 1810 1396 1813 1693
rect 1818 1603 1821 1616
rect 1826 1603 1829 1666
rect 1834 1613 1837 1686
rect 1842 1536 1845 1823
rect 1850 1753 1853 1806
rect 1866 1736 1869 1806
rect 1874 1793 1877 1816
rect 1882 1736 1885 1833
rect 1890 1813 1893 1826
rect 1854 1733 1869 1736
rect 1874 1733 1885 1736
rect 1854 1646 1857 1733
rect 1866 1653 1869 1726
rect 1850 1643 1857 1646
rect 1850 1623 1853 1643
rect 1874 1626 1877 1733
rect 1890 1713 1893 1756
rect 1898 1733 1901 1866
rect 1906 1783 1909 1816
rect 1914 1803 1917 1866
rect 1922 1746 1925 1846
rect 1930 1813 1933 1826
rect 1914 1743 1925 1746
rect 1898 1686 1901 1726
rect 1866 1623 1877 1626
rect 1882 1683 1901 1686
rect 1834 1533 1845 1536
rect 1818 1436 1821 1526
rect 1834 1466 1837 1533
rect 1834 1463 1845 1466
rect 1842 1443 1845 1463
rect 1818 1433 1837 1436
rect 1826 1403 1829 1426
rect 1810 1393 1829 1396
rect 1786 1333 1797 1336
rect 1786 1283 1789 1333
rect 1802 1313 1813 1316
rect 1818 1303 1821 1336
rect 1794 1256 1797 1266
rect 1718 1123 1725 1126
rect 1690 1073 1697 1076
rect 1694 1006 1697 1073
rect 1690 1003 1697 1006
rect 1682 893 1685 916
rect 1634 793 1677 796
rect 1682 793 1685 806
rect 1626 733 1629 746
rect 1634 733 1637 793
rect 1618 696 1621 716
rect 1618 693 1629 696
rect 1626 636 1629 693
rect 1606 583 1613 586
rect 1618 633 1629 636
rect 1578 563 1597 566
rect 1562 533 1569 536
rect 1546 523 1557 526
rect 1546 493 1549 523
rect 1554 486 1557 516
rect 1562 506 1565 533
rect 1570 513 1581 516
rect 1562 503 1581 506
rect 1586 503 1589 546
rect 1538 483 1557 486
rect 1538 413 1541 446
rect 1554 383 1557 406
rect 1562 393 1565 486
rect 1570 346 1573 446
rect 1546 323 1549 346
rect 1554 343 1573 346
rect 1530 313 1541 316
rect 1538 256 1541 313
rect 1554 263 1557 343
rect 1562 283 1565 316
rect 1538 253 1549 256
rect 1538 213 1541 226
rect 1546 203 1549 253
rect 1570 226 1573 336
rect 1578 253 1581 503
rect 1586 413 1589 426
rect 1586 323 1589 386
rect 1594 326 1597 563
rect 1606 526 1609 583
rect 1618 533 1621 633
rect 1606 523 1613 526
rect 1602 393 1605 406
rect 1610 383 1613 523
rect 1626 456 1629 526
rect 1642 513 1645 786
rect 1650 613 1653 736
rect 1658 723 1661 746
rect 1658 703 1661 716
rect 1666 603 1669 766
rect 1690 746 1693 1003
rect 1706 943 1709 1106
rect 1718 1026 1721 1123
rect 1730 1033 1733 1116
rect 1738 1093 1741 1136
rect 1762 1126 1765 1256
rect 1786 1253 1797 1256
rect 1778 1153 1781 1216
rect 1770 1133 1781 1136
rect 1746 1086 1749 1126
rect 1762 1123 1781 1126
rect 1778 1113 1781 1123
rect 1786 1106 1789 1253
rect 1794 1223 1821 1226
rect 1794 1173 1797 1216
rect 1802 1133 1805 1216
rect 1818 1206 1821 1223
rect 1826 1213 1829 1393
rect 1834 1376 1837 1433
rect 1850 1416 1853 1526
rect 1866 1436 1869 1623
rect 1882 1616 1885 1683
rect 1874 1613 1885 1616
rect 1890 1603 1893 1626
rect 1906 1613 1909 1636
rect 1914 1623 1917 1743
rect 1922 1733 1933 1736
rect 1938 1733 1941 1873
rect 1946 1873 1965 1876
rect 1946 1726 1949 1873
rect 1954 1813 1957 1826
rect 1962 1793 1965 1856
rect 1962 1743 1965 1756
rect 1974 1746 1977 1983
rect 1986 1973 1989 2016
rect 1994 2003 1997 2036
rect 1986 1803 1989 1826
rect 1994 1813 1997 1916
rect 2010 1863 2013 1926
rect 2002 1793 2005 1806
rect 2018 1803 2021 1946
rect 2034 1933 2037 2043
rect 2042 1996 2045 2206
rect 2050 2163 2053 2216
rect 2058 2193 2061 2216
rect 2066 2156 2069 2233
rect 2050 2153 2069 2156
rect 2050 2053 2053 2153
rect 2058 2003 2061 2126
rect 2066 2123 2069 2146
rect 2042 1993 2061 1996
rect 2066 1986 2069 2116
rect 2074 2033 2077 2266
rect 2082 2116 2085 2306
rect 2090 2296 2093 2313
rect 2090 2293 2101 2296
rect 2098 2226 2101 2293
rect 2090 2223 2101 2226
rect 2090 2206 2093 2223
rect 2114 2213 2117 2326
rect 2162 2303 2165 2336
rect 2178 2333 2205 2336
rect 2170 2256 2173 2326
rect 2146 2253 2173 2256
rect 2122 2206 2125 2216
rect 2090 2203 2125 2206
rect 2090 2133 2101 2136
rect 2114 2133 2117 2156
rect 2122 2146 2125 2203
rect 2122 2143 2133 2146
rect 2082 2113 2089 2116
rect 2086 2046 2089 2113
rect 2106 2103 2109 2126
rect 2122 2093 2125 2136
rect 2130 2056 2133 2143
rect 2082 2043 2089 2046
rect 2098 2053 2133 2056
rect 2074 1993 2077 2016
rect 2082 2006 2085 2043
rect 2090 2013 2093 2026
rect 2082 2003 2093 2006
rect 2066 1983 2077 1986
rect 2066 1936 2069 1946
rect 2058 1933 2069 1936
rect 2026 1813 2029 1876
rect 2034 1843 2037 1926
rect 2058 1916 2061 1933
rect 2074 1923 2077 1983
rect 2082 1933 2085 1956
rect 2090 1926 2093 2003
rect 2098 1963 2101 2053
rect 2138 2046 2141 2236
rect 2146 2196 2149 2253
rect 2178 2246 2181 2326
rect 2202 2323 2205 2333
rect 2202 2303 2205 2316
rect 2154 2243 2181 2246
rect 2154 2213 2157 2243
rect 2162 2213 2165 2226
rect 2178 2223 2181 2236
rect 2194 2233 2197 2246
rect 2146 2193 2157 2196
rect 2154 2126 2157 2193
rect 2150 2123 2157 2126
rect 2178 2123 2181 2136
rect 2186 2126 2189 2226
rect 2218 2156 2221 2366
rect 2242 2333 2245 2346
rect 2250 2333 2253 2366
rect 2274 2333 2277 2383
rect 2314 2346 2317 2416
rect 2330 2413 2349 2416
rect 2330 2403 2333 2413
rect 2282 2333 2285 2346
rect 2306 2343 2317 2346
rect 2258 2306 2261 2326
rect 2250 2303 2261 2306
rect 2250 2236 2253 2303
rect 2250 2233 2261 2236
rect 2226 2193 2229 2226
rect 2234 2213 2245 2216
rect 2258 2196 2261 2233
rect 2274 2226 2277 2316
rect 2306 2246 2309 2343
rect 2306 2243 2317 2246
rect 2266 2223 2277 2226
rect 2282 2206 2285 2216
rect 2306 2213 2309 2226
rect 2250 2193 2261 2196
rect 2266 2203 2285 2206
rect 2266 2193 2269 2203
rect 2210 2153 2221 2156
rect 2186 2123 2197 2126
rect 2150 2066 2153 2123
rect 2194 2113 2197 2123
rect 2122 2043 2141 2046
rect 2146 2063 2153 2066
rect 2146 2043 2149 2063
rect 2098 1933 2101 1946
rect 2082 1923 2093 1926
rect 2042 1913 2061 1916
rect 2042 1803 2045 1913
rect 1970 1743 1977 1746
rect 1930 1723 1949 1726
rect 1874 1543 1877 1576
rect 1882 1516 1885 1566
rect 1898 1533 1901 1576
rect 1878 1513 1885 1516
rect 1878 1456 1881 1513
rect 1878 1453 1885 1456
rect 1866 1433 1877 1436
rect 1850 1413 1869 1416
rect 1842 1393 1845 1406
rect 1850 1386 1853 1406
rect 1850 1383 1857 1386
rect 1834 1373 1845 1376
rect 1834 1246 1837 1326
rect 1842 1323 1845 1373
rect 1854 1316 1857 1383
rect 1850 1313 1857 1316
rect 1850 1263 1853 1313
rect 1866 1296 1869 1413
rect 1862 1293 1869 1296
rect 1834 1243 1845 1246
rect 1814 1203 1821 1206
rect 1814 1146 1817 1203
rect 1814 1143 1821 1146
rect 1818 1123 1821 1143
rect 1826 1133 1829 1206
rect 1842 1156 1845 1243
rect 1862 1196 1865 1293
rect 1874 1233 1877 1433
rect 1882 1353 1885 1453
rect 1890 1443 1893 1516
rect 1898 1496 1901 1526
rect 1906 1503 1909 1606
rect 1914 1533 1917 1616
rect 1922 1533 1925 1596
rect 1930 1563 1933 1723
rect 1946 1696 1949 1716
rect 1942 1693 1949 1696
rect 1914 1496 1917 1526
rect 1942 1516 1945 1693
rect 1954 1523 1957 1666
rect 1962 1603 1965 1626
rect 1970 1613 1973 1743
rect 1978 1696 1981 1726
rect 1986 1703 1989 1746
rect 1994 1713 1997 1726
rect 1978 1693 2001 1696
rect 1942 1513 1949 1516
rect 1962 1513 1965 1586
rect 1970 1553 1973 1606
rect 1898 1493 1917 1496
rect 1898 1453 1933 1456
rect 1890 1403 1893 1426
rect 1898 1423 1901 1453
rect 1906 1413 1909 1446
rect 1930 1413 1933 1453
rect 1898 1373 1901 1406
rect 1890 1333 1893 1346
rect 1898 1326 1901 1336
rect 1890 1323 1901 1326
rect 1906 1323 1909 1406
rect 1914 1323 1925 1326
rect 1890 1313 1893 1323
rect 1914 1316 1917 1323
rect 1898 1313 1917 1316
rect 1862 1193 1869 1196
rect 1834 1153 1845 1156
rect 1738 1083 1749 1086
rect 1778 1103 1789 1106
rect 1714 1023 1721 1026
rect 1714 1006 1717 1023
rect 1722 1013 1733 1016
rect 1714 1003 1721 1006
rect 1718 916 1721 1003
rect 1730 983 1733 1006
rect 1718 913 1725 916
rect 1698 853 1701 906
rect 1682 743 1693 746
rect 1698 746 1701 786
rect 1706 763 1709 816
rect 1698 743 1705 746
rect 1682 716 1685 743
rect 1678 713 1685 716
rect 1678 596 1681 713
rect 1674 593 1681 596
rect 1650 513 1653 536
rect 1658 533 1661 546
rect 1674 536 1677 593
rect 1682 543 1685 566
rect 1666 533 1685 536
rect 1626 453 1661 456
rect 1634 436 1637 446
rect 1634 433 1653 436
rect 1618 403 1621 416
rect 1634 413 1637 433
rect 1626 326 1629 406
rect 1642 403 1645 426
rect 1650 413 1653 433
rect 1650 356 1653 406
rect 1658 396 1661 453
rect 1666 413 1669 533
rect 1658 393 1665 396
rect 1642 353 1653 356
rect 1594 323 1613 326
rect 1626 323 1637 326
rect 1642 323 1645 353
rect 1662 346 1665 393
rect 1674 386 1677 526
rect 1682 513 1685 533
rect 1690 503 1693 736
rect 1702 646 1705 743
rect 1698 643 1705 646
rect 1698 436 1701 643
rect 1714 616 1717 896
rect 1722 723 1725 913
rect 1730 803 1733 966
rect 1730 723 1733 766
rect 1706 613 1717 616
rect 1706 603 1709 613
rect 1714 563 1717 606
rect 1722 603 1725 636
rect 1730 576 1733 716
rect 1738 703 1741 1083
rect 1778 1026 1781 1103
rect 1826 1063 1829 1126
rect 1834 1096 1837 1153
rect 1858 1136 1861 1176
rect 1842 1113 1845 1136
rect 1850 1133 1861 1136
rect 1834 1093 1845 1096
rect 1842 1036 1845 1093
rect 1774 1023 1781 1026
rect 1762 1003 1765 1016
rect 1746 913 1749 976
rect 1774 966 1777 1023
rect 1826 1016 1829 1036
rect 1786 983 1789 1016
rect 1794 1013 1805 1016
rect 1810 1013 1829 1016
rect 1834 1033 1845 1036
rect 1754 913 1757 946
rect 1746 646 1749 866
rect 1754 803 1757 906
rect 1762 853 1765 966
rect 1774 963 1781 966
rect 1754 723 1757 796
rect 1762 733 1765 826
rect 1770 726 1773 946
rect 1762 723 1773 726
rect 1746 643 1753 646
rect 1738 613 1741 636
rect 1722 573 1733 576
rect 1722 526 1725 573
rect 1706 493 1709 526
rect 1718 523 1725 526
rect 1718 466 1721 523
rect 1718 463 1725 466
rect 1698 433 1709 436
rect 1682 393 1685 416
rect 1698 403 1701 426
rect 1674 383 1685 386
rect 1658 343 1665 346
rect 1682 346 1685 383
rect 1682 343 1693 346
rect 1594 303 1597 323
rect 1570 223 1597 226
rect 1586 213 1597 216
rect 1586 206 1589 213
rect 1498 193 1509 196
rect 1498 143 1509 146
rect 1562 133 1565 206
rect 1570 203 1589 206
rect 1594 193 1597 206
rect 1602 203 1605 316
rect 1610 303 1613 323
rect 1618 303 1621 316
rect 1634 253 1637 323
rect 1658 213 1661 343
rect 1690 323 1693 336
rect 1690 213 1693 256
rect 1706 213 1709 433
rect 1714 413 1717 446
rect 1722 233 1725 463
rect 1730 386 1733 516
rect 1738 513 1741 606
rect 1750 546 1753 643
rect 1762 596 1765 723
rect 1770 613 1773 656
rect 1778 603 1781 963
rect 1786 933 1789 946
rect 1794 943 1797 1013
rect 1786 813 1789 916
rect 1802 893 1805 1006
rect 1810 876 1813 1013
rect 1818 983 1821 1006
rect 1826 946 1829 1006
rect 1802 873 1813 876
rect 1818 943 1829 946
rect 1786 783 1789 806
rect 1802 796 1805 873
rect 1818 863 1821 943
rect 1826 833 1829 936
rect 1818 813 1829 816
rect 1802 793 1813 796
rect 1802 733 1805 776
rect 1810 736 1813 793
rect 1818 763 1821 796
rect 1810 733 1821 736
rect 1826 733 1829 813
rect 1794 723 1805 726
rect 1810 713 1813 726
rect 1818 716 1821 733
rect 1818 713 1825 716
rect 1786 616 1789 686
rect 1802 623 1805 656
rect 1786 613 1805 616
rect 1762 593 1789 596
rect 1746 543 1753 546
rect 1738 423 1741 466
rect 1738 393 1741 416
rect 1746 406 1749 543
rect 1770 526 1773 536
rect 1778 526 1781 536
rect 1754 523 1781 526
rect 1754 413 1757 523
rect 1786 516 1789 593
rect 1762 433 1765 506
rect 1746 403 1757 406
rect 1730 383 1749 386
rect 1738 293 1741 326
rect 1658 166 1661 206
rect 1666 193 1677 196
rect 1658 163 1717 166
rect 1594 143 1597 156
rect 1506 123 1525 126
rect 1618 86 1621 126
rect 1634 103 1637 136
rect 1658 86 1661 126
rect 1714 123 1717 163
rect 1722 133 1725 206
rect 1730 196 1733 206
rect 1746 203 1749 383
rect 1754 356 1757 403
rect 1770 363 1773 516
rect 1778 513 1789 516
rect 1778 403 1781 513
rect 1794 446 1797 566
rect 1810 496 1813 706
rect 1822 616 1825 713
rect 1822 613 1829 616
rect 1818 516 1821 606
rect 1826 573 1829 613
rect 1834 603 1837 1033
rect 1866 1016 1869 1193
rect 1874 1153 1877 1226
rect 1850 1013 1869 1016
rect 1842 933 1845 976
rect 1842 893 1845 926
rect 1850 826 1853 1013
rect 1882 1006 1885 1306
rect 1890 1113 1893 1236
rect 1898 1213 1909 1216
rect 1914 1213 1917 1236
rect 1898 1146 1901 1196
rect 1898 1143 1917 1146
rect 1890 1013 1893 1026
rect 1898 1006 1901 1143
rect 1906 1116 1909 1136
rect 1906 1113 1913 1116
rect 1866 1003 1885 1006
rect 1890 1003 1901 1006
rect 1858 893 1861 956
rect 1866 913 1869 1003
rect 1890 996 1893 1003
rect 1874 993 1893 996
rect 1898 983 1901 1003
rect 1910 966 1913 1113
rect 1906 963 1913 966
rect 1906 946 1909 963
rect 1922 956 1925 1266
rect 1930 1123 1933 1366
rect 1938 1343 1941 1436
rect 1938 1203 1941 1316
rect 1946 1233 1949 1513
rect 1954 1423 1957 1436
rect 1962 1423 1965 1506
rect 1970 1493 1973 1516
rect 1954 1343 1957 1416
rect 1954 1226 1957 1336
rect 1962 1303 1965 1376
rect 1970 1313 1973 1416
rect 1978 1303 1981 1646
rect 1986 1603 1989 1686
rect 1998 1626 2001 1693
rect 1998 1623 2005 1626
rect 2002 1603 2005 1623
rect 2010 1613 2013 1706
rect 2018 1703 2021 1766
rect 2050 1726 2053 1846
rect 2066 1813 2069 1876
rect 2074 1836 2077 1916
rect 2082 1853 2085 1923
rect 2074 1833 2081 1836
rect 2066 1793 2069 1806
rect 2078 1786 2081 1833
rect 2090 1803 2093 1916
rect 2098 1903 2101 1926
rect 2098 1813 2101 1846
rect 2106 1816 2109 2026
rect 2114 2003 2117 2026
rect 2106 1813 2117 1816
rect 2098 1803 2109 1806
rect 2074 1783 2081 1786
rect 2026 1683 2029 1726
rect 2038 1723 2053 1726
rect 2038 1676 2041 1723
rect 2034 1673 2041 1676
rect 2034 1626 2037 1673
rect 2018 1623 2037 1626
rect 2050 1623 2053 1716
rect 1986 1523 1989 1566
rect 1994 1456 1997 1526
rect 2002 1513 2005 1536
rect 1994 1453 2001 1456
rect 2010 1453 2013 1606
rect 1986 1423 1989 1446
rect 1986 1393 1989 1406
rect 1998 1386 2001 1453
rect 2018 1446 2021 1623
rect 2026 1613 2053 1616
rect 2026 1493 2029 1613
rect 2058 1606 2061 1746
rect 2074 1726 2077 1783
rect 2066 1723 2077 1726
rect 2066 1696 2069 1723
rect 2082 1716 2085 1736
rect 2074 1713 2085 1716
rect 2066 1693 2073 1696
rect 2070 1626 2073 1693
rect 2070 1623 2077 1626
rect 2034 1596 2037 1606
rect 2042 1603 2061 1606
rect 2066 1596 2069 1616
rect 2034 1593 2069 1596
rect 2074 1596 2077 1623
rect 2082 1613 2085 1696
rect 2074 1593 2085 1596
rect 1994 1383 2001 1386
rect 2010 1443 2021 1446
rect 1986 1293 1989 1336
rect 1994 1263 1997 1383
rect 1946 1203 1949 1226
rect 1954 1223 1973 1226
rect 1962 1173 1965 1216
rect 1970 1193 1973 1223
rect 1986 1213 1989 1256
rect 2002 1246 2005 1356
rect 2010 1293 2013 1443
rect 2018 1413 2021 1436
rect 2026 1403 2029 1416
rect 2034 1386 2037 1586
rect 2058 1583 2077 1586
rect 2058 1536 2061 1583
rect 2082 1576 2085 1593
rect 2090 1583 2093 1746
rect 2098 1683 2101 1796
rect 2114 1786 2117 1813
rect 2110 1783 2117 1786
rect 2122 1783 2125 2043
rect 2130 2016 2133 2036
rect 2138 2033 2157 2036
rect 2130 2013 2157 2016
rect 2130 1956 2133 1976
rect 2162 1956 2165 2106
rect 2210 2056 2213 2153
rect 2210 2053 2221 2056
rect 2170 2023 2173 2036
rect 2194 2033 2213 2036
rect 2130 1953 2141 1956
rect 2138 1836 2141 1953
rect 2154 1953 2165 1956
rect 2154 1866 2157 1953
rect 2170 1913 2173 1946
rect 2178 1906 2181 2026
rect 2202 1936 2205 2026
rect 2210 2013 2213 2033
rect 2218 1983 2221 2053
rect 2226 1996 2229 2146
rect 2250 2133 2253 2193
rect 2314 2186 2317 2243
rect 2322 2196 2325 2336
rect 2330 2333 2349 2336
rect 2354 2333 2357 2406
rect 2370 2346 2373 2406
rect 2386 2393 2389 2426
rect 2402 2413 2405 2453
rect 2418 2403 2421 2436
rect 2442 2413 2445 2453
rect 2498 2396 2501 2416
rect 2490 2393 2501 2396
rect 2370 2343 2381 2346
rect 2330 2283 2333 2333
rect 2338 2286 2341 2326
rect 2346 2323 2349 2333
rect 2362 2293 2365 2326
rect 2370 2286 2373 2336
rect 2338 2283 2373 2286
rect 2338 2203 2341 2226
rect 2322 2193 2341 2196
rect 2314 2183 2325 2186
rect 2290 2173 2317 2176
rect 2242 2023 2245 2126
rect 2226 1993 2245 1996
rect 2194 1933 2205 1936
rect 2250 1936 2253 2126
rect 2258 2123 2261 2146
rect 2290 2133 2293 2173
rect 2314 2143 2317 2173
rect 2298 2106 2301 2126
rect 2294 2103 2301 2106
rect 2258 2006 2261 2056
rect 2266 2013 2269 2046
rect 2294 2036 2297 2103
rect 2258 2003 2269 2006
rect 2250 1933 2261 1936
rect 2186 1913 2189 1926
rect 2178 1903 2197 1906
rect 2154 1863 2173 1866
rect 2130 1833 2141 1836
rect 2110 1716 2113 1783
rect 2130 1736 2133 1833
rect 2138 1793 2141 1816
rect 2154 1803 2157 1816
rect 2162 1813 2165 1856
rect 2170 1806 2173 1863
rect 2162 1803 2173 1806
rect 2122 1733 2133 1736
rect 2146 1733 2149 1756
rect 2110 1713 2117 1716
rect 2106 1653 2109 1696
rect 2042 1533 2061 1536
rect 2066 1533 2069 1576
rect 2074 1573 2085 1576
rect 2042 1516 2045 1533
rect 2050 1523 2061 1526
rect 2042 1513 2053 1516
rect 2066 1513 2069 1526
rect 2042 1393 2045 1416
rect 2018 1383 2037 1386
rect 2018 1283 2021 1383
rect 2026 1333 2029 1376
rect 2050 1356 2053 1513
rect 2074 1506 2077 1573
rect 2066 1503 2077 1506
rect 2058 1413 2061 1446
rect 2058 1383 2061 1406
rect 2034 1333 2037 1356
rect 2042 1353 2053 1356
rect 1994 1243 2005 1246
rect 1994 1206 1997 1243
rect 1978 1203 1997 1206
rect 1954 1123 1965 1126
rect 1938 1003 1941 1056
rect 1954 1003 1957 1016
rect 1962 1013 1965 1076
rect 1970 996 1973 1136
rect 1978 1093 1981 1203
rect 1986 1123 1989 1186
rect 1978 1023 1981 1086
rect 1986 1013 1989 1116
rect 1962 983 1965 996
rect 1970 993 1981 996
rect 1922 953 1949 956
rect 1898 943 1909 946
rect 1874 923 1877 936
rect 1882 846 1885 926
rect 1890 923 1893 936
rect 1898 883 1901 943
rect 1866 843 1885 846
rect 1850 823 1857 826
rect 1842 773 1845 816
rect 1854 766 1857 823
rect 1866 796 1869 843
rect 1874 806 1877 836
rect 1906 826 1909 936
rect 1914 933 1925 936
rect 1914 893 1917 926
rect 1930 923 1933 936
rect 1938 933 1941 946
rect 1890 823 1909 826
rect 1874 803 1885 806
rect 1866 793 1885 796
rect 1854 763 1877 766
rect 1842 613 1845 706
rect 1826 523 1829 566
rect 1850 526 1853 736
rect 1874 703 1877 763
rect 1882 716 1885 793
rect 1890 763 1893 823
rect 1898 793 1901 806
rect 1906 786 1909 816
rect 1898 783 1909 786
rect 1898 723 1901 783
rect 1882 713 1897 716
rect 1858 616 1861 636
rect 1858 613 1869 616
rect 1874 613 1877 676
rect 1866 606 1869 613
rect 1858 533 1861 606
rect 1866 603 1877 606
rect 1882 603 1885 686
rect 1850 523 1861 526
rect 1818 513 1837 516
rect 1834 503 1837 513
rect 1842 496 1845 516
rect 1810 493 1845 496
rect 1850 493 1853 516
rect 1786 443 1797 446
rect 1786 403 1789 443
rect 1794 423 1845 426
rect 1818 413 1829 416
rect 1754 353 1773 356
rect 1754 203 1757 326
rect 1762 246 1765 336
rect 1770 273 1773 353
rect 1794 333 1797 346
rect 1810 333 1813 366
rect 1818 343 1821 406
rect 1826 263 1829 413
rect 1834 393 1837 406
rect 1842 403 1845 423
rect 1842 323 1845 356
rect 1858 316 1861 523
rect 1866 506 1869 576
rect 1874 523 1877 603
rect 1894 546 1897 713
rect 1914 686 1917 856
rect 1922 823 1925 886
rect 1906 683 1917 686
rect 1894 543 1901 546
rect 1882 523 1885 536
rect 1898 526 1901 543
rect 1906 533 1909 683
rect 1922 653 1925 796
rect 1922 623 1925 636
rect 1930 613 1933 836
rect 1938 593 1941 886
rect 1946 836 1949 953
rect 1954 843 1957 936
rect 1946 833 1957 836
rect 1946 763 1949 826
rect 1954 813 1957 833
rect 1946 723 1957 726
rect 1954 693 1957 723
rect 1946 576 1949 666
rect 1942 573 1949 576
rect 1898 523 1909 526
rect 1890 513 1901 516
rect 1866 503 1877 506
rect 1874 436 1877 503
rect 1866 433 1877 436
rect 1866 413 1869 433
rect 1890 413 1893 426
rect 1898 393 1901 406
rect 1906 376 1909 523
rect 1914 486 1917 526
rect 1922 503 1925 566
rect 1930 513 1933 526
rect 1914 483 1925 486
rect 1922 426 1925 483
rect 1942 456 1945 573
rect 1942 453 1949 456
rect 1946 433 1949 453
rect 1922 423 1949 426
rect 1914 396 1917 406
rect 1930 403 1933 416
rect 1914 393 1925 396
rect 1938 393 1941 406
rect 1842 313 1861 316
rect 1762 243 1781 246
rect 1762 196 1765 226
rect 1730 193 1765 196
rect 1770 143 1773 156
rect 1778 143 1781 243
rect 1794 243 1829 246
rect 1794 213 1797 243
rect 1802 193 1805 216
rect 1818 213 1821 236
rect 1770 126 1773 136
rect 1810 133 1813 206
rect 1826 203 1829 243
rect 1746 123 1773 126
rect 1794 113 1797 126
rect 1842 103 1845 313
rect 1866 193 1869 336
rect 1874 333 1877 376
rect 1882 373 1909 376
rect 1874 313 1877 326
rect 1882 303 1885 373
rect 1890 323 1893 366
rect 1898 286 1901 346
rect 1906 323 1909 336
rect 1890 283 1901 286
rect 1890 236 1893 283
rect 1890 233 1901 236
rect 1898 213 1901 233
rect 1906 213 1909 306
rect 1914 283 1917 386
rect 1922 343 1925 393
rect 1946 356 1949 423
rect 1954 363 1957 616
rect 1962 513 1965 976
rect 1978 926 1981 993
rect 1994 933 1997 1196
rect 1970 923 1981 926
rect 1994 906 1997 926
rect 1990 903 1997 906
rect 1970 803 1973 826
rect 1978 813 1981 836
rect 1990 826 1993 903
rect 1990 823 1997 826
rect 2002 823 2005 1236
rect 2010 1176 2013 1276
rect 2018 1183 2021 1206
rect 2010 1173 2021 1176
rect 2010 1123 2013 1156
rect 2018 1143 2021 1173
rect 2026 1136 2029 1326
rect 2042 1233 2045 1353
rect 2058 1333 2061 1356
rect 2066 1306 2069 1503
rect 2082 1496 2085 1546
rect 2098 1536 2101 1606
rect 2106 1566 2109 1606
rect 2114 1576 2117 1713
rect 2122 1663 2125 1733
rect 2130 1723 2141 1726
rect 2154 1723 2157 1736
rect 2162 1716 2165 1803
rect 2178 1763 2181 1826
rect 2186 1803 2189 1826
rect 2194 1746 2197 1903
rect 2250 1843 2253 1926
rect 2266 1923 2269 2003
rect 2274 1933 2277 2006
rect 2282 2003 2285 2036
rect 2294 2033 2301 2036
rect 2290 1933 2293 2016
rect 2298 1996 2301 2033
rect 2306 2013 2309 2136
rect 2322 2126 2325 2183
rect 2362 2166 2365 2206
rect 2354 2163 2365 2166
rect 2370 2163 2373 2216
rect 2318 2123 2325 2126
rect 2318 2046 2321 2123
rect 2318 2043 2325 2046
rect 2314 2013 2317 2026
rect 2298 1993 2309 1996
rect 2306 1926 2309 1993
rect 2282 1916 2285 1926
rect 2258 1913 2285 1916
rect 2298 1923 2309 1926
rect 2322 1923 2325 2043
rect 2202 1823 2237 1826
rect 2210 1813 2213 1823
rect 2186 1743 2197 1746
rect 2122 1623 2125 1656
rect 2138 1603 2141 1686
rect 2146 1623 2149 1716
rect 2158 1713 2165 1716
rect 2158 1656 2161 1713
rect 2154 1653 2161 1656
rect 2114 1573 2133 1576
rect 2130 1566 2133 1573
rect 2106 1563 2117 1566
rect 2130 1563 2141 1566
rect 2074 1493 2085 1496
rect 2090 1533 2101 1536
rect 2074 1333 2077 1493
rect 2090 1486 2093 1533
rect 2098 1493 2101 1526
rect 2114 1523 2117 1563
rect 2122 1533 2125 1556
rect 2082 1483 2093 1486
rect 2082 1336 2085 1483
rect 2090 1413 2093 1446
rect 2090 1343 2093 1356
rect 2082 1333 2093 1336
rect 2066 1303 2073 1306
rect 2050 1223 2053 1246
rect 2034 1213 2045 1216
rect 2018 1133 2029 1136
rect 2042 1136 2045 1213
rect 2042 1133 2053 1136
rect 2010 996 2013 1086
rect 2018 1003 2021 1133
rect 2026 1113 2029 1126
rect 2050 1123 2053 1133
rect 2058 1106 2061 1296
rect 2070 1216 2073 1303
rect 2070 1213 2077 1216
rect 2066 1183 2069 1206
rect 2010 993 2021 996
rect 2010 853 2013 986
rect 2018 846 2021 993
rect 2010 843 2021 846
rect 1994 806 1997 823
rect 1978 796 1981 806
rect 1994 803 2005 806
rect 1994 796 1997 803
rect 1978 793 1997 796
rect 1970 673 1973 746
rect 1978 723 1981 786
rect 1986 716 1989 766
rect 1994 743 1997 756
rect 2010 743 2013 843
rect 2018 783 2021 836
rect 1978 713 1989 716
rect 1970 603 1973 656
rect 1970 426 1973 526
rect 1978 433 1981 713
rect 2010 706 2013 736
rect 2002 703 2013 706
rect 1986 616 1989 676
rect 2002 646 2005 703
rect 2018 666 2021 726
rect 2026 676 2029 1106
rect 2050 1103 2061 1106
rect 2034 803 2037 1096
rect 2050 1046 2053 1103
rect 2050 1043 2061 1046
rect 2058 1026 2061 1043
rect 2050 1023 2061 1026
rect 2050 1013 2053 1023
rect 2042 983 2045 1006
rect 2050 933 2053 996
rect 2042 893 2045 926
rect 2042 813 2045 876
rect 2058 833 2061 1023
rect 2066 993 2069 1146
rect 2074 1023 2077 1213
rect 2074 973 2077 1006
rect 2066 953 2077 956
rect 2034 683 2037 736
rect 2026 673 2037 676
rect 2018 663 2029 666
rect 2026 653 2029 663
rect 2002 643 2021 646
rect 1994 623 2005 626
rect 1986 613 1997 616
rect 1970 423 1981 426
rect 1962 413 1973 416
rect 1938 353 1949 356
rect 1938 333 1941 353
rect 1946 343 1957 346
rect 1946 333 1957 336
rect 1946 303 1949 333
rect 1954 323 1973 326
rect 1978 316 1981 423
rect 1986 406 1989 546
rect 1994 413 1997 613
rect 2002 573 2005 616
rect 2010 533 2013 636
rect 2018 603 2021 643
rect 2034 596 2037 673
rect 2042 633 2045 786
rect 2018 593 2037 596
rect 2018 493 2021 593
rect 2042 583 2045 616
rect 2034 536 2037 576
rect 2050 573 2053 816
rect 2066 813 2069 953
rect 2082 883 2085 1306
rect 2090 1143 2093 1333
rect 2098 1276 2101 1486
rect 2114 1426 2117 1506
rect 2138 1503 2141 1563
rect 2146 1523 2149 1536
rect 2146 1483 2149 1516
rect 2106 1423 2117 1426
rect 2106 1293 2109 1423
rect 2114 1403 2117 1416
rect 2130 1373 2133 1416
rect 2154 1413 2157 1653
rect 2162 1613 2165 1636
rect 2170 1613 2173 1736
rect 2186 1676 2189 1743
rect 2186 1673 2197 1676
rect 2178 1593 2181 1606
rect 2186 1583 2189 1656
rect 2162 1516 2165 1576
rect 2194 1566 2197 1673
rect 2202 1573 2205 1806
rect 2210 1733 2213 1746
rect 2218 1723 2221 1823
rect 2226 1783 2229 1816
rect 2242 1813 2245 1836
rect 2250 1746 2253 1836
rect 2226 1743 2253 1746
rect 2210 1646 2213 1666
rect 2210 1643 2217 1646
rect 2214 1586 2217 1643
rect 2226 1603 2229 1743
rect 2234 1653 2237 1736
rect 2242 1733 2253 1736
rect 2242 1683 2245 1726
rect 2242 1613 2245 1676
rect 2210 1583 2217 1586
rect 2210 1566 2213 1583
rect 2186 1563 2197 1566
rect 2202 1563 2213 1566
rect 2162 1513 2173 1516
rect 2186 1496 2189 1563
rect 2098 1273 2105 1276
rect 2102 1156 2105 1273
rect 2098 1153 2105 1156
rect 2114 1153 2117 1366
rect 2090 1003 2093 1136
rect 2098 946 2101 1153
rect 2122 1136 2125 1326
rect 2138 1323 2141 1336
rect 2146 1326 2149 1406
rect 2162 1336 2165 1496
rect 2178 1493 2189 1496
rect 2170 1413 2173 1436
rect 2178 1343 2181 1493
rect 2202 1426 2205 1563
rect 2234 1543 2237 1606
rect 2218 1533 2253 1536
rect 2218 1526 2221 1533
rect 2210 1523 2221 1526
rect 2210 1513 2213 1523
rect 2218 1446 2221 1516
rect 2226 1513 2229 1526
rect 2226 1503 2237 1506
rect 2242 1503 2245 1516
rect 2218 1443 2237 1446
rect 2186 1413 2189 1426
rect 2202 1423 2221 1426
rect 2186 1383 2189 1406
rect 2194 1376 2197 1406
rect 2186 1373 2197 1376
rect 2162 1333 2173 1336
rect 2146 1323 2165 1326
rect 2130 1313 2141 1316
rect 2130 1206 2133 1296
rect 2138 1223 2141 1313
rect 2130 1203 2137 1206
rect 2134 1136 2137 1203
rect 2146 1173 2149 1206
rect 2154 1186 2157 1286
rect 2170 1283 2173 1333
rect 2186 1313 2189 1373
rect 2202 1356 2205 1423
rect 2210 1413 2221 1416
rect 2218 1403 2221 1413
rect 2226 1393 2229 1436
rect 2234 1386 2237 1443
rect 2194 1353 2205 1356
rect 2218 1383 2237 1386
rect 2162 1213 2165 1236
rect 2154 1183 2161 1186
rect 2106 1133 2125 1136
rect 2130 1133 2137 1136
rect 2106 1063 2109 1126
rect 2114 1093 2117 1126
rect 2130 1116 2133 1133
rect 2130 1113 2141 1116
rect 2106 953 2109 1026
rect 2122 1023 2125 1106
rect 2114 983 2117 996
rect 2122 993 2125 1016
rect 2130 976 2133 1066
rect 2146 1026 2149 1136
rect 2158 1126 2161 1183
rect 2170 1153 2173 1246
rect 2186 1213 2189 1246
rect 2194 1206 2197 1353
rect 2202 1333 2205 1346
rect 2218 1343 2221 1383
rect 2250 1356 2253 1416
rect 2258 1413 2261 1913
rect 2266 1833 2269 1886
rect 2290 1846 2293 1866
rect 2282 1843 2293 1846
rect 2282 1766 2285 1843
rect 2298 1803 2301 1923
rect 2322 1836 2325 1866
rect 2306 1833 2325 1836
rect 2306 1796 2309 1826
rect 2298 1793 2309 1796
rect 2282 1763 2293 1766
rect 2266 1723 2269 1736
rect 2274 1733 2277 1746
rect 2274 1626 2277 1726
rect 2282 1713 2285 1726
rect 2290 1676 2293 1763
rect 2298 1703 2301 1793
rect 2306 1726 2309 1786
rect 2314 1733 2317 1826
rect 2322 1803 2325 1833
rect 2330 1823 2333 2146
rect 2338 2123 2349 2126
rect 2354 2116 2357 2163
rect 2378 2136 2381 2343
rect 2386 2203 2389 2326
rect 2394 2316 2397 2336
rect 2418 2333 2421 2346
rect 2434 2333 2437 2346
rect 2394 2313 2401 2316
rect 2398 2236 2401 2313
rect 2410 2296 2413 2326
rect 2434 2313 2437 2326
rect 2410 2293 2421 2296
rect 2394 2233 2401 2236
rect 2394 2213 2397 2233
rect 2418 2216 2421 2293
rect 2410 2213 2421 2216
rect 2410 2193 2413 2213
rect 2442 2196 2445 2216
rect 2458 2203 2461 2236
rect 2370 2133 2381 2136
rect 2338 2113 2357 2116
rect 2338 2013 2341 2113
rect 2386 2106 2389 2146
rect 2402 2133 2413 2136
rect 2402 2113 2405 2133
rect 2346 2103 2357 2106
rect 2382 2103 2389 2106
rect 2346 2033 2349 2103
rect 2354 2006 2357 2026
rect 2354 2003 2365 2006
rect 2370 1996 2373 2086
rect 2382 2036 2385 2103
rect 2394 2086 2397 2106
rect 2394 2083 2405 2086
rect 2402 2036 2405 2083
rect 2434 2046 2437 2196
rect 2442 2193 2453 2196
rect 2466 2193 2469 2206
rect 2450 2136 2453 2193
rect 2474 2143 2477 2336
rect 2490 2316 2493 2393
rect 2506 2323 2509 2406
rect 2514 2343 2517 2416
rect 2546 2406 2549 2416
rect 2522 2386 2525 2396
rect 2538 2393 2541 2406
rect 2546 2403 2557 2406
rect 2562 2403 2565 2416
rect 2546 2386 2549 2396
rect 2522 2383 2549 2386
rect 2490 2313 2501 2316
rect 2482 2213 2485 2226
rect 2446 2133 2453 2136
rect 2446 2066 2449 2133
rect 2446 2063 2453 2066
rect 2434 2043 2445 2046
rect 2382 2033 2389 2036
rect 2362 1993 2373 1996
rect 2346 1933 2349 1956
rect 2362 1933 2365 1993
rect 2378 1933 2381 2016
rect 2386 1996 2389 2033
rect 2394 2033 2405 2036
rect 2394 2013 2397 2033
rect 2418 2023 2437 2026
rect 2418 2003 2421 2023
rect 2386 1993 2405 1996
rect 2402 1976 2405 1993
rect 2402 1973 2413 1976
rect 2386 1933 2389 1956
rect 2394 1926 2397 1946
rect 2330 1753 2333 1816
rect 2346 1746 2349 1816
rect 2354 1813 2357 1866
rect 2362 1773 2365 1806
rect 2322 1743 2349 1746
rect 2322 1733 2325 1743
rect 2338 1733 2349 1736
rect 2306 1723 2317 1726
rect 2290 1673 2309 1676
rect 2274 1623 2285 1626
rect 2266 1503 2269 1566
rect 2274 1486 2277 1616
rect 2282 1583 2285 1623
rect 2306 1613 2309 1673
rect 2314 1613 2317 1723
rect 2322 1713 2325 1726
rect 2330 1676 2333 1726
rect 2346 1703 2349 1726
rect 2354 1713 2357 1736
rect 2370 1723 2373 1926
rect 2386 1923 2397 1926
rect 2386 1906 2389 1923
rect 2410 1916 2413 1973
rect 2434 1923 2437 2023
rect 2442 2006 2445 2043
rect 2450 2013 2453 2063
rect 2458 2036 2461 2126
rect 2466 2123 2469 2136
rect 2474 2053 2477 2126
rect 2482 2046 2485 2136
rect 2474 2043 2485 2046
rect 2458 2033 2469 2036
rect 2458 2006 2461 2026
rect 2442 2003 2461 2006
rect 2458 1953 2461 2003
rect 2382 1903 2389 1906
rect 2394 1913 2413 1916
rect 2442 1913 2445 1936
rect 2466 1923 2469 2033
rect 2474 2003 2477 2043
rect 2490 2036 2493 2206
rect 2482 2033 2493 2036
rect 2482 1923 2485 2033
rect 2498 2016 2501 2313
rect 2506 2196 2509 2216
rect 2514 2206 2517 2336
rect 2538 2316 2541 2336
rect 2530 2313 2541 2316
rect 2530 2256 2533 2313
rect 2530 2253 2541 2256
rect 2530 2223 2533 2236
rect 2514 2203 2525 2206
rect 2506 2193 2517 2196
rect 2530 2193 2533 2216
rect 2538 2213 2541 2253
rect 2546 2206 2549 2383
rect 2554 2333 2557 2403
rect 2570 2383 2573 2416
rect 2618 2413 2629 2416
rect 2618 2353 2621 2406
rect 2634 2393 2637 2406
rect 2578 2333 2581 2346
rect 2562 2313 2565 2326
rect 2570 2283 2573 2326
rect 2586 2293 2589 2326
rect 2594 2313 2597 2336
rect 2634 2316 2637 2336
rect 2626 2313 2637 2316
rect 2626 2256 2629 2313
rect 2642 2276 2645 2386
rect 2658 2356 2661 2426
rect 2658 2353 2669 2356
rect 2650 2323 2653 2346
rect 2642 2273 2653 2276
rect 2626 2253 2637 2256
rect 2514 2176 2517 2193
rect 2514 2173 2521 2176
rect 2538 2173 2541 2206
rect 2546 2203 2581 2206
rect 2586 2176 2589 2236
rect 2594 2223 2597 2236
rect 2554 2173 2589 2176
rect 2506 2083 2509 2146
rect 2518 2096 2521 2173
rect 2538 2133 2541 2146
rect 2554 2133 2557 2173
rect 2562 2126 2565 2166
rect 2530 2123 2541 2126
rect 2546 2113 2549 2126
rect 2554 2123 2565 2126
rect 2570 2123 2573 2173
rect 2514 2093 2521 2096
rect 2514 2076 2517 2093
rect 2494 2013 2501 2016
rect 2506 2073 2517 2076
rect 2382 1836 2385 1903
rect 2382 1833 2389 1836
rect 2322 1673 2333 1676
rect 2290 1553 2293 1596
rect 2322 1556 2325 1673
rect 2314 1553 2325 1556
rect 2282 1543 2309 1546
rect 2282 1523 2285 1543
rect 2290 1506 2293 1536
rect 2298 1523 2301 1536
rect 2314 1533 2317 1553
rect 2322 1533 2325 1546
rect 2330 1513 2333 1666
rect 2370 1623 2373 1666
rect 2378 1623 2381 1806
rect 2386 1773 2389 1833
rect 2394 1823 2397 1913
rect 2402 1833 2405 1886
rect 2418 1806 2421 1826
rect 2386 1693 2389 1736
rect 2338 1593 2341 1606
rect 2346 1603 2381 1606
rect 2346 1516 2349 1526
rect 2354 1523 2357 1586
rect 2370 1533 2373 1556
rect 2346 1513 2373 1516
rect 2378 1513 2381 1536
rect 2270 1483 2277 1486
rect 2246 1353 2253 1356
rect 2218 1293 2221 1336
rect 2226 1323 2237 1326
rect 2226 1276 2229 1316
rect 2218 1273 2229 1276
rect 2218 1256 2221 1273
rect 2214 1253 2221 1256
rect 2202 1213 2205 1236
rect 2178 1126 2181 1206
rect 2186 1203 2197 1206
rect 2186 1133 2189 1203
rect 2214 1196 2217 1253
rect 2226 1203 2229 1266
rect 2214 1193 2221 1196
rect 2202 1133 2205 1146
rect 2158 1123 2173 1126
rect 2178 1123 2197 1126
rect 2154 1033 2157 1066
rect 2146 1023 2157 1026
rect 2126 973 2133 976
rect 2098 943 2109 946
rect 2098 916 2101 936
rect 2094 913 2101 916
rect 2074 873 2085 876
rect 2082 813 2085 873
rect 2094 846 2097 913
rect 2106 856 2109 943
rect 2114 873 2117 936
rect 2126 906 2129 973
rect 2138 913 2141 1006
rect 2146 983 2149 1016
rect 2154 956 2157 1023
rect 2162 963 2165 1116
rect 2170 1056 2173 1123
rect 2210 1093 2213 1126
rect 2218 1076 2221 1193
rect 2194 1073 2221 1076
rect 2170 1053 2189 1056
rect 2170 1003 2173 1046
rect 2154 953 2173 956
rect 2146 933 2157 936
rect 2126 903 2133 906
rect 2106 853 2113 856
rect 2094 843 2101 846
rect 2058 783 2061 806
rect 2066 803 2077 806
rect 2090 803 2093 826
rect 2058 553 2061 746
rect 2066 733 2069 756
rect 2066 696 2069 726
rect 2074 723 2077 776
rect 2082 723 2085 736
rect 2066 693 2077 696
rect 2074 626 2077 693
rect 2090 663 2093 726
rect 2098 713 2101 843
rect 2110 776 2113 853
rect 2106 773 2113 776
rect 2066 623 2077 626
rect 2066 603 2069 623
rect 2034 533 2045 536
rect 2034 513 2037 526
rect 2042 503 2045 533
rect 2066 506 2069 586
rect 2082 583 2085 606
rect 2090 566 2093 636
rect 2098 603 2101 616
rect 2074 563 2093 566
rect 2074 516 2077 563
rect 2082 523 2085 556
rect 2090 533 2101 536
rect 2106 526 2109 773
rect 2114 733 2117 756
rect 2122 743 2125 886
rect 2122 703 2125 726
rect 2130 686 2133 903
rect 2146 893 2149 926
rect 2154 923 2165 926
rect 2138 803 2141 876
rect 2146 783 2149 806
rect 2138 733 2149 736
rect 2138 693 2141 733
rect 2130 683 2141 686
rect 2114 533 2117 576
rect 2122 536 2125 606
rect 2130 593 2133 616
rect 2122 533 2133 536
rect 2098 516 2101 526
rect 2106 523 2117 526
rect 2074 513 2101 516
rect 2066 503 2085 506
rect 2002 413 2005 436
rect 2010 406 2013 426
rect 1986 403 2013 406
rect 1986 333 1989 403
rect 2018 386 2021 446
rect 2034 413 2037 446
rect 2042 433 2061 436
rect 2050 406 2053 426
rect 2058 423 2061 433
rect 2066 423 2069 496
rect 2082 406 2085 503
rect 2114 466 2117 523
rect 2114 463 2125 466
rect 2090 413 2093 446
rect 2010 383 2021 386
rect 2026 403 2053 406
rect 2010 326 2013 383
rect 2026 333 2029 403
rect 1962 313 1981 316
rect 1938 153 1941 196
rect 1866 113 1869 126
rect 1946 123 1949 206
rect 1954 113 1957 136
rect 1962 123 1965 313
rect 1994 293 1997 326
rect 2010 323 2021 326
rect 1970 206 1973 216
rect 1978 213 1981 246
rect 2010 213 2013 226
rect 2018 213 2021 323
rect 2050 273 2053 326
rect 2058 293 2061 336
rect 2066 323 2069 406
rect 2082 403 2093 406
rect 2090 376 2093 403
rect 2082 373 2093 376
rect 2082 326 2085 373
rect 2114 366 2117 426
rect 2122 403 2125 463
rect 2098 333 2101 366
rect 2106 363 2117 366
rect 2106 333 2109 363
rect 2130 353 2133 533
rect 2138 413 2141 683
rect 2146 633 2149 726
rect 2146 523 2149 616
rect 2154 593 2157 916
rect 2162 883 2165 923
rect 2170 903 2173 953
rect 2162 823 2173 826
rect 2162 703 2165 726
rect 2170 713 2173 823
rect 2178 786 2181 1016
rect 2186 843 2189 1053
rect 2186 803 2189 816
rect 2178 783 2185 786
rect 2170 683 2173 706
rect 2182 676 2185 783
rect 2178 673 2185 676
rect 2170 583 2173 596
rect 2170 533 2173 546
rect 2178 486 2181 673
rect 2186 603 2189 616
rect 2194 576 2197 1073
rect 2202 1013 2205 1026
rect 2210 996 2213 1006
rect 2218 1003 2221 1066
rect 2226 996 2229 1126
rect 2234 1083 2237 1316
rect 2246 1256 2249 1353
rect 2258 1313 2261 1346
rect 2270 1296 2273 1483
rect 2282 1413 2285 1506
rect 2290 1503 2301 1506
rect 2298 1436 2301 1503
rect 2290 1433 2301 1436
rect 2282 1323 2285 1406
rect 2270 1293 2277 1296
rect 2246 1253 2253 1256
rect 2242 1213 2245 1236
rect 2242 1036 2245 1136
rect 2210 993 2229 996
rect 2238 1033 2245 1036
rect 2202 623 2205 946
rect 2210 933 2213 966
rect 2218 933 2221 993
rect 2238 986 2241 1033
rect 2234 983 2241 986
rect 2210 866 2213 926
rect 2226 913 2229 926
rect 2210 863 2221 866
rect 2202 586 2205 616
rect 2210 596 2213 856
rect 2218 813 2221 863
rect 2226 856 2229 876
rect 2234 863 2237 983
rect 2250 953 2253 1253
rect 2258 1223 2261 1276
rect 2274 1273 2277 1293
rect 2282 1183 2285 1206
rect 2282 1133 2285 1166
rect 2258 1093 2261 1126
rect 2258 1003 2261 1076
rect 2242 893 2245 926
rect 2258 913 2261 936
rect 2258 886 2261 906
rect 2254 883 2261 886
rect 2226 853 2237 856
rect 2234 806 2237 853
rect 2254 826 2257 883
rect 2266 833 2269 1086
rect 2274 1073 2277 1126
rect 2290 1116 2293 1433
rect 2386 1426 2389 1526
rect 2394 1493 2397 1806
rect 2410 1803 2421 1806
rect 2410 1736 2413 1803
rect 2410 1733 2421 1736
rect 2410 1696 2413 1716
rect 2402 1693 2413 1696
rect 2402 1623 2405 1693
rect 2418 1636 2421 1733
rect 2426 1696 2429 1846
rect 2494 1836 2497 2013
rect 2506 1973 2509 2073
rect 2514 1996 2517 2036
rect 2530 2023 2549 2026
rect 2530 1996 2533 2006
rect 2514 1993 2533 1996
rect 2538 1983 2541 1996
rect 2506 1933 2509 1946
rect 2506 1883 2509 1926
rect 2546 1916 2549 2023
rect 2554 2013 2557 2123
rect 2570 2016 2573 2116
rect 2562 2013 2573 2016
rect 2514 1913 2549 1916
rect 2442 1833 2461 1836
rect 2490 1833 2497 1836
rect 2538 1833 2541 1906
rect 2554 1896 2557 1936
rect 2550 1893 2557 1896
rect 2550 1836 2553 1893
rect 2550 1833 2557 1836
rect 2434 1753 2437 1816
rect 2450 1736 2453 1826
rect 2466 1783 2469 1826
rect 2474 1753 2477 1816
rect 2490 1766 2493 1833
rect 2506 1823 2533 1826
rect 2490 1763 2501 1766
rect 2434 1733 2453 1736
rect 2434 1716 2437 1726
rect 2458 1716 2461 1746
rect 2474 1723 2477 1736
rect 2490 1733 2493 1746
rect 2498 1726 2501 1763
rect 2506 1733 2509 1823
rect 2522 1786 2525 1816
rect 2530 1803 2533 1823
rect 2554 1813 2557 1833
rect 2530 1793 2541 1796
rect 2554 1793 2557 1806
rect 2522 1783 2541 1786
rect 2522 1733 2525 1756
rect 2538 1733 2541 1783
rect 2562 1746 2565 2013
rect 2586 1956 2589 2066
rect 2594 2056 2597 2216
rect 2602 2203 2613 2206
rect 2602 2183 2605 2203
rect 2618 2173 2621 2236
rect 2626 2223 2629 2236
rect 2610 2133 2613 2146
rect 2634 2123 2637 2253
rect 2650 2176 2653 2273
rect 2646 2173 2653 2176
rect 2594 2053 2613 2056
rect 2610 1996 2613 2053
rect 2634 2013 2637 2116
rect 2646 2096 2649 2173
rect 2666 2166 2669 2353
rect 2658 2163 2669 2166
rect 2658 2136 2661 2163
rect 2658 2133 2669 2136
rect 2658 2113 2661 2126
rect 2646 2093 2653 2096
rect 2570 1953 2589 1956
rect 2602 1993 2613 1996
rect 2570 1866 2573 1953
rect 2578 1933 2581 1946
rect 2594 1936 2597 1946
rect 2586 1933 2597 1936
rect 2602 1923 2605 1993
rect 2650 1966 2653 2093
rect 2666 2036 2669 2133
rect 2642 1963 2653 1966
rect 2662 2033 2669 2036
rect 2642 1866 2645 1963
rect 2662 1956 2665 2033
rect 2658 1953 2665 1956
rect 2570 1863 2589 1866
rect 2642 1863 2653 1866
rect 2578 1836 2581 1856
rect 2570 1833 2581 1836
rect 2562 1743 2569 1746
rect 2578 1743 2581 1756
rect 2490 1723 2501 1726
rect 2506 1723 2533 1726
rect 2434 1713 2461 1716
rect 2426 1693 2433 1696
rect 2410 1633 2421 1636
rect 2410 1616 2413 1633
rect 2430 1626 2433 1693
rect 2402 1613 2413 1616
rect 2418 1613 2421 1626
rect 2426 1623 2433 1626
rect 2402 1453 2405 1613
rect 2410 1496 2413 1606
rect 2418 1553 2421 1606
rect 2418 1513 2421 1526
rect 2410 1493 2417 1496
rect 2354 1423 2389 1426
rect 2298 1413 2309 1416
rect 2354 1413 2357 1423
rect 2378 1413 2389 1416
rect 2298 1396 2301 1406
rect 2306 1403 2317 1406
rect 2322 1396 2325 1406
rect 2298 1393 2325 1396
rect 2298 1373 2341 1376
rect 2298 1333 2301 1373
rect 2322 1353 2333 1356
rect 2330 1323 2333 1353
rect 2314 1296 2317 1316
rect 2338 1313 2341 1373
rect 2346 1323 2349 1406
rect 2386 1363 2389 1413
rect 2394 1403 2397 1426
rect 2402 1413 2405 1436
rect 2414 1426 2417 1493
rect 2410 1423 2417 1426
rect 2402 1306 2405 1326
rect 2306 1293 2317 1296
rect 2330 1293 2333 1306
rect 2394 1303 2405 1306
rect 2410 1306 2413 1423
rect 2418 1323 2421 1406
rect 2426 1366 2429 1623
rect 2434 1563 2437 1606
rect 2442 1586 2445 1706
rect 2450 1693 2453 1706
rect 2490 1636 2493 1723
rect 2474 1633 2493 1636
rect 2450 1593 2453 1606
rect 2442 1583 2453 1586
rect 2434 1506 2437 1536
rect 2442 1533 2445 1546
rect 2434 1503 2441 1506
rect 2438 1436 2441 1503
rect 2434 1433 2441 1436
rect 2434 1413 2437 1433
rect 2450 1416 2453 1583
rect 2442 1413 2453 1416
rect 2434 1383 2437 1396
rect 2426 1363 2433 1366
rect 2430 1316 2433 1363
rect 2426 1313 2433 1316
rect 2410 1303 2417 1306
rect 2286 1113 2293 1116
rect 2286 1056 2289 1113
rect 2298 1103 2301 1176
rect 2274 1053 2289 1056
rect 2254 823 2261 826
rect 2218 713 2221 806
rect 2234 803 2253 806
rect 2218 703 2229 706
rect 2234 703 2237 716
rect 2218 603 2221 703
rect 2242 696 2245 746
rect 2250 723 2253 803
rect 2258 763 2261 823
rect 2266 746 2269 826
rect 2258 743 2269 746
rect 2274 743 2277 1053
rect 2282 986 2285 1046
rect 2306 1043 2309 1293
rect 2314 1183 2317 1216
rect 2314 1123 2317 1146
rect 2314 1103 2317 1116
rect 2314 1033 2317 1066
rect 2290 1003 2317 1006
rect 2282 983 2289 986
rect 2286 866 2289 983
rect 2306 973 2309 996
rect 2298 933 2309 936
rect 2298 903 2301 926
rect 2306 916 2309 926
rect 2314 923 2317 1003
rect 2322 916 2325 1286
rect 2394 1256 2397 1303
rect 2394 1253 2405 1256
rect 2330 1203 2333 1246
rect 2338 1233 2389 1236
rect 2338 1223 2341 1233
rect 2346 1223 2357 1226
rect 2338 1193 2341 1206
rect 2306 913 2325 916
rect 2330 896 2333 1166
rect 2346 1113 2349 1146
rect 2354 1136 2357 1223
rect 2362 1213 2373 1216
rect 2386 1213 2389 1233
rect 2402 1213 2405 1253
rect 2414 1236 2417 1303
rect 2410 1233 2417 1236
rect 2362 1193 2365 1206
rect 2394 1176 2397 1206
rect 2370 1173 2397 1176
rect 2354 1133 2365 1136
rect 2370 1133 2373 1173
rect 2362 1126 2365 1133
rect 2338 1043 2341 1106
rect 2354 1093 2357 1126
rect 2362 1123 2381 1126
rect 2362 1096 2365 1116
rect 2362 1093 2369 1096
rect 2346 1036 2349 1086
rect 2338 1033 2349 1036
rect 2338 1023 2341 1033
rect 2354 1016 2357 1046
rect 2338 1013 2357 1016
rect 2338 983 2341 1013
rect 2366 1006 2369 1093
rect 2362 1003 2369 1006
rect 2282 863 2289 866
rect 2326 893 2333 896
rect 2282 846 2285 863
rect 2282 843 2317 846
rect 2282 833 2285 843
rect 2226 693 2245 696
rect 2226 623 2229 693
rect 2250 683 2253 706
rect 2258 616 2261 743
rect 2266 693 2269 716
rect 2274 703 2277 716
rect 2282 636 2285 716
rect 2290 693 2293 766
rect 2274 633 2285 636
rect 2298 633 2301 836
rect 2314 766 2317 843
rect 2306 763 2317 766
rect 2306 683 2309 763
rect 2326 746 2329 893
rect 2338 813 2341 936
rect 2346 913 2349 966
rect 2362 946 2365 1003
rect 2354 943 2365 946
rect 2346 813 2349 826
rect 2314 743 2329 746
rect 2338 803 2349 806
rect 2234 613 2261 616
rect 2210 593 2237 596
rect 2202 583 2213 586
rect 2194 573 2205 576
rect 2186 496 2189 526
rect 2194 513 2197 546
rect 2202 523 2205 573
rect 2210 516 2213 583
rect 2202 513 2213 516
rect 2186 493 2197 496
rect 2178 483 2189 486
rect 2146 413 2149 426
rect 2170 406 2173 466
rect 2186 413 2189 483
rect 2154 403 2173 406
rect 2170 346 2173 403
rect 2178 363 2181 406
rect 2194 383 2197 493
rect 2114 343 2141 346
rect 2082 323 2093 326
rect 2090 223 2093 323
rect 1970 203 2029 206
rect 2074 203 2093 206
rect 2002 103 2005 136
rect 2026 123 2029 203
rect 2034 123 2037 196
rect 2082 113 2085 126
rect 2090 113 2093 203
rect 2098 103 2101 216
rect 2106 186 2109 216
rect 2114 193 2117 343
rect 2138 336 2141 343
rect 2130 323 2133 336
rect 2138 333 2157 336
rect 2138 303 2141 326
rect 2130 213 2133 296
rect 2146 263 2149 326
rect 2162 323 2165 346
rect 2170 343 2181 346
rect 2170 303 2173 336
rect 2178 323 2181 336
rect 2202 306 2205 513
rect 2234 506 2237 593
rect 2242 513 2245 526
rect 2250 513 2253 536
rect 2210 503 2229 506
rect 2234 503 2245 506
rect 2242 426 2245 503
rect 2258 433 2261 613
rect 2266 623 2293 626
rect 2266 606 2269 623
rect 2266 603 2273 606
rect 2270 526 2273 603
rect 2266 523 2273 526
rect 2282 523 2285 616
rect 2298 586 2301 606
rect 2294 583 2301 586
rect 2294 526 2297 583
rect 2306 533 2309 646
rect 2314 606 2317 743
rect 2338 736 2341 803
rect 2322 733 2333 736
rect 2338 733 2349 736
rect 2322 713 2325 733
rect 2354 716 2357 943
rect 2346 713 2357 716
rect 2322 613 2325 696
rect 2330 613 2333 706
rect 2346 646 2349 713
rect 2346 643 2353 646
rect 2362 643 2365 866
rect 2370 803 2373 936
rect 2378 933 2381 1123
rect 2386 1003 2389 1116
rect 2394 1103 2397 1173
rect 2402 1113 2405 1196
rect 2410 1053 2413 1233
rect 2426 1226 2429 1313
rect 2426 1223 2437 1226
rect 2418 1213 2429 1216
rect 2418 1046 2421 1196
rect 2434 1116 2437 1223
rect 2442 1193 2445 1413
rect 2450 1373 2453 1406
rect 2450 1213 2453 1226
rect 2450 1133 2453 1206
rect 2458 1203 2461 1566
rect 2466 1513 2469 1536
rect 2474 1503 2477 1633
rect 2482 1613 2485 1626
rect 2490 1613 2493 1633
rect 2482 1543 2485 1556
rect 2490 1516 2493 1606
rect 2498 1583 2501 1606
rect 2506 1563 2509 1723
rect 2554 1683 2557 1736
rect 2566 1696 2569 1743
rect 2586 1736 2589 1863
rect 2562 1693 2569 1696
rect 2578 1733 2589 1736
rect 2634 1733 2637 1816
rect 2642 1733 2645 1746
rect 2562 1673 2565 1693
rect 2514 1603 2517 1626
rect 2522 1613 2525 1636
rect 2506 1523 2509 1546
rect 2490 1513 2501 1516
rect 2498 1436 2501 1513
rect 2514 1446 2517 1576
rect 2522 1533 2525 1546
rect 2514 1443 2521 1446
rect 2498 1433 2509 1436
rect 2466 1413 2469 1426
rect 2482 1413 2501 1416
rect 2506 1406 2509 1433
rect 2466 1393 2469 1406
rect 2482 1393 2485 1406
rect 2498 1403 2509 1406
rect 2474 1213 2477 1366
rect 2498 1316 2501 1403
rect 2518 1396 2521 1443
rect 2530 1413 2533 1646
rect 2578 1636 2581 1733
rect 2586 1723 2605 1726
rect 2578 1633 2589 1636
rect 2538 1603 2541 1626
rect 2578 1543 2581 1586
rect 2586 1536 2589 1633
rect 2634 1603 2637 1616
rect 2546 1523 2549 1536
rect 2570 1533 2589 1536
rect 2642 1533 2645 1546
rect 2514 1393 2521 1396
rect 2514 1336 2517 1393
rect 2530 1373 2533 1406
rect 2538 1346 2541 1506
rect 2554 1413 2557 1426
rect 2562 1413 2565 1446
rect 2570 1436 2573 1533
rect 2578 1523 2597 1526
rect 2570 1433 2589 1436
rect 2546 1356 2549 1406
rect 2554 1393 2557 1406
rect 2546 1353 2565 1356
rect 2538 1343 2549 1346
rect 2506 1333 2517 1336
rect 2514 1323 2533 1326
rect 2498 1313 2533 1316
rect 2466 1193 2469 1206
rect 2482 1203 2485 1226
rect 2498 1196 2501 1313
rect 2538 1263 2541 1336
rect 2546 1326 2549 1343
rect 2546 1323 2553 1326
rect 2550 1266 2553 1323
rect 2546 1263 2553 1266
rect 2482 1193 2501 1196
rect 2458 1116 2461 1136
rect 2402 1043 2421 1046
rect 2394 983 2397 1016
rect 2402 1013 2405 1043
rect 2426 1013 2429 1116
rect 2434 1113 2445 1116
rect 2450 1113 2461 1116
rect 2434 1083 2437 1106
rect 2442 1076 2445 1113
rect 2466 1106 2469 1166
rect 2462 1103 2469 1106
rect 2442 1073 2453 1076
rect 2442 1013 2445 1066
rect 2402 973 2405 1006
rect 2418 1003 2429 1006
rect 2434 983 2437 1006
rect 2442 956 2445 1006
rect 2450 963 2453 1073
rect 2462 1026 2465 1103
rect 2458 1023 2465 1026
rect 2458 1003 2461 1023
rect 2466 983 2469 1006
rect 2442 953 2453 956
rect 2378 903 2381 926
rect 2402 913 2405 936
rect 2426 906 2429 926
rect 2434 923 2437 946
rect 2418 903 2429 906
rect 2418 846 2421 903
rect 2418 843 2429 846
rect 2378 773 2381 816
rect 2394 736 2397 766
rect 2402 746 2405 816
rect 2402 743 2413 746
rect 2370 693 2373 726
rect 2378 646 2381 736
rect 2386 733 2397 736
rect 2370 643 2381 646
rect 2394 686 2397 726
rect 2402 693 2405 736
rect 2410 733 2413 743
rect 2418 686 2421 826
rect 2426 803 2429 843
rect 2426 783 2429 796
rect 2426 723 2429 746
rect 2394 683 2421 686
rect 2338 613 2341 626
rect 2314 603 2333 606
rect 2330 533 2333 603
rect 2338 533 2341 606
rect 2350 596 2353 643
rect 2362 603 2365 626
rect 2350 593 2357 596
rect 2294 523 2301 526
rect 2314 523 2325 526
rect 2266 433 2269 523
rect 2210 423 2245 426
rect 2210 326 2213 423
rect 2234 403 2237 416
rect 2242 413 2245 423
rect 2250 423 2269 426
rect 2250 406 2253 423
rect 2242 403 2253 406
rect 2242 396 2245 403
rect 2226 393 2245 396
rect 2218 333 2221 386
rect 2266 356 2269 423
rect 2282 403 2285 516
rect 2298 383 2301 523
rect 2338 513 2341 526
rect 2314 416 2317 506
rect 2310 413 2317 416
rect 2266 353 2277 356
rect 2274 333 2277 353
rect 2282 333 2285 356
rect 2310 336 2313 413
rect 2322 386 2325 486
rect 2354 426 2357 593
rect 2370 583 2373 643
rect 2378 593 2381 636
rect 2394 626 2397 683
rect 2434 676 2437 896
rect 2442 813 2445 906
rect 2450 893 2453 953
rect 2474 886 2477 1156
rect 2482 1116 2485 1193
rect 2482 1113 2493 1116
rect 2490 1066 2493 1113
rect 2506 1093 2509 1126
rect 2514 1116 2517 1196
rect 2530 1193 2533 1216
rect 2538 1213 2541 1236
rect 2546 1146 2549 1263
rect 2562 1246 2565 1353
rect 2554 1243 2565 1246
rect 2554 1206 2557 1243
rect 2562 1213 2565 1226
rect 2554 1203 2565 1206
rect 2562 1146 2565 1203
rect 2586 1163 2589 1433
rect 2610 1413 2613 1426
rect 2610 1323 2613 1336
rect 2610 1213 2613 1226
rect 2578 1153 2605 1156
rect 2522 1123 2525 1146
rect 2546 1143 2553 1146
rect 2562 1143 2573 1146
rect 2530 1133 2541 1136
rect 2530 1116 2533 1126
rect 2514 1113 2533 1116
rect 2538 1073 2541 1133
rect 2550 1086 2553 1143
rect 2546 1083 2553 1086
rect 2546 1066 2549 1083
rect 2482 1063 2493 1066
rect 2530 1063 2549 1066
rect 2482 1043 2485 1063
rect 2490 1013 2501 1016
rect 2482 983 2485 996
rect 2490 973 2493 1006
rect 2506 1003 2509 1026
rect 2514 966 2517 1056
rect 2530 986 2533 1063
rect 2538 1013 2557 1016
rect 2562 1013 2565 1136
rect 2570 1116 2573 1143
rect 2578 1123 2581 1153
rect 2570 1113 2589 1116
rect 2594 1113 2597 1146
rect 2602 1123 2605 1153
rect 2610 1133 2613 1146
rect 2618 1136 2621 1416
rect 2650 1336 2653 1863
rect 2658 1506 2661 1953
rect 2674 1943 2677 2016
rect 2674 1793 2677 1816
rect 2674 1723 2677 1736
rect 2666 1613 2669 1626
rect 2666 1523 2669 1606
rect 2658 1503 2669 1506
rect 2666 1436 2669 1503
rect 2658 1433 2669 1436
rect 2658 1403 2661 1433
rect 2666 1393 2669 1416
rect 2642 1333 2653 1336
rect 2642 1266 2645 1333
rect 2642 1263 2653 1266
rect 2650 1246 2653 1263
rect 2650 1243 2657 1246
rect 2654 1176 2657 1243
rect 2666 1213 2669 1326
rect 2650 1173 2657 1176
rect 2618 1133 2629 1136
rect 2634 1133 2637 1146
rect 2586 1026 2589 1113
rect 2618 1046 2621 1133
rect 2578 1023 2589 1026
rect 2610 1043 2621 1046
rect 2634 1046 2637 1116
rect 2634 1043 2645 1046
rect 2538 993 2541 1006
rect 2530 983 2549 986
rect 2498 946 2501 966
rect 2514 963 2521 966
rect 2494 943 2501 946
rect 2482 903 2485 926
rect 2454 883 2477 886
rect 2494 886 2497 943
rect 2518 886 2521 963
rect 2530 913 2533 926
rect 2494 883 2501 886
rect 2454 816 2457 883
rect 2450 813 2457 816
rect 2466 816 2469 836
rect 2498 816 2501 883
rect 2466 813 2477 816
rect 2442 723 2445 766
rect 2418 673 2437 676
rect 2386 623 2397 626
rect 2338 413 2341 426
rect 2354 423 2361 426
rect 2330 403 2341 406
rect 2346 403 2349 416
rect 2322 383 2333 386
rect 2330 336 2333 383
rect 2358 366 2361 423
rect 2370 403 2373 526
rect 2378 513 2381 526
rect 2386 496 2389 623
rect 2382 493 2389 496
rect 2354 363 2361 366
rect 2310 333 2317 336
rect 2210 323 2221 326
rect 2218 306 2221 323
rect 2194 303 2205 306
rect 2214 303 2221 306
rect 2106 183 2141 186
rect 2114 103 2117 126
rect 2138 123 2141 183
rect 2146 133 2149 256
rect 2194 236 2197 303
rect 2214 236 2217 303
rect 2234 296 2237 326
rect 2194 233 2205 236
rect 2178 203 2181 216
rect 2178 183 2181 196
rect 2202 183 2205 233
rect 2210 233 2217 236
rect 2226 293 2237 296
rect 2210 213 2213 233
rect 2218 203 2221 226
rect 2226 173 2229 293
rect 2266 286 2269 326
rect 2282 303 2285 316
rect 2314 313 2317 333
rect 2322 333 2333 336
rect 2322 313 2325 333
rect 2234 283 2269 286
rect 2234 213 2237 283
rect 2242 223 2253 226
rect 2314 216 2317 226
rect 2250 203 2253 216
rect 2282 213 2317 216
rect 2274 196 2277 206
rect 2282 203 2285 213
rect 2298 196 2301 206
rect 2314 203 2317 213
rect 2274 193 2301 196
rect 2346 186 2349 356
rect 2354 343 2357 363
rect 2382 356 2385 493
rect 2382 353 2389 356
rect 2362 333 2381 336
rect 2362 303 2365 333
rect 2386 326 2389 353
rect 2378 323 2389 326
rect 2370 303 2373 316
rect 2234 143 2253 146
rect 2242 123 2253 126
rect 2258 123 2261 136
rect 2274 126 2277 186
rect 2330 183 2349 186
rect 2354 186 2357 216
rect 2362 203 2365 216
rect 2378 213 2381 323
rect 2394 223 2397 616
rect 2402 586 2405 656
rect 2418 603 2421 673
rect 2402 583 2413 586
rect 2402 463 2405 536
rect 2410 503 2413 583
rect 2418 566 2421 586
rect 2418 563 2425 566
rect 2422 496 2425 563
rect 2434 503 2437 516
rect 2442 513 2445 596
rect 2450 563 2453 813
rect 2458 743 2461 796
rect 2474 746 2477 813
rect 2466 743 2477 746
rect 2490 813 2501 816
rect 2514 883 2521 886
rect 2514 813 2517 883
rect 2490 746 2493 813
rect 2506 766 2509 806
rect 2514 793 2517 806
rect 2522 803 2525 816
rect 2538 813 2541 916
rect 2538 783 2541 806
rect 2506 763 2517 766
rect 2490 743 2501 746
rect 2466 653 2469 743
rect 2482 646 2485 706
rect 2490 673 2493 726
rect 2482 643 2489 646
rect 2466 526 2469 616
rect 2486 566 2489 643
rect 2498 576 2501 743
rect 2506 703 2509 726
rect 2506 613 2509 626
rect 2514 593 2517 616
rect 2522 576 2525 776
rect 2530 733 2541 736
rect 2546 726 2549 983
rect 2554 893 2557 1006
rect 2562 993 2565 1006
rect 2562 923 2565 946
rect 2578 936 2581 1023
rect 2594 946 2597 1016
rect 2610 1013 2613 1043
rect 2610 983 2613 1006
rect 2594 943 2613 946
rect 2578 933 2589 936
rect 2562 886 2565 906
rect 2554 823 2557 886
rect 2562 883 2569 886
rect 2578 883 2581 916
rect 2566 816 2569 883
rect 2578 823 2581 836
rect 2562 813 2569 816
rect 2554 733 2557 766
rect 2538 723 2549 726
rect 2538 616 2541 723
rect 2498 573 2509 576
rect 2486 563 2493 566
rect 2474 543 2477 556
rect 2466 523 2477 526
rect 2418 493 2425 496
rect 2410 403 2413 416
rect 2418 386 2421 493
rect 2426 456 2429 476
rect 2426 453 2433 456
rect 2410 383 2421 386
rect 2410 316 2413 383
rect 2430 356 2433 453
rect 2426 353 2433 356
rect 2426 323 2429 353
rect 2410 313 2421 316
rect 2370 193 2373 206
rect 2386 186 2389 206
rect 2418 203 2421 313
rect 2442 306 2445 416
rect 2434 303 2445 306
rect 2450 316 2453 346
rect 2458 333 2461 506
rect 2466 503 2469 516
rect 2474 413 2477 523
rect 2482 413 2485 516
rect 2466 323 2469 336
rect 2474 316 2477 336
rect 2450 313 2477 316
rect 2434 236 2437 303
rect 2450 256 2453 313
rect 2482 306 2485 396
rect 2490 376 2493 563
rect 2506 506 2509 573
rect 2498 503 2509 506
rect 2518 573 2525 576
rect 2530 613 2541 616
rect 2554 613 2557 646
rect 2498 483 2501 503
rect 2518 476 2521 573
rect 2530 486 2533 613
rect 2538 593 2541 606
rect 2546 593 2557 596
rect 2546 553 2549 593
rect 2538 493 2541 526
rect 2546 523 2549 536
rect 2530 483 2549 486
rect 2498 473 2521 476
rect 2498 393 2501 473
rect 2530 423 2533 436
rect 2546 426 2549 483
rect 2554 433 2557 586
rect 2562 503 2565 813
rect 2578 803 2581 816
rect 2570 506 2573 796
rect 2586 773 2589 933
rect 2594 903 2597 926
rect 2594 733 2597 896
rect 2602 806 2605 936
rect 2610 916 2613 943
rect 2618 933 2621 1036
rect 2626 1023 2629 1036
rect 2610 913 2617 916
rect 2614 846 2617 913
rect 2610 843 2617 846
rect 2610 813 2613 843
rect 2626 826 2629 946
rect 2634 943 2637 1026
rect 2642 1013 2645 1043
rect 2618 823 2629 826
rect 2618 806 2621 823
rect 2602 803 2621 806
rect 2578 713 2581 726
rect 2602 643 2605 803
rect 2610 743 2613 776
rect 2626 753 2629 816
rect 2642 813 2645 826
rect 2634 756 2637 806
rect 2650 796 2653 1173
rect 2658 1023 2661 1036
rect 2666 1006 2669 1126
rect 2662 1003 2669 1006
rect 2662 826 2665 1003
rect 2662 823 2669 826
rect 2666 803 2669 823
rect 2650 793 2669 796
rect 2634 753 2653 756
rect 2578 513 2581 536
rect 2570 503 2581 506
rect 2578 433 2581 503
rect 2586 426 2589 616
rect 2618 613 2621 726
rect 2634 713 2637 736
rect 2642 733 2645 746
rect 2650 726 2653 753
rect 2650 723 2661 726
rect 2666 703 2669 793
rect 2666 593 2669 616
rect 2642 536 2645 556
rect 2594 513 2597 536
rect 2626 516 2629 536
rect 2618 513 2629 516
rect 2638 533 2645 536
rect 2594 486 2597 506
rect 2594 483 2605 486
rect 2602 426 2605 483
rect 2618 456 2621 513
rect 2618 453 2629 456
rect 2538 406 2541 426
rect 2546 423 2557 426
rect 2506 403 2541 406
rect 2490 373 2497 376
rect 2494 316 2497 373
rect 2506 323 2509 403
rect 2530 333 2533 356
rect 2514 316 2517 326
rect 2546 316 2549 336
rect 2494 313 2517 316
rect 2474 303 2485 306
rect 2450 253 2461 256
rect 2434 233 2445 236
rect 2354 183 2389 186
rect 2282 133 2285 166
rect 2274 123 2285 126
rect 2290 123 2293 136
rect 2298 123 2301 136
rect 2330 126 2333 183
rect 2394 176 2397 196
rect 2434 193 2437 216
rect 2442 203 2445 233
rect 2450 203 2453 216
rect 2346 173 2397 176
rect 2346 133 2349 173
rect 2330 123 2341 126
rect 2354 123 2357 146
rect 2362 133 2365 166
rect 2410 133 2413 156
rect 2434 143 2437 186
rect 2154 113 2189 116
rect 2338 103 2341 123
rect 2370 103 2373 126
rect 2458 123 2461 253
rect 2474 236 2477 303
rect 2466 233 2477 236
rect 2466 163 2469 233
rect 2514 226 2517 313
rect 2538 313 2549 316
rect 2514 223 2521 226
rect 2474 213 2493 216
rect 2490 206 2493 213
rect 2490 203 2501 206
rect 2498 163 2501 196
rect 2482 113 2485 136
rect 2506 123 2509 216
rect 2518 156 2521 223
rect 2538 216 2541 313
rect 2554 216 2557 423
rect 2578 423 2589 426
rect 2594 423 2605 426
rect 2618 423 2621 436
rect 2538 213 2549 216
rect 2554 213 2565 216
rect 2546 196 2549 213
rect 2530 193 2549 196
rect 2554 193 2557 206
rect 2562 166 2565 213
rect 2514 153 2521 156
rect 2554 163 2565 166
rect 2514 133 2517 153
rect 2554 143 2557 163
rect 2562 123 2565 156
rect 2578 113 2581 423
rect 2594 253 2597 423
rect 2626 413 2629 453
rect 2638 386 2641 533
rect 2638 383 2645 386
rect 2602 343 2605 366
rect 2618 333 2621 356
rect 2634 346 2637 366
rect 2626 343 2637 346
rect 2642 336 2645 383
rect 2650 346 2653 526
rect 2658 513 2661 526
rect 2674 473 2677 1256
rect 2658 423 2661 436
rect 2658 363 2661 406
rect 2650 343 2661 346
rect 2626 333 2645 336
rect 2626 323 2629 333
rect 2642 293 2645 326
rect 2658 286 2661 343
rect 2650 283 2661 286
rect 2586 223 2605 226
rect 2586 213 2589 223
rect 2594 203 2597 216
rect 2602 203 2605 223
rect 2610 213 2613 236
rect 2650 203 2653 283
rect 2594 133 2629 136
rect 2618 113 2621 126
rect 1618 83 1661 86
rect 1162 73 1189 76
rect 2686 37 2706 2503
rect 2710 13 2730 2527
<< metal3 >>
rect 1769 2452 2046 2457
rect 209 2442 294 2447
rect 1401 2442 1526 2447
rect 1769 2437 1774 2452
rect 2041 2437 2046 2452
rect 2089 2452 2214 2457
rect 2089 2437 2094 2452
rect 81 2432 166 2437
rect 241 2432 310 2437
rect 521 2432 654 2437
rect 1625 2432 1774 2437
rect 1841 2432 1926 2437
rect 2041 2432 2094 2437
rect 2209 2437 2214 2452
rect 2233 2442 2310 2447
rect 2329 2442 2398 2447
rect 2329 2437 2334 2442
rect 2209 2432 2334 2437
rect 2393 2437 2398 2442
rect 2441 2442 2638 2447
rect 2393 2432 2422 2437
rect 1841 2427 1846 2432
rect 1153 2422 1222 2427
rect 1785 2422 1846 2427
rect 1921 2427 1926 2432
rect 2441 2427 2446 2442
rect 1921 2422 2446 2427
rect 2633 2427 2638 2442
rect 2633 2422 2662 2427
rect 265 2412 302 2417
rect 673 2412 742 2417
rect 673 2407 678 2412
rect 633 2402 678 2407
rect 737 2407 742 2412
rect 1489 2412 1606 2417
rect 1857 2412 1910 2417
rect 2217 2412 2270 2417
rect 2289 2412 2318 2417
rect 737 2402 766 2407
rect 1257 2402 1374 2407
rect 1393 2402 1470 2407
rect 1257 2397 1262 2402
rect 97 2392 174 2397
rect 537 2392 1262 2397
rect 1369 2397 1374 2402
rect 1489 2397 1494 2412
rect 1369 2392 1494 2397
rect 1601 2397 1606 2412
rect 2289 2407 2294 2412
rect 1673 2402 1758 2407
rect 1809 2402 2294 2407
rect 2313 2407 2318 2412
rect 2457 2412 2622 2417
rect 2457 2407 2462 2412
rect 2313 2402 2462 2407
rect 2505 2402 2566 2407
rect 1601 2392 1630 2397
rect 2153 2392 2294 2397
rect 2537 2392 2638 2397
rect 1873 2387 2158 2392
rect 2289 2387 2294 2392
rect 521 2382 750 2387
rect 1377 2382 1446 2387
rect 649 2372 798 2377
rect 1273 2372 1358 2377
rect 1377 2367 1382 2382
rect 1441 2377 1446 2382
rect 1537 2382 1878 2387
rect 2177 2382 2270 2387
rect 2289 2382 2646 2387
rect 1537 2377 1542 2382
rect 1441 2372 1542 2377
rect 1569 2372 1710 2377
rect 1825 2372 1974 2377
rect 1993 2372 2062 2377
rect 1993 2367 1998 2372
rect 417 2362 670 2367
rect 1153 2362 1238 2367
rect 1313 2362 1382 2367
rect 1561 2362 1782 2367
rect 1945 2362 1998 2367
rect 2057 2367 2062 2372
rect 2057 2362 2254 2367
rect 1313 2357 1318 2362
rect 785 2352 870 2357
rect 1025 2352 1134 2357
rect 1025 2347 1030 2352
rect 497 2342 598 2347
rect 905 2342 1030 2347
rect 1129 2347 1134 2352
rect 1233 2352 1318 2357
rect 1329 2352 1422 2357
rect 1585 2352 1846 2357
rect 1937 2352 2046 2357
rect 1233 2347 1238 2352
rect 1129 2342 1238 2347
rect 1249 2342 1302 2347
rect 1321 2342 1446 2347
rect 1601 2342 1654 2347
rect 1665 2342 1750 2347
rect 1769 2342 1806 2347
rect 2065 2342 2222 2347
rect 2241 2342 2286 2347
rect 2305 2342 2374 2347
rect 2417 2342 2518 2347
rect 2577 2342 2654 2347
rect 1249 2337 1254 2342
rect 1649 2337 1654 2342
rect 1969 2337 2070 2342
rect 2217 2337 2222 2342
rect 2305 2337 2310 2342
rect 849 2332 918 2337
rect 969 2332 1038 2337
rect 1185 2332 1254 2337
rect 1265 2332 1398 2337
rect 1465 2332 1566 2337
rect 1649 2332 1974 2337
rect 2217 2332 2310 2337
rect 2369 2337 2374 2342
rect 2369 2332 2558 2337
rect 1185 2327 1190 2332
rect 1465 2327 1470 2332
rect 137 2322 190 2327
rect 361 2322 462 2327
rect 897 2322 950 2327
rect 1041 2322 1190 2327
rect 1209 2322 1470 2327
rect 1561 2327 1566 2332
rect 1561 2322 1710 2327
rect 1985 2322 2206 2327
rect 2297 2322 2390 2327
rect 1041 2317 1046 2322
rect 1705 2317 1990 2322
rect 2201 2317 2302 2322
rect 897 2312 1046 2317
rect 1057 2312 1534 2317
rect 1649 2312 1686 2317
rect 2009 2312 2110 2317
rect 2321 2312 2438 2317
rect 2561 2312 2598 2317
rect 329 2302 374 2307
rect 769 2302 1390 2307
rect 1481 2302 1574 2307
rect 1705 2302 1958 2307
rect 1977 2302 2086 2307
rect 2161 2302 2206 2307
rect 1705 2297 1710 2302
rect 833 2292 1390 2297
rect 1401 2292 1510 2297
rect 1521 2292 1598 2297
rect 1681 2292 1710 2297
rect 1953 2297 1958 2302
rect 2225 2297 2342 2302
rect 1953 2292 2230 2297
rect 2337 2292 2590 2297
rect 1657 2282 2102 2287
rect 953 2277 1086 2282
rect 1129 2277 1262 2282
rect 2097 2277 2102 2282
rect 2305 2282 2358 2287
rect 929 2272 958 2277
rect 1081 2272 1134 2277
rect 1257 2272 1342 2277
rect 1433 2272 1638 2277
rect 2097 2272 2198 2277
rect 417 2262 526 2267
rect 417 2257 422 2262
rect 89 2252 238 2257
rect 369 2252 422 2257
rect 521 2257 526 2262
rect 729 2262 886 2267
rect 729 2257 734 2262
rect 521 2252 734 2257
rect 881 2257 886 2262
rect 929 2257 934 2272
rect 1433 2267 1438 2272
rect 945 2262 982 2267
rect 1017 2262 1438 2267
rect 1633 2267 1638 2272
rect 1777 2267 1846 2272
rect 2193 2267 2198 2272
rect 2305 2267 2310 2282
rect 1633 2262 1782 2267
rect 1841 2262 2078 2267
rect 2193 2262 2310 2267
rect 2353 2267 2358 2282
rect 2545 2282 2574 2287
rect 2545 2267 2550 2282
rect 2353 2262 2550 2267
rect 881 2252 934 2257
rect 977 2257 982 2262
rect 1513 2257 1606 2262
rect 977 2252 1062 2257
rect 1345 2252 1518 2257
rect 1601 2252 1622 2257
rect 1793 2252 1830 2257
rect 2097 2252 2174 2257
rect 1057 2247 1350 2252
rect 1617 2247 1798 2252
rect 2001 2247 2102 2252
rect 2169 2247 2174 2252
rect 225 2242 510 2247
rect 785 2242 862 2247
rect 961 2242 1038 2247
rect 1473 2242 1590 2247
rect 1817 2242 1846 2247
rect 1905 2242 2006 2247
rect 2169 2242 2198 2247
rect 785 2237 790 2242
rect 857 2237 942 2242
rect 1369 2237 1454 2242
rect 1905 2237 1910 2242
rect 217 2232 382 2237
rect 745 2232 790 2237
rect 937 2232 1374 2237
rect 1449 2232 1910 2237
rect 1937 2232 2142 2237
rect 2217 2232 2318 2237
rect 2457 2232 2534 2237
rect 2593 2232 2630 2237
rect 2217 2227 2222 2232
rect 73 2222 118 2227
rect 177 2222 342 2227
rect 545 2222 646 2227
rect 801 2222 958 2227
rect 1089 2222 1118 2227
rect 1385 2222 1526 2227
rect 1881 2222 2038 2227
rect 2177 2222 2222 2227
rect 2313 2227 2318 2232
rect 2313 2222 2342 2227
rect 545 2217 550 2222
rect 953 2217 1094 2222
rect 1153 2217 1366 2222
rect 185 2212 230 2217
rect 241 2212 334 2217
rect 441 2212 550 2217
rect 1129 2212 1158 2217
rect 1361 2212 1462 2217
rect 1665 2212 1798 2217
rect 1841 2212 1966 2217
rect 2121 2212 2246 2217
rect 2305 2212 2510 2217
rect 2537 2212 2598 2217
rect 1665 2207 1670 2212
rect 377 2202 486 2207
rect 993 2202 1430 2207
rect 1449 2202 1670 2207
rect 1793 2207 1798 2212
rect 1793 2202 2046 2207
rect 81 2192 230 2197
rect 417 2192 518 2197
rect 889 2192 966 2197
rect 1145 2192 1182 2197
rect 1265 2192 1358 2197
rect 1457 2192 1902 2197
rect 2033 2192 2062 2197
rect 2225 2192 2270 2197
rect 2409 2192 2470 2197
rect 2489 2192 2534 2197
rect 1001 2182 1238 2187
rect 1265 2177 1270 2192
rect 1897 2187 2038 2192
rect 2465 2187 2470 2192
rect 1321 2182 1630 2187
rect 1705 2182 1878 2187
rect 2289 2182 2390 2187
rect 2465 2182 2606 2187
rect 2289 2177 2294 2182
rect 305 2172 398 2177
rect 1089 2172 1270 2177
rect 1345 2172 1446 2177
rect 1753 2172 1798 2177
rect 1969 2172 2038 2177
rect 2081 2172 2198 2177
rect 2217 2172 2294 2177
rect 2385 2177 2390 2182
rect 2385 2172 2622 2177
rect 305 2167 310 2172
rect 281 2162 310 2167
rect 393 2167 398 2172
rect 2081 2167 2086 2172
rect 393 2162 470 2167
rect 673 2162 734 2167
rect 1257 2162 1326 2167
rect 1353 2162 1542 2167
rect 1641 2162 2086 2167
rect 2193 2167 2198 2172
rect 2193 2162 2222 2167
rect 2305 2162 2398 2167
rect 2537 2162 2566 2167
rect 2217 2157 2310 2162
rect 2393 2157 2542 2162
rect 217 2152 390 2157
rect 953 2152 1078 2157
rect 1297 2152 1390 2157
rect 1873 2152 1974 2157
rect 1985 2152 2118 2157
rect 1297 2147 1302 2152
rect 1441 2147 1670 2152
rect 209 2142 294 2147
rect 505 2142 590 2147
rect 705 2142 830 2147
rect 1073 2142 1198 2147
rect 1233 2142 1302 2147
rect 1417 2142 1446 2147
rect 1665 2142 1694 2147
rect 1777 2142 1862 2147
rect 1977 2142 2334 2147
rect 2385 2142 2478 2147
rect 2537 2142 2614 2147
rect 505 2137 510 2142
rect 257 2132 510 2137
rect 585 2137 590 2142
rect 849 2137 974 2142
rect 1857 2137 1982 2142
rect 585 2132 614 2137
rect 721 2132 854 2137
rect 969 2132 998 2137
rect 1249 2132 1342 2137
rect 1393 2132 1670 2137
rect 2001 2132 2094 2137
rect 2177 2132 2254 2137
rect 161 2122 238 2127
rect 161 2117 166 2122
rect 233 2117 326 2122
rect 721 2117 726 2132
rect 745 2122 942 2127
rect 1017 2122 1110 2127
rect 1129 2122 1262 2127
rect 1017 2117 1022 2122
rect 113 2112 166 2117
rect 321 2112 350 2117
rect 521 2112 726 2117
rect 969 2112 1022 2117
rect 1105 2117 1110 2122
rect 1393 2117 1398 2132
rect 1569 2122 1614 2127
rect 1929 2122 2006 2127
rect 2249 2122 2342 2127
rect 2465 2122 2534 2127
rect 1569 2117 1574 2122
rect 2001 2117 2006 2122
rect 1105 2112 1398 2117
rect 1409 2112 1574 2117
rect 1593 2112 1614 2117
rect 1681 2112 1782 2117
rect 1801 2112 1910 2117
rect 2001 2112 2070 2117
rect 2489 2112 2550 2117
rect 2633 2112 2662 2117
rect 817 2107 950 2112
rect 1801 2107 1806 2112
rect 177 2102 270 2107
rect 329 2102 414 2107
rect 713 2102 782 2107
rect 793 2102 822 2107
rect 945 2102 1094 2107
rect 1273 2102 1358 2107
rect 1513 2102 1558 2107
rect 1769 2102 1806 2107
rect 1905 2107 1910 2112
rect 1905 2102 2166 2107
rect 1089 2097 1278 2102
rect 193 2092 310 2097
rect 345 2092 446 2097
rect 521 2092 694 2097
rect 825 2092 998 2097
rect 1297 2092 1374 2097
rect 1569 2092 1670 2097
rect 1689 2092 1998 2097
rect 521 2087 526 2092
rect 689 2087 782 2092
rect 1993 2087 1998 2092
rect 2097 2092 2126 2097
rect 2393 2092 2470 2097
rect 2097 2087 2102 2092
rect 2393 2087 2398 2092
rect 497 2082 526 2087
rect 777 2082 1094 2087
rect 1113 2082 1214 2087
rect 1393 2082 1494 2087
rect 1585 2082 1702 2087
rect 1801 2082 1918 2087
rect 1993 2082 2102 2087
rect 2369 2082 2398 2087
rect 2465 2087 2470 2092
rect 2465 2082 2510 2087
rect 1113 2077 1118 2082
rect 473 2072 702 2077
rect 737 2072 766 2077
rect 761 2067 766 2072
rect 857 2072 1118 2077
rect 1209 2077 1214 2082
rect 1313 2077 1398 2082
rect 1489 2077 1494 2082
rect 1209 2072 1318 2077
rect 1489 2072 1662 2077
rect 1761 2072 1974 2077
rect 2241 2072 2350 2077
rect 857 2067 862 2072
rect 2241 2067 2246 2072
rect 537 2062 638 2067
rect 761 2062 862 2067
rect 905 2062 1054 2067
rect 1161 2062 1198 2067
rect 1329 2062 1566 2067
rect 1857 2062 1982 2067
rect 2073 2062 2246 2067
rect 2345 2067 2350 2072
rect 2345 2062 2590 2067
rect 1049 2057 1142 2062
rect 1217 2057 1334 2062
rect 2073 2057 2078 2062
rect 137 2052 206 2057
rect 913 2052 1030 2057
rect 1137 2052 1222 2057
rect 1353 2052 1382 2057
rect 1529 2052 1766 2057
rect 1825 2052 1846 2057
rect 1929 2052 2078 2057
rect 2257 2052 2334 2057
rect 137 2047 142 2052
rect 81 2042 142 2047
rect 201 2047 206 2052
rect 1377 2047 1534 2052
rect 2329 2047 2334 2052
rect 2449 2052 2478 2057
rect 2449 2047 2454 2052
rect 201 2042 574 2047
rect 657 2042 734 2047
rect 881 2042 902 2047
rect 1049 2042 1334 2047
rect 1553 2042 1894 2047
rect 1961 2042 2014 2047
rect 2057 2042 2270 2047
rect 2329 2042 2454 2047
rect 153 2032 198 2037
rect 825 2032 910 2037
rect 929 2032 1030 2037
rect 1145 2032 1454 2037
rect 1505 2032 1534 2037
rect 929 2027 934 2032
rect 1025 2027 1126 2032
rect 1553 2027 1558 2042
rect 1577 2032 1606 2037
rect 633 2022 678 2027
rect 849 2022 934 2027
rect 1121 2022 1558 2027
rect 1601 2027 1606 2032
rect 1689 2032 1798 2037
rect 1897 2032 1998 2037
rect 2073 2032 2134 2037
rect 2169 2032 2286 2037
rect 1689 2027 1694 2032
rect 1601 2022 1694 2027
rect 1713 2022 1758 2027
rect 1817 2022 1878 2027
rect 1905 2022 1982 2027
rect 2001 2022 2094 2027
rect 2113 2022 2454 2027
rect 185 2012 350 2017
rect 609 2012 758 2017
rect 849 2007 854 2022
rect 2001 2017 2006 2022
rect 865 2012 934 2017
rect 945 2012 1014 2017
rect 1033 2012 1166 2017
rect 1185 2012 1270 2017
rect 1393 2012 1462 2017
rect 1881 2012 2006 2017
rect 2177 2012 2318 2017
rect 393 2002 494 2007
rect 625 2002 854 2007
rect 1009 2007 1014 2012
rect 1665 2007 1862 2012
rect 2025 2007 2094 2012
rect 1009 2002 1062 2007
rect 1521 2002 1670 2007
rect 1857 2002 1910 2007
rect 1969 2002 2030 2007
rect 2089 2002 2270 2007
rect 393 1997 398 2002
rect 201 1992 262 1997
rect 369 1992 398 1997
rect 489 1997 494 2002
rect 1057 1997 1062 2002
rect 1217 1997 1318 2002
rect 1521 1997 1526 2002
rect 489 1992 518 1997
rect 633 1992 670 1997
rect 689 1992 822 1997
rect 889 1992 950 1997
rect 1009 1992 1038 1997
rect 1057 1992 1222 1997
rect 1313 1992 1446 1997
rect 1473 1992 1526 1997
rect 1537 1992 1590 1997
rect 1681 1992 1814 1997
rect 1841 1992 2078 1997
rect 2113 1987 2198 1992
rect 73 1982 494 1987
rect 529 1982 654 1987
rect 953 1982 1094 1987
rect 1233 1982 1358 1987
rect 1465 1982 1574 1987
rect 1657 1982 1750 1987
rect 1905 1982 2014 1987
rect 2089 1982 2118 1987
rect 2193 1982 2222 1987
rect 2329 1982 2478 1987
rect 2537 1982 2606 1987
rect 1113 1977 1214 1982
rect 1769 1977 1886 1982
rect 2009 1977 2094 1982
rect 2329 1977 2334 1982
rect 377 1972 486 1977
rect 657 1972 742 1977
rect 921 1972 1118 1977
rect 1209 1972 1678 1977
rect 1729 1972 1774 1977
rect 1881 1972 1926 1977
rect 1945 1972 1990 1977
rect 2129 1972 2158 1977
rect 2153 1967 2158 1972
rect 2233 1972 2334 1977
rect 2473 1977 2478 1982
rect 2473 1972 2510 1977
rect 2233 1967 2238 1972
rect 673 1962 742 1967
rect 1001 1962 1350 1967
rect 1425 1962 2102 1967
rect 2153 1962 2238 1967
rect 1425 1957 1430 1962
rect 185 1952 270 1957
rect 857 1952 1262 1957
rect 1361 1952 1430 1957
rect 1449 1952 1702 1957
rect 1793 1952 1822 1957
rect 1865 1952 2110 1957
rect 2345 1952 2390 1957
rect 2417 1952 2462 1957
rect 721 1947 838 1952
rect 1257 1947 1366 1952
rect 1697 1947 1782 1952
rect 2417 1947 2422 1952
rect 145 1942 222 1947
rect 465 1942 566 1947
rect 697 1942 726 1947
rect 833 1942 1166 1947
rect 1409 1942 1510 1947
rect 1777 1942 2022 1947
rect 2033 1942 2334 1947
rect 2393 1942 2422 1947
rect 2433 1942 2510 1947
rect 2577 1942 2678 1947
rect 1529 1937 1670 1942
rect 2033 1937 2038 1942
rect 2329 1937 2398 1942
rect 401 1932 430 1937
rect 513 1932 542 1937
rect 641 1932 1006 1937
rect 1113 1932 1294 1937
rect 1377 1932 1534 1937
rect 1665 1932 2038 1937
rect 2553 1932 2590 1937
rect 425 1927 518 1932
rect 2057 1927 2230 1932
rect 145 1922 182 1927
rect 545 1922 630 1927
rect 777 1922 918 1927
rect 1009 1922 1070 1927
rect 1137 1922 1318 1927
rect 1337 1922 1414 1927
rect 1473 1922 1654 1927
rect 1737 1922 2062 1927
rect 2225 1922 2470 1927
rect 201 1912 238 1917
rect 393 1912 494 1917
rect 393 1907 398 1912
rect 169 1902 286 1907
rect 369 1902 398 1907
rect 489 1907 494 1912
rect 545 1907 550 1922
rect 625 1917 782 1922
rect 801 1912 878 1917
rect 1001 1912 1158 1917
rect 1209 1912 1294 1917
rect 1401 1912 1430 1917
rect 1513 1912 1582 1917
rect 1801 1912 1854 1917
rect 1897 1912 2078 1917
rect 2089 1912 2174 1917
rect 2185 1912 2214 1917
rect 2209 1907 2214 1912
rect 2417 1912 2446 1917
rect 2417 1907 2422 1912
rect 489 1902 550 1907
rect 649 1902 822 1907
rect 841 1902 886 1907
rect 1089 1902 1494 1907
rect 1513 1902 1574 1907
rect 1601 1902 1678 1907
rect 2033 1902 2102 1907
rect 2209 1902 2422 1907
rect 817 1897 822 1902
rect 905 1897 1070 1902
rect 1601 1897 1606 1902
rect 393 1892 670 1897
rect 817 1892 910 1897
rect 1065 1892 1430 1897
rect 1561 1892 1606 1897
rect 1673 1897 1678 1902
rect 1673 1892 1702 1897
rect 1721 1892 2014 1897
rect 305 1887 398 1892
rect 689 1887 798 1892
rect 1449 1887 1542 1892
rect 1721 1887 1726 1892
rect 2009 1887 2086 1892
rect 73 1882 294 1887
rect 89 1872 118 1877
rect 113 1857 118 1872
rect 305 1857 310 1887
rect 417 1882 694 1887
rect 793 1882 1110 1887
rect 1257 1882 1342 1887
rect 1417 1882 1454 1887
rect 1537 1882 1726 1887
rect 2081 1882 2510 1887
rect 1105 1877 1262 1882
rect 1745 1877 1990 1882
rect 433 1872 814 1877
rect 809 1867 814 1872
rect 905 1872 990 1877
rect 1049 1872 1086 1877
rect 1281 1872 1606 1877
rect 1641 1872 1750 1877
rect 1985 1872 2070 1877
rect 905 1867 910 1872
rect 1281 1867 1286 1872
rect 2169 1867 2270 1872
rect 561 1862 790 1867
rect 809 1862 910 1867
rect 929 1862 1286 1867
rect 1305 1862 1902 1867
rect 1913 1862 2014 1867
rect 2145 1862 2174 1867
rect 2265 1862 2294 1867
rect 2321 1862 2358 1867
rect 2377 1862 2446 1867
rect 2145 1857 2150 1862
rect 2377 1857 2382 1862
rect 113 1852 310 1857
rect 545 1852 646 1857
rect 657 1852 686 1857
rect 1241 1852 1550 1857
rect 1577 1852 1694 1857
rect 1761 1852 1798 1857
rect 1961 1852 2150 1857
rect 2161 1852 2382 1857
rect 2441 1857 2446 1862
rect 2441 1852 2582 1857
rect 873 1847 1022 1852
rect 369 1842 470 1847
rect 537 1842 702 1847
rect 849 1842 878 1847
rect 1017 1842 1174 1847
rect 1217 1842 1406 1847
rect 1545 1842 2038 1847
rect 2049 1842 2102 1847
rect 2249 1842 2430 1847
rect 369 1837 374 1842
rect 345 1832 374 1837
rect 465 1837 470 1842
rect 1217 1837 1222 1842
rect 1401 1837 1550 1842
rect 465 1832 494 1837
rect 529 1832 686 1837
rect 833 1832 1222 1837
rect 1233 1832 1382 1837
rect 1569 1832 1638 1837
rect 1713 1832 2358 1837
rect 1569 1827 1574 1832
rect 2353 1827 2358 1832
rect 2441 1832 2542 1837
rect 2441 1827 2446 1832
rect 289 1822 318 1827
rect 385 1822 486 1827
rect 521 1822 582 1827
rect 881 1822 926 1827
rect 985 1822 1022 1827
rect 1137 1822 1214 1827
rect 1249 1822 1310 1827
rect 1329 1822 1398 1827
rect 1425 1822 1574 1827
rect 1585 1822 1750 1827
rect 1761 1822 1934 1827
rect 313 1817 390 1822
rect 1425 1817 1430 1822
rect 585 1812 646 1817
rect 713 1812 1430 1817
rect 1441 1812 1574 1817
rect 1713 1807 1718 1817
rect 537 1802 694 1807
rect 737 1802 846 1807
rect 865 1802 1206 1807
rect 1217 1802 1270 1807
rect 1385 1802 1718 1807
rect 1745 1807 1750 1822
rect 1953 1817 1958 1827
rect 1985 1822 2190 1827
rect 2305 1822 2334 1827
rect 2353 1822 2446 1827
rect 1873 1812 1958 1817
rect 2017 1812 2158 1817
rect 1953 1807 1958 1812
rect 1745 1802 1910 1807
rect 1953 1802 2206 1807
rect 2297 1802 2398 1807
rect 2417 1802 2486 1807
rect 2417 1797 2422 1802
rect 121 1792 478 1797
rect 529 1792 614 1797
rect 761 1792 934 1797
rect 961 1792 1302 1797
rect 1353 1792 1406 1797
rect 1449 1792 1550 1797
rect 1609 1792 1670 1797
rect 1713 1792 1758 1797
rect 1897 1792 2006 1797
rect 2065 1792 2142 1797
rect 2353 1792 2422 1797
rect 2481 1797 2486 1802
rect 2481 1792 2542 1797
rect 2553 1792 2678 1797
rect 2353 1787 2358 1792
rect 673 1782 838 1787
rect 905 1782 974 1787
rect 1025 1782 1350 1787
rect 1377 1782 1398 1787
rect 1409 1782 1478 1787
rect 1905 1782 2126 1787
rect 2225 1782 2358 1787
rect 2377 1782 2470 1787
rect 769 1772 854 1777
rect 929 1772 2054 1777
rect 2361 1772 2390 1777
rect 617 1762 806 1767
rect 1049 1762 1502 1767
rect 1905 1762 2182 1767
rect 801 1757 1014 1762
rect 1521 1757 1630 1762
rect 73 1752 430 1757
rect 1009 1752 1038 1757
rect 1129 1752 1166 1757
rect 1177 1752 1238 1757
rect 1249 1752 1526 1757
rect 1625 1752 1654 1757
rect 1673 1752 1750 1757
rect 1849 1752 1894 1757
rect 1673 1747 1678 1752
rect 177 1742 294 1747
rect 729 1742 782 1747
rect 849 1742 1678 1747
rect 1745 1747 1750 1752
rect 1745 1742 1774 1747
rect 1905 1737 1910 1762
rect 1961 1752 2150 1757
rect 2289 1752 2478 1757
rect 2521 1752 2582 1757
rect 2289 1747 2294 1752
rect 1985 1742 2062 1747
rect 2089 1742 2182 1747
rect 2209 1742 2294 1747
rect 2489 1742 2518 1747
rect 2177 1737 2182 1742
rect 2513 1737 2518 1742
rect 2593 1742 2646 1747
rect 2593 1737 2598 1742
rect 729 1732 950 1737
rect 977 1732 1126 1737
rect 1137 1732 1254 1737
rect 1265 1732 1390 1737
rect 1497 1732 1558 1737
rect 1617 1732 1910 1737
rect 1921 1732 2158 1737
rect 2177 1732 2246 1737
rect 2265 1732 2318 1737
rect 2345 1732 2478 1737
rect 2513 1732 2598 1737
rect 2633 1732 2678 1737
rect 697 1722 886 1727
rect 1105 1722 1134 1727
rect 1185 1722 1214 1727
rect 1377 1722 2374 1727
rect 961 1717 1086 1722
rect 1281 1717 1382 1722
rect 185 1712 278 1717
rect 561 1712 662 1717
rect 937 1712 966 1717
rect 1081 1712 1262 1717
rect 1281 1707 1286 1717
rect 1401 1712 1654 1717
rect 1745 1712 2286 1717
rect 2321 1712 2358 1717
rect 137 1702 222 1707
rect 537 1702 574 1707
rect 641 1702 742 1707
rect 761 1702 814 1707
rect 881 1702 1102 1707
rect 1145 1702 1246 1707
rect 1257 1702 1286 1707
rect 1313 1702 1606 1707
rect 1865 1702 1990 1707
rect 2009 1702 2446 1707
rect 1745 1697 1846 1702
rect 201 1692 230 1697
rect 225 1687 230 1692
rect 289 1692 366 1697
rect 841 1692 878 1697
rect 289 1687 294 1692
rect 225 1682 294 1687
rect 873 1687 878 1692
rect 937 1692 1118 1697
rect 1289 1692 1470 1697
rect 1553 1692 1702 1697
rect 1721 1692 1750 1697
rect 1841 1692 1862 1697
rect 1961 1692 2086 1697
rect 2105 1692 2334 1697
rect 2385 1692 2454 1697
rect 937 1687 942 1692
rect 1137 1687 1270 1692
rect 1857 1687 1966 1692
rect 873 1682 942 1687
rect 1089 1682 1142 1687
rect 1265 1682 1670 1687
rect 1769 1682 1838 1687
rect 1985 1682 2030 1687
rect 2097 1682 2142 1687
rect 2241 1682 2558 1687
rect 721 1672 854 1677
rect 1073 1672 1782 1677
rect 1937 1672 2398 1677
rect 2537 1672 2566 1677
rect 1937 1667 1942 1672
rect 2393 1667 2542 1672
rect 753 1662 806 1667
rect 1297 1662 1406 1667
rect 1441 1662 1622 1667
rect 1665 1662 1686 1667
rect 1705 1662 1942 1667
rect 1953 1662 2126 1667
rect 2161 1662 2374 1667
rect 1017 1657 1182 1662
rect 1681 1657 1686 1662
rect 2161 1657 2166 1662
rect 873 1652 974 1657
rect 993 1652 1022 1657
rect 1177 1652 1662 1657
rect 1681 1652 1726 1657
rect 1737 1652 1870 1657
rect 1969 1652 2110 1657
rect 2121 1652 2166 1657
rect 2185 1652 2238 1657
rect 2393 1652 2510 1657
rect 873 1647 878 1652
rect 849 1642 878 1647
rect 969 1647 974 1652
rect 2257 1647 2398 1652
rect 2505 1647 2510 1652
rect 969 1642 1166 1647
rect 1345 1642 1422 1647
rect 1505 1642 1574 1647
rect 1689 1642 1758 1647
rect 1913 1642 1982 1647
rect 2137 1642 2262 1647
rect 2505 1642 2534 1647
rect 1777 1637 1886 1642
rect 2033 1637 2142 1642
rect 201 1632 278 1637
rect 601 1632 630 1637
rect 1009 1632 1494 1637
rect 1585 1632 1782 1637
rect 1881 1632 1910 1637
rect 2033 1632 2038 1637
rect 2161 1632 2526 1637
rect 1489 1627 1590 1632
rect 1929 1627 2038 1632
rect 129 1622 222 1627
rect 417 1622 518 1627
rect 593 1622 654 1627
rect 721 1622 774 1627
rect 865 1622 974 1627
rect 1337 1622 1470 1627
rect 1649 1622 1934 1627
rect 2049 1622 2198 1627
rect 2297 1622 2470 1627
rect 2481 1622 2518 1627
rect 2537 1622 2670 1627
rect 241 1612 350 1617
rect 241 1607 246 1612
rect 217 1602 246 1607
rect 345 1607 350 1612
rect 401 1607 406 1617
rect 345 1602 406 1607
rect 129 1592 334 1597
rect 417 1592 422 1622
rect 993 1617 1246 1622
rect 2193 1617 2302 1622
rect 497 1612 686 1617
rect 889 1612 998 1617
rect 1241 1612 1302 1617
rect 1361 1612 1438 1617
rect 1521 1612 1758 1617
rect 1785 1612 1822 1617
rect 1913 1612 2174 1617
rect 2321 1607 2398 1612
rect 2465 1607 2470 1622
rect 489 1602 558 1607
rect 657 1602 718 1607
rect 793 1602 862 1607
rect 969 1602 998 1607
rect 1009 1602 1230 1607
rect 1377 1602 1662 1607
rect 1961 1602 2086 1607
rect 2105 1602 2326 1607
rect 2393 1602 2422 1607
rect 2465 1602 2494 1607
rect 2633 1602 2670 1607
rect 857 1597 974 1602
rect 1225 1597 1382 1602
rect 1681 1597 1750 1602
rect 2081 1597 2086 1602
rect 497 1592 534 1597
rect 1073 1592 1206 1597
rect 1401 1592 1454 1597
rect 1497 1592 1686 1597
rect 1745 1592 1926 1597
rect 2081 1592 2182 1597
rect 2337 1592 2454 1597
rect 265 1582 310 1587
rect 385 1582 582 1587
rect 697 1582 774 1587
rect 809 1582 838 1587
rect 937 1582 1030 1587
rect 1305 1582 1734 1587
rect 1873 1582 1966 1587
rect 2033 1582 2190 1587
rect 2281 1582 2358 1587
rect 2497 1582 2582 1587
rect 305 1577 310 1582
rect 577 1577 582 1582
rect 937 1577 942 1582
rect 1025 1577 1286 1582
rect 1873 1577 1878 1582
rect 2377 1577 2478 1582
rect 305 1572 454 1577
rect 577 1572 646 1577
rect 721 1572 782 1577
rect 849 1572 942 1577
rect 1281 1572 1878 1577
rect 1897 1572 2166 1577
rect 2201 1572 2382 1577
rect 2473 1572 2518 1577
rect 777 1567 854 1572
rect 953 1562 1014 1567
rect 1081 1562 1934 1567
rect 1985 1562 2134 1567
rect 2265 1562 2438 1567
rect 2457 1562 2510 1567
rect 593 1557 758 1562
rect 513 1552 598 1557
rect 753 1552 782 1557
rect 801 1552 870 1557
rect 913 1552 1030 1557
rect 1145 1552 1574 1557
rect 1609 1552 1646 1557
rect 1969 1552 2126 1557
rect 801 1547 806 1552
rect 209 1527 214 1547
rect 609 1542 678 1547
rect 705 1542 742 1547
rect 761 1542 806 1547
rect 865 1547 870 1552
rect 1025 1547 1126 1552
rect 1737 1547 1822 1552
rect 2289 1547 2294 1557
rect 2369 1552 2486 1557
rect 865 1542 894 1547
rect 1121 1542 1166 1547
rect 1217 1542 1534 1547
rect 1577 1542 1638 1547
rect 1713 1542 1742 1547
rect 1817 1542 1990 1547
rect 2081 1542 2238 1547
rect 2273 1542 2294 1547
rect 2305 1542 2326 1547
rect 2441 1542 2510 1547
rect 2521 1542 2646 1547
rect 473 1537 574 1542
rect 2273 1537 2278 1542
rect 449 1532 478 1537
rect 569 1532 598 1537
rect 593 1527 598 1532
rect 665 1532 958 1537
rect 1089 1532 1198 1537
rect 1273 1532 1318 1537
rect 1385 1532 1454 1537
rect 1521 1532 1590 1537
rect 1617 1532 1750 1537
rect 1769 1532 1806 1537
rect 2001 1532 2022 1537
rect 2145 1532 2302 1537
rect 2313 1532 2438 1537
rect 665 1527 670 1532
rect 977 1527 1070 1532
rect 193 1522 214 1527
rect 497 1522 542 1527
rect 593 1522 670 1527
rect 689 1522 774 1527
rect 857 1522 982 1527
rect 1065 1522 1998 1527
rect 2017 1517 2022 1532
rect 2057 1522 2550 1527
rect 729 1512 1078 1517
rect 1089 1512 1502 1517
rect 1593 1512 2006 1517
rect 2017 1512 2070 1517
rect 2001 1507 2006 1512
rect 2137 1507 2142 1517
rect 2169 1512 2382 1517
rect 2417 1512 2470 1517
rect 217 1502 998 1507
rect 1065 1502 1230 1507
rect 1345 1502 1374 1507
rect 1409 1502 1742 1507
rect 1777 1502 1910 1507
rect 2001 1502 2118 1507
rect 2137 1502 2230 1507
rect 2241 1502 2270 1507
rect 2281 1502 2542 1507
rect 705 1492 918 1497
rect 937 1492 1062 1497
rect 1145 1492 1214 1497
rect 1265 1492 1654 1497
rect 1801 1492 2102 1497
rect 2161 1492 2190 1497
rect 913 1487 918 1492
rect 2185 1487 2190 1492
rect 2369 1492 2398 1497
rect 2369 1487 2374 1492
rect 473 1482 862 1487
rect 913 1482 1006 1487
rect 1169 1482 1710 1487
rect 1769 1482 2150 1487
rect 2185 1482 2374 1487
rect 657 1472 1038 1477
rect 1097 1472 1854 1477
rect 1953 1467 2030 1472
rect 2097 1467 2198 1472
rect 337 1462 742 1467
rect 977 1462 1350 1467
rect 1425 1462 1566 1467
rect 1617 1462 1694 1467
rect 1753 1462 1958 1467
rect 2025 1462 2102 1467
rect 2193 1462 2222 1467
rect 2241 1462 2382 1467
rect 737 1457 982 1462
rect 2241 1457 2246 1462
rect 249 1452 374 1457
rect 577 1452 606 1457
rect 689 1452 718 1457
rect 1001 1452 1558 1457
rect 1569 1452 1806 1457
rect 1969 1452 2014 1457
rect 2113 1452 2246 1457
rect 2377 1457 2382 1462
rect 2377 1452 2406 1457
rect 601 1447 694 1452
rect 1553 1447 1558 1452
rect 1969 1447 1974 1452
rect 809 1442 1014 1447
rect 1105 1442 1278 1447
rect 1345 1442 1390 1447
rect 1425 1442 1462 1447
rect 1473 1442 1526 1447
rect 1553 1442 1582 1447
rect 1633 1442 1846 1447
rect 1889 1442 1974 1447
rect 1985 1442 2062 1447
rect 2089 1442 2566 1447
rect 1633 1437 1638 1442
rect 305 1432 526 1437
rect 617 1432 862 1437
rect 1073 1432 1398 1437
rect 1529 1432 1638 1437
rect 1713 1432 2006 1437
rect 2017 1432 2230 1437
rect 2401 1432 2454 1437
rect 305 1427 310 1432
rect 209 1422 310 1427
rect 521 1427 526 1432
rect 2001 1427 2006 1432
rect 521 1422 550 1427
rect 769 1422 814 1427
rect 825 1422 910 1427
rect 1049 1422 1086 1427
rect 1137 1417 1142 1427
rect 1161 1422 1262 1427
rect 1297 1422 1334 1427
rect 1361 1422 1614 1427
rect 1721 1422 1774 1427
rect 1889 1422 1966 1427
rect 2001 1422 2358 1427
rect 2393 1422 2470 1427
rect 2553 1422 2614 1427
rect 321 1412 454 1417
rect 633 1412 1142 1417
rect 1201 1412 1974 1417
rect 2113 1407 2118 1417
rect 2185 1412 2214 1417
rect 2249 1412 2302 1417
rect 2377 1412 2438 1417
rect 2529 1412 2622 1417
rect 321 1402 358 1407
rect 441 1402 862 1407
rect 1041 1402 1102 1407
rect 1281 1402 1558 1407
rect 1649 1402 1766 1407
rect 1777 1402 2118 1407
rect 2281 1402 2310 1407
rect 2321 1402 2486 1407
rect 2545 1402 2662 1407
rect 353 1397 358 1402
rect 129 1392 174 1397
rect 297 1392 334 1397
rect 353 1392 526 1397
rect 609 1392 654 1397
rect 737 1392 982 1397
rect 993 1392 1086 1397
rect 1193 1392 1430 1397
rect 1465 1392 1638 1397
rect 1841 1392 1990 1397
rect 2041 1392 2470 1397
rect 2553 1392 2582 1397
rect 609 1387 614 1392
rect 2577 1387 2582 1392
rect 2641 1392 2670 1397
rect 2641 1387 2646 1392
rect 81 1382 134 1387
rect 337 1382 614 1387
rect 641 1382 726 1387
rect 753 1382 806 1387
rect 841 1382 1030 1387
rect 1249 1382 1622 1387
rect 1745 1382 2062 1387
rect 2185 1382 2214 1387
rect 2409 1382 2438 1387
rect 2577 1382 2646 1387
rect 1049 1377 1158 1382
rect 2209 1377 2414 1382
rect 81 1372 454 1377
rect 577 1372 1054 1377
rect 1153 1372 1302 1377
rect 1425 1372 1726 1377
rect 1897 1372 1966 1377
rect 2025 1372 2134 1377
rect 2449 1372 2534 1377
rect 1297 1367 1430 1372
rect 169 1362 198 1367
rect 321 1362 822 1367
rect 841 1362 886 1367
rect 1001 1362 1142 1367
rect 1209 1362 1278 1367
rect 1449 1362 1518 1367
rect 1561 1362 1934 1367
rect 2113 1362 2286 1367
rect 193 1357 326 1362
rect 345 1352 542 1357
rect 585 1352 726 1357
rect 817 1347 822 1362
rect 2281 1357 2286 1362
rect 2361 1362 2478 1367
rect 2361 1357 2366 1362
rect 849 1352 942 1357
rect 953 1352 1054 1357
rect 1081 1352 1134 1357
rect 1257 1352 1326 1357
rect 1385 1352 1670 1357
rect 1737 1352 1790 1357
rect 1881 1352 2038 1357
rect 2057 1352 2094 1357
rect 2281 1352 2366 1357
rect 113 1342 230 1347
rect 521 1342 574 1347
rect 649 1342 718 1347
rect 769 1342 798 1347
rect 817 1342 894 1347
rect 945 1342 1366 1347
rect 1393 1342 1574 1347
rect 1617 1342 1702 1347
rect 1889 1342 1942 1347
rect 1953 1342 2182 1347
rect 2201 1342 2262 1347
rect 345 1337 502 1342
rect 1617 1337 1622 1342
rect 1721 1337 1870 1342
rect 1953 1337 1958 1342
rect 2177 1337 2182 1342
rect 201 1332 254 1337
rect 321 1332 350 1337
rect 497 1332 686 1337
rect 937 1332 966 1337
rect 1057 1332 1622 1337
rect 1673 1332 1726 1337
rect 1865 1332 1958 1337
rect 1985 1332 2142 1337
rect 2177 1332 2222 1337
rect 1057 1327 1062 1332
rect 289 1322 422 1327
rect 441 1322 502 1327
rect 641 1322 694 1327
rect 705 1322 1062 1327
rect 1073 1322 1342 1327
rect 1425 1322 1550 1327
rect 1561 1322 1614 1327
rect 1657 1322 1758 1327
rect 1769 1322 2350 1327
rect 2609 1322 2670 1327
rect 417 1317 422 1322
rect 705 1317 710 1322
rect 1073 1317 1078 1322
rect 313 1312 390 1317
rect 417 1312 446 1317
rect 481 1312 662 1317
rect 689 1312 710 1317
rect 889 1312 1078 1317
rect 1113 1312 1806 1317
rect 1833 1312 1894 1317
rect 1937 1312 2238 1317
rect 393 1302 414 1307
rect 457 1302 518 1307
rect 833 1302 1822 1307
rect 1881 1302 1966 1307
rect 1977 1302 2086 1307
rect 545 1297 814 1302
rect 521 1292 550 1297
rect 809 1292 1062 1297
rect 1289 1292 1350 1297
rect 1417 1292 1438 1297
rect 1457 1292 1646 1297
rect 1761 1292 1990 1297
rect 2009 1292 2062 1297
rect 2105 1292 2134 1297
rect 2217 1292 2334 1297
rect 1081 1287 1270 1292
rect 1641 1287 1766 1292
rect 409 1282 1086 1287
rect 1265 1282 1318 1287
rect 1337 1282 1470 1287
rect 1577 1282 1622 1287
rect 1785 1282 1814 1287
rect 1929 1282 1958 1287
rect 2017 1282 2158 1287
rect 2169 1282 2326 1287
rect 2353 1282 2518 1287
rect 1809 1277 1934 1282
rect 449 1272 526 1277
rect 633 1272 662 1277
rect 761 1272 1230 1277
rect 1249 1272 1342 1277
rect 1425 1272 1686 1277
rect 2009 1272 2278 1277
rect 657 1267 766 1272
rect 1425 1267 1430 1272
rect 2353 1267 2358 1282
rect 257 1262 478 1267
rect 785 1262 854 1267
rect 873 1262 1430 1267
rect 1449 1262 1598 1267
rect 1609 1262 1782 1267
rect 1793 1262 1854 1267
rect 1921 1262 1998 1267
rect 2137 1262 2358 1267
rect 2513 1267 2518 1282
rect 2513 1262 2542 1267
rect 1777 1257 1782 1262
rect 2017 1257 2118 1262
rect 417 1252 774 1257
rect 1089 1252 1142 1257
rect 1233 1252 1766 1257
rect 1777 1252 2022 1257
rect 2113 1252 2678 1257
rect 769 1247 1078 1252
rect 1137 1247 1238 1252
rect 345 1242 462 1247
rect 457 1237 462 1242
rect 537 1242 566 1247
rect 1073 1242 1118 1247
rect 1257 1242 1398 1247
rect 1417 1242 1630 1247
rect 1721 1242 2054 1247
rect 2065 1242 2174 1247
rect 2185 1242 2334 1247
rect 537 1237 542 1242
rect 1625 1237 1726 1242
rect 2065 1237 2070 1242
rect 2433 1237 2518 1242
rect 353 1232 438 1237
rect 457 1232 542 1237
rect 697 1232 814 1237
rect 849 1232 958 1237
rect 1033 1232 1230 1237
rect 1273 1232 1606 1237
rect 1745 1232 1918 1237
rect 1945 1232 2006 1237
rect 2041 1232 2070 1237
rect 2161 1232 2206 1237
rect 2241 1232 2438 1237
rect 2513 1232 2542 1237
rect 113 1222 230 1227
rect 641 1222 678 1227
rect 969 1222 1422 1227
rect 1433 1222 1510 1227
rect 1553 1222 2350 1227
rect 2449 1222 2486 1227
rect 2561 1222 2614 1227
rect 273 1217 358 1222
rect 201 1212 278 1217
rect 353 1212 382 1217
rect 409 1212 510 1217
rect 521 1212 574 1217
rect 641 1207 646 1222
rect 673 1212 918 1217
rect 961 1212 1102 1217
rect 1113 1212 1518 1217
rect 1665 1212 1806 1217
rect 1905 1212 2422 1217
rect 1537 1207 1646 1212
rect 289 1202 342 1207
rect 569 1202 598 1207
rect 617 1202 646 1207
rect 1209 1202 1542 1207
rect 1641 1202 2462 1207
rect 825 1197 910 1202
rect 985 1197 1190 1202
rect 273 1192 462 1197
rect 657 1192 830 1197
rect 905 1192 990 1197
rect 1185 1192 1222 1197
rect 1377 1192 1686 1197
rect 1705 1192 2342 1197
rect 2361 1192 2406 1197
rect 2417 1192 2446 1197
rect 2465 1192 2534 1197
rect 1233 1187 1382 1192
rect 265 1182 486 1187
rect 553 1182 718 1187
rect 801 1182 894 1187
rect 1001 1182 1054 1187
rect 1097 1182 1150 1187
rect 1193 1182 1238 1187
rect 1401 1182 1494 1187
rect 1537 1182 1990 1187
rect 2017 1182 2070 1187
rect 2281 1182 2318 1187
rect 889 1177 1006 1182
rect 2169 1177 2262 1182
rect 201 1172 254 1177
rect 337 1172 390 1177
rect 513 1172 566 1177
rect 745 1172 870 1177
rect 1025 1172 1110 1177
rect 1129 1172 1286 1177
rect 1313 1172 1430 1177
rect 1473 1172 1798 1177
rect 1825 1172 1862 1177
rect 1961 1172 2030 1177
rect 2145 1172 2174 1177
rect 2257 1172 2374 1177
rect 217 1162 334 1167
rect 441 1162 630 1167
rect 761 1162 1030 1167
rect 1089 1162 1414 1167
rect 1481 1162 2334 1167
rect 2465 1162 2590 1167
rect 1025 1157 1030 1162
rect 81 1152 214 1157
rect 249 1152 326 1157
rect 457 1152 534 1157
rect 545 1152 1014 1157
rect 1025 1152 1134 1157
rect 1225 1152 1254 1157
rect 1337 1152 1526 1157
rect 1577 1152 1878 1157
rect 2009 1152 2118 1157
rect 2169 1152 2478 1157
rect 1009 1147 1014 1152
rect 1249 1147 1342 1152
rect 193 1142 286 1147
rect 361 1142 390 1147
rect 417 1142 470 1147
rect 545 1142 662 1147
rect 769 1142 966 1147
rect 1009 1142 1214 1147
rect 1441 1142 1998 1147
rect 2065 1142 2206 1147
rect 2313 1142 2350 1147
rect 2521 1142 2598 1147
rect 2609 1142 2638 1147
rect 681 1137 774 1142
rect 1209 1137 1214 1142
rect 1361 1137 1446 1142
rect 1993 1137 2070 1142
rect 489 1132 582 1137
rect 601 1132 686 1137
rect 785 1132 870 1137
rect 953 1132 1070 1137
rect 1209 1132 1366 1137
rect 1465 1132 1590 1137
rect 1641 1132 1774 1137
rect 1801 1132 1846 1137
rect 2089 1132 2630 1137
rect 305 1122 822 1127
rect 945 1122 998 1127
rect 1105 1122 1166 1127
rect 1385 1122 1558 1127
rect 1633 1122 1958 1127
rect 1985 1122 2230 1127
rect 2289 1122 2406 1127
rect 2289 1117 2294 1122
rect 129 1112 198 1117
rect 561 1112 686 1117
rect 801 1112 830 1117
rect 849 1112 958 1117
rect 1017 1112 1366 1117
rect 1425 1112 1990 1117
rect 2025 1112 2086 1117
rect 2137 1112 2166 1117
rect 2265 1112 2294 1117
rect 2361 1112 2430 1117
rect 2449 1112 2526 1117
rect 681 1107 806 1112
rect 1361 1107 1366 1112
rect 2161 1107 2270 1112
rect 2289 1107 2294 1112
rect 2449 1107 2454 1112
rect 113 1102 142 1107
rect 281 1102 382 1107
rect 449 1102 662 1107
rect 841 1102 1174 1107
rect 1185 1102 1230 1107
rect 1361 1102 1486 1107
rect 1545 1102 1638 1107
rect 1681 1102 2126 1107
rect 2289 1102 2318 1107
rect 2377 1102 2454 1107
rect 2521 1107 2526 1112
rect 2521 1102 2638 1107
rect 1185 1097 1190 1102
rect 217 1092 270 1097
rect 265 1077 270 1092
rect 441 1092 494 1097
rect 585 1092 1190 1097
rect 1209 1092 1742 1097
rect 1977 1092 2038 1097
rect 2113 1092 2214 1097
rect 2257 1092 2358 1097
rect 2385 1092 2510 1097
rect 441 1077 446 1092
rect 465 1087 470 1092
rect 1785 1087 1958 1092
rect 465 1082 686 1087
rect 881 1082 1006 1087
rect 1057 1082 1086 1087
rect 1281 1082 1502 1087
rect 1553 1082 1614 1087
rect 1633 1082 1790 1087
rect 1953 1082 2014 1087
rect 2233 1082 2270 1087
rect 2345 1082 2438 1087
rect 705 1077 830 1082
rect 1081 1077 1286 1082
rect 2089 1077 2214 1082
rect 265 1072 446 1077
rect 625 1072 710 1077
rect 825 1072 854 1077
rect 1425 1072 1638 1077
rect 1801 1072 1966 1077
rect 2017 1072 2094 1077
rect 2209 1072 2262 1077
rect 2273 1072 2542 1077
rect 897 1067 1030 1072
rect 1305 1067 1406 1072
rect 1633 1067 1806 1072
rect 2017 1067 2022 1072
rect 673 1062 902 1067
rect 1025 1062 1054 1067
rect 1129 1062 1262 1067
rect 1281 1062 1310 1067
rect 1401 1062 1614 1067
rect 1825 1062 2022 1067
rect 2105 1062 2134 1067
rect 2153 1062 2446 1067
rect 673 1057 678 1062
rect 1129 1057 1134 1062
rect 497 1052 678 1057
rect 697 1052 790 1057
rect 865 1052 1046 1057
rect 1089 1052 1134 1057
rect 1257 1057 1262 1062
rect 1257 1052 1606 1057
rect 1633 1052 1750 1057
rect 1937 1052 2518 1057
rect 1041 1047 1046 1052
rect 1633 1047 1638 1052
rect 401 1042 478 1047
rect 897 1042 982 1047
rect 1041 1042 1078 1047
rect 1145 1042 1262 1047
rect 1417 1042 1486 1047
rect 1505 1042 1638 1047
rect 1745 1047 1750 1052
rect 1809 1047 1918 1052
rect 1745 1042 1814 1047
rect 1913 1042 2174 1047
rect 2281 1042 2342 1047
rect 2353 1042 2486 1047
rect 1073 1037 1078 1042
rect 1257 1037 1422 1042
rect 225 1032 294 1037
rect 617 1032 686 1037
rect 617 1027 622 1032
rect 273 1022 390 1027
rect 73 1012 294 1017
rect 305 997 310 1022
rect 385 1017 390 1022
rect 489 1022 622 1027
rect 681 1027 686 1032
rect 769 1032 1054 1037
rect 1073 1032 1238 1037
rect 1497 1032 1734 1037
rect 1825 1032 2406 1037
rect 2625 1032 2662 1037
rect 769 1027 774 1032
rect 681 1022 774 1027
rect 785 1022 966 1027
rect 1193 1022 1222 1027
rect 489 1017 494 1022
rect 977 1017 1198 1022
rect 1233 1017 1238 1032
rect 1273 1022 1342 1027
rect 1361 1022 1534 1027
rect 1705 1022 1894 1027
rect 1905 1022 1982 1027
rect 2073 1022 2110 1027
rect 2201 1022 2510 1027
rect 1273 1017 1278 1022
rect 385 1012 494 1017
rect 633 1012 982 1017
rect 1233 1012 1278 1017
rect 1337 1017 1342 1022
rect 1529 1017 1710 1022
rect 1905 1017 1910 1022
rect 1337 1012 1398 1017
rect 1729 1012 1766 1017
rect 1801 1012 1910 1017
rect 1953 1012 2494 1017
rect 2609 1012 2638 1017
rect 1393 1007 1510 1012
rect 521 1002 630 1007
rect 841 1002 894 1007
rect 1025 1002 1046 1007
rect 1057 1002 1126 1007
rect 1289 1002 1374 1007
rect 1505 1002 1614 1007
rect 1705 1002 1854 1007
rect 2025 1002 2142 1007
rect 2257 1002 2390 1007
rect 2425 1002 2542 1007
rect 729 997 822 1002
rect 1609 997 1614 1002
rect 1849 997 2030 1002
rect 289 992 310 997
rect 553 992 662 997
rect 705 992 734 997
rect 817 992 1486 997
rect 1609 992 1830 997
rect 2049 992 2070 997
rect 2121 992 2566 997
rect 425 982 934 987
rect 1001 982 1510 987
rect 1521 982 1598 987
rect 1665 982 1734 987
rect 1785 982 1822 987
rect 1897 982 1966 987
rect 2041 982 2118 987
rect 2145 982 2342 987
rect 2393 982 2438 987
rect 2465 982 2614 987
rect 457 972 486 977
rect 673 972 782 977
rect 897 972 1062 977
rect 1097 972 1582 977
rect 1745 972 1846 977
rect 1961 972 2078 977
rect 2193 972 2310 977
rect 2401 972 2494 977
rect 481 967 486 972
rect 569 967 678 972
rect 2193 967 2198 972
rect 481 962 574 967
rect 697 962 806 967
rect 1089 962 1174 967
rect 1193 962 1734 967
rect 1761 962 2198 967
rect 2209 962 2350 967
rect 2449 962 2502 967
rect 1089 957 1094 962
rect 233 952 286 957
rect 593 952 614 957
rect 745 952 966 957
rect 993 952 1118 957
rect 1249 952 1382 957
rect 1489 952 2254 957
rect 321 942 430 947
rect 609 942 638 947
rect 665 942 710 947
rect 929 942 966 947
rect 1025 942 1166 947
rect 745 937 910 942
rect 1025 937 1030 942
rect 1249 937 1254 952
rect 1489 947 1494 952
rect 1265 942 1342 947
rect 1377 942 1494 947
rect 1513 942 1574 947
rect 1705 942 1758 947
rect 1769 942 1798 947
rect 1809 942 1942 947
rect 1993 942 2206 947
rect 2561 942 2638 947
rect 1569 937 1686 942
rect 377 932 518 937
rect 569 932 598 937
rect 593 927 598 932
rect 665 932 750 937
rect 905 932 1030 937
rect 1137 932 1254 937
rect 1681 932 1790 937
rect 665 927 670 932
rect 1313 927 1550 932
rect 1809 927 1814 942
rect 1873 932 1918 937
rect 1937 932 1942 942
rect 1953 932 2158 937
rect 2305 932 2342 937
rect 2209 927 2286 932
rect 497 922 558 927
rect 593 922 670 927
rect 761 922 894 927
rect 1025 922 1182 927
rect 1265 922 1318 927
rect 1545 922 1638 927
rect 1785 922 1814 927
rect 1889 922 1934 927
rect 1969 922 2214 927
rect 2281 922 2438 927
rect 377 917 478 922
rect 1177 917 1270 922
rect 1697 917 1790 922
rect 105 912 166 917
rect 289 912 382 917
rect 473 912 510 917
rect 833 912 1158 917
rect 1329 912 1366 917
rect 1425 912 1702 917
rect 1865 912 2158 917
rect 2225 912 2262 917
rect 2401 912 2534 917
rect 393 902 630 907
rect 745 902 822 907
rect 929 902 958 907
rect 1049 902 1326 907
rect 1321 897 1326 902
rect 1417 902 2262 907
rect 2297 902 2382 907
rect 2441 902 2486 907
rect 2537 902 2598 907
rect 1417 897 1422 902
rect 385 892 590 897
rect 825 892 1150 897
rect 1321 892 1422 897
rect 1465 892 1718 897
rect 1801 892 1846 897
rect 1857 892 1918 897
rect 2017 892 2046 897
rect 2145 892 2246 897
rect 2433 892 2454 897
rect 2553 892 2598 897
rect 313 882 438 887
rect 481 882 638 887
rect 953 882 1094 887
rect 1153 882 1190 887
rect 1209 882 1302 887
rect 1897 882 1926 887
rect 1937 882 2086 887
rect 2121 882 2166 887
rect 2553 882 2582 887
rect 809 877 934 882
rect 1209 877 1214 882
rect 473 872 526 877
rect 545 872 574 877
rect 649 872 710 877
rect 785 872 814 877
rect 929 872 1214 877
rect 1297 877 1302 882
rect 1393 877 1766 882
rect 1801 877 1878 882
rect 1297 872 1398 877
rect 1761 872 1806 877
rect 1873 872 2006 877
rect 2041 872 2078 877
rect 2113 872 2230 877
rect 497 857 502 872
rect 569 867 654 872
rect 713 862 1062 867
rect 1073 862 1286 867
rect 1409 862 1510 867
rect 1545 862 1750 867
rect 1817 862 2366 867
rect 713 857 718 862
rect 1073 857 1078 862
rect 137 852 206 857
rect 497 852 718 857
rect 937 852 1078 857
rect 1209 852 1254 857
rect 1313 852 1366 857
rect 1505 852 1510 862
rect 1641 852 1766 857
rect 1913 852 1990 857
rect 2009 852 2214 857
rect 137 847 142 852
rect 113 842 142 847
rect 201 847 206 852
rect 737 847 942 852
rect 1097 847 1190 852
rect 1505 847 1622 852
rect 1809 847 1894 852
rect 1985 847 1990 852
rect 201 842 230 847
rect 281 842 366 847
rect 737 837 742 847
rect 961 842 1102 847
rect 1185 842 1310 847
rect 1409 842 1438 847
rect 1449 842 1486 847
rect 1617 842 1678 847
rect 1777 842 1814 847
rect 1889 842 1958 847
rect 1985 842 2190 847
rect 2489 842 2558 847
rect 1673 837 1782 842
rect 2489 837 2494 842
rect 241 832 310 837
rect 449 832 742 837
rect 753 832 806 837
rect 865 832 1542 837
rect 1601 832 1654 837
rect 1825 832 1878 837
rect 1929 832 1982 837
rect 2017 832 2062 837
rect 2265 832 2302 837
rect 2465 832 2494 837
rect 2553 837 2558 842
rect 2553 832 2582 837
rect 89 827 158 832
rect 345 827 454 832
rect 801 827 806 832
rect 1601 827 1606 832
rect 65 822 94 827
rect 153 822 230 827
rect 321 822 350 827
rect 593 822 614 827
rect 625 822 662 827
rect 801 822 1254 827
rect 1289 822 1406 827
rect 225 817 326 822
rect 473 817 574 822
rect 81 812 142 817
rect 361 812 478 817
rect 569 812 838 817
rect 1001 812 1038 817
rect 1081 812 1190 817
rect 865 807 982 812
rect 1201 807 1206 817
rect 1353 812 1382 817
rect 1425 807 1430 827
rect 1489 822 1606 827
rect 1673 822 1806 827
rect 1921 822 1950 827
rect 1969 822 2094 827
rect 2169 822 2350 827
rect 2417 822 2646 827
rect 1673 817 1678 822
rect 1577 812 1678 817
rect 1801 817 1806 822
rect 1801 812 2262 817
rect 2377 812 2550 817
rect 193 802 414 807
rect 433 802 486 807
rect 513 802 558 807
rect 577 802 638 807
rect 673 802 702 807
rect 577 797 582 802
rect 81 792 166 797
rect 185 792 262 797
rect 465 792 582 797
rect 697 797 702 802
rect 841 802 870 807
rect 977 802 1094 807
rect 1113 802 1206 807
rect 1305 802 1446 807
rect 841 797 846 802
rect 1089 797 1094 802
rect 1441 797 1446 802
rect 1665 802 1790 807
rect 1897 802 1974 807
rect 2001 802 2070 807
rect 2121 802 2190 807
rect 1665 797 1670 802
rect 1969 797 1974 802
rect 2257 797 2262 812
rect 2345 802 2430 807
rect 2521 802 2582 807
rect 697 792 846 797
rect 889 792 942 797
rect 961 792 1006 797
rect 1033 792 1070 797
rect 1089 792 1430 797
rect 1441 792 1670 797
rect 1681 792 1958 797
rect 1969 792 2182 797
rect 2257 792 2574 797
rect 1953 787 1958 792
rect 2177 787 2182 792
rect 169 782 286 787
rect 385 782 486 787
rect 537 782 590 787
rect 865 782 886 787
rect 1073 782 1134 787
rect 1145 782 1550 787
rect 1625 782 1646 787
rect 1665 782 1702 787
rect 1785 782 1926 787
rect 1953 782 1982 787
rect 2017 782 2046 787
rect 2057 782 2150 787
rect 2177 782 2430 787
rect 2457 782 2542 787
rect 1665 777 1670 782
rect 2401 777 2406 782
rect 73 772 654 777
rect 665 772 710 777
rect 737 772 918 777
rect 985 772 1446 777
rect 1521 772 1670 777
rect 1801 772 1846 777
rect 1881 772 2142 777
rect 737 767 742 772
rect 2137 767 2142 772
rect 2233 772 2382 777
rect 2401 772 2614 777
rect 2233 767 2238 772
rect 177 762 406 767
rect 561 762 742 767
rect 849 762 998 767
rect 1009 762 1270 767
rect 1281 762 1390 767
rect 1425 762 1550 767
rect 1617 762 1710 767
rect 1729 762 1798 767
rect 1817 762 1894 767
rect 1945 762 1990 767
rect 2137 762 2238 767
rect 2257 762 2294 767
rect 2393 762 2446 767
rect 2513 762 2558 767
rect 401 757 550 762
rect 849 757 854 762
rect 1793 757 1798 762
rect 161 752 294 757
rect 545 752 574 757
rect 753 752 854 757
rect 897 752 998 757
rect 1113 752 1190 757
rect 1201 752 1262 757
rect 1361 752 1782 757
rect 1793 752 2054 757
rect 2065 752 2118 757
rect 2401 752 2502 757
rect 2569 752 2630 757
rect 569 747 758 752
rect 993 747 1118 752
rect 1201 747 1206 752
rect 97 727 102 747
rect 369 742 550 747
rect 369 737 374 742
rect 545 737 550 742
rect 817 742 910 747
rect 817 737 822 742
rect 1137 737 1142 747
rect 1169 742 1206 747
rect 1217 742 1294 747
rect 1337 742 1510 747
rect 1625 742 1702 747
rect 2009 742 2062 747
rect 2241 742 2278 747
rect 1697 737 1702 742
rect 1785 737 1918 742
rect 2089 737 2222 742
rect 2401 737 2406 752
rect 2497 747 2574 752
rect 201 732 374 737
rect 385 732 414 737
rect 497 732 526 737
rect 545 732 822 737
rect 841 732 1046 737
rect 1137 732 1198 737
rect 1353 732 1390 737
rect 1409 732 1438 737
rect 1593 732 1654 737
rect 1697 732 1790 737
rect 1913 732 2014 737
rect 2065 732 2094 737
rect 2217 732 2406 737
rect 2537 732 2646 737
rect 409 727 502 732
rect 2065 727 2070 732
rect 97 722 118 727
rect 1305 722 1470 727
rect 1681 722 1734 727
rect 1801 722 1902 727
rect 1025 717 1262 722
rect 1681 717 1686 722
rect 1897 717 1902 722
rect 2041 722 2070 727
rect 2081 722 2430 727
rect 2041 717 2046 722
rect 97 712 190 717
rect 441 712 646 717
rect 737 712 806 717
rect 865 712 1030 717
rect 1257 712 1294 717
rect 1353 712 1598 717
rect 1617 712 1686 717
rect 1729 712 1814 717
rect 1897 712 2046 717
rect 2065 712 2102 717
rect 2217 712 2286 717
rect 2577 712 2638 717
rect 1289 707 1358 712
rect 2353 707 2422 712
rect 273 702 438 707
rect 433 697 438 702
rect 553 702 582 707
rect 1041 702 1246 707
rect 1377 702 1558 707
rect 1569 702 1662 707
rect 1737 702 1814 707
rect 1841 702 1878 707
rect 2121 702 2166 707
rect 2233 702 2278 707
rect 2329 702 2358 707
rect 2417 702 2566 707
rect 553 697 558 702
rect 433 692 558 697
rect 609 692 790 697
rect 1217 692 1366 697
rect 609 687 614 692
rect 385 682 414 687
rect 409 677 414 682
rect 593 682 614 687
rect 785 687 790 692
rect 977 687 1198 692
rect 1377 687 1382 702
rect 2561 697 2566 702
rect 2641 702 2670 707
rect 2641 697 2646 702
rect 1393 692 1414 697
rect 1537 692 2022 697
rect 2137 692 2270 697
rect 2289 692 2326 697
rect 2369 692 2406 697
rect 2561 692 2646 697
rect 785 682 814 687
rect 849 682 982 687
rect 1193 682 1382 687
rect 1465 682 1542 687
rect 1553 682 1590 687
rect 1665 682 1886 687
rect 2033 682 2174 687
rect 2249 682 2310 687
rect 593 677 598 682
rect 409 672 598 677
rect 617 672 726 677
rect 769 672 838 677
rect 833 667 838 672
rect 993 672 1022 677
rect 1033 672 1878 677
rect 1969 672 2494 677
rect 993 667 998 672
rect 689 662 710 667
rect 793 662 814 667
rect 833 662 998 667
rect 1097 662 1134 667
rect 1257 662 1646 667
rect 1745 662 2094 667
rect 1665 657 1750 662
rect 2113 657 2238 662
rect 2289 657 2382 662
rect 553 652 646 657
rect 665 652 798 657
rect 1025 652 1302 657
rect 1361 652 1670 657
rect 1769 652 1806 657
rect 1921 652 1974 657
rect 2025 652 2118 657
rect 2233 652 2294 657
rect 2377 652 2470 657
rect 553 647 558 652
rect 425 642 510 647
rect 529 642 558 647
rect 641 647 646 652
rect 641 642 846 647
rect 961 642 998 647
rect 1065 642 1310 647
rect 1377 642 1398 647
rect 1417 642 1582 647
rect 1641 642 2222 647
rect 2305 642 2366 647
rect 2553 642 2606 647
rect 425 637 430 642
rect 361 632 430 637
rect 505 637 510 642
rect 993 637 998 642
rect 505 632 622 637
rect 657 632 982 637
rect 993 632 1166 637
rect 1201 632 1726 637
rect 1737 632 2014 637
rect 2041 632 2094 637
rect 2145 632 2382 637
rect 2401 632 2486 637
rect 2401 627 2406 632
rect 97 622 150 627
rect 161 622 190 627
rect 457 622 566 627
rect 585 622 670 627
rect 753 622 782 627
rect 801 622 886 627
rect 937 622 1998 627
rect 2201 622 2230 627
rect 2313 622 2342 627
rect 2361 622 2406 627
rect 2481 627 2486 632
rect 2481 622 2510 627
rect 561 617 566 622
rect 665 617 758 622
rect 2225 617 2318 622
rect 265 612 334 617
rect 361 612 470 617
rect 561 612 646 617
rect 777 612 1390 617
rect 1409 612 1494 617
rect 1593 612 1934 617
rect 2017 612 2102 617
rect 2417 612 2446 617
rect 2521 612 2590 617
rect 2441 607 2526 612
rect 433 602 566 607
rect 593 602 726 607
rect 737 602 894 607
rect 1089 602 1286 607
rect 1361 602 1670 607
rect 1705 602 1742 607
rect 1833 602 2126 607
rect 2185 602 2342 607
rect 721 597 726 602
rect 921 597 1054 602
rect 1665 597 1670 602
rect 721 592 926 597
rect 1049 592 1078 597
rect 1209 592 1278 597
rect 1465 592 1494 597
rect 1665 592 2134 597
rect 2153 592 2198 597
rect 2345 592 2518 597
rect 2537 592 2670 597
rect 2193 587 2350 592
rect 2513 587 2518 592
rect 153 582 270 587
rect 689 582 766 587
rect 937 582 1390 587
rect 1441 582 1478 587
rect 1801 582 1894 587
rect 1977 582 2070 587
rect 2081 582 2174 587
rect 2369 582 2422 587
rect 2513 582 2558 587
rect 841 577 918 582
rect 1665 577 1806 582
rect 1889 577 1982 582
rect 209 572 278 577
rect 393 572 430 577
rect 465 572 518 577
rect 633 572 846 577
rect 913 572 1094 577
rect 1249 572 1598 577
rect 1665 567 1670 577
rect 1825 572 1870 577
rect 2001 572 2038 577
rect 2049 572 2118 577
rect 2193 572 2294 577
rect 2193 567 2198 572
rect 521 562 606 567
rect 625 562 654 567
rect 857 562 886 567
rect 937 562 1102 567
rect 1169 562 1222 567
rect 1353 562 1670 567
rect 1681 562 1718 567
rect 1793 562 1830 567
rect 1921 562 2198 567
rect 2289 567 2294 572
rect 2289 562 2454 567
rect 649 557 862 562
rect 145 552 230 557
rect 297 552 366 557
rect 385 552 502 557
rect 969 552 1782 557
rect 1841 552 2086 557
rect 2137 552 2278 557
rect 385 547 390 552
rect 89 542 158 547
rect 177 542 310 547
rect 321 542 390 547
rect 497 547 502 552
rect 1777 547 1846 552
rect 2273 547 2278 552
rect 2385 552 2646 557
rect 2385 547 2390 552
rect 497 542 542 547
rect 561 542 774 547
rect 793 542 998 547
rect 1073 542 1126 547
rect 1193 542 1262 547
rect 1353 542 1486 547
rect 1497 542 1590 547
rect 1657 542 1686 547
rect 1985 542 2014 547
rect 305 537 310 542
rect 561 537 566 542
rect 305 532 382 537
rect 409 532 566 537
rect 769 537 774 542
rect 2009 537 2014 542
rect 2073 542 2198 547
rect 2273 542 2390 547
rect 2073 537 2078 542
rect 769 532 1518 537
rect 1769 532 1862 537
rect 2009 532 2078 537
rect 2097 532 2174 537
rect 2201 532 2254 537
rect 2409 532 2598 537
rect 585 527 750 532
rect 1513 527 1654 532
rect 89 522 118 527
rect 201 522 294 527
rect 353 522 590 527
rect 745 522 950 527
rect 1049 522 1222 527
rect 1265 522 1334 527
rect 1345 522 1494 527
rect 1649 522 1886 527
rect 2241 522 2294 527
rect 2313 522 2374 527
rect 2545 522 2662 527
rect 945 517 1054 522
rect 1329 517 1334 522
rect 2289 517 2294 522
rect 113 512 174 517
rect 449 512 622 517
rect 633 512 662 517
rect 689 512 774 517
rect 849 512 926 517
rect 1073 512 1118 517
rect 1193 512 1246 517
rect 1329 512 1414 517
rect 1465 512 1654 517
rect 1897 512 1934 517
rect 1961 512 2038 517
rect 2289 512 2342 517
rect 2377 512 2582 517
rect 1673 507 1878 512
rect 2161 507 2270 512
rect 177 502 390 507
rect 425 502 1678 507
rect 1873 502 1926 507
rect 2041 502 2166 507
rect 2265 502 2318 507
rect 2433 502 2470 507
rect 2561 502 2598 507
rect 385 487 390 502
rect 401 492 494 497
rect 521 492 550 497
rect 737 492 862 497
rect 1185 492 1382 497
rect 1481 492 1550 497
rect 1593 492 1750 497
rect 1761 492 2070 497
rect 2177 492 2542 497
rect 545 487 742 492
rect 881 487 1166 492
rect 1745 487 1750 492
rect 385 482 462 487
rect 761 482 886 487
rect 1161 482 1366 487
rect 1457 482 1566 487
rect 1745 482 1790 487
rect 1961 482 1990 487
rect 2321 482 2502 487
rect 1785 477 1966 482
rect 2153 477 2278 482
rect 513 472 750 477
rect 817 472 990 477
rect 1049 472 1118 477
rect 1129 472 1198 477
rect 1225 472 1766 477
rect 1761 467 1766 472
rect 2001 472 2158 477
rect 2273 472 2454 477
rect 2001 467 2006 472
rect 2449 467 2454 472
rect 2553 472 2678 477
rect 2553 467 2558 472
rect 793 462 974 467
rect 1105 462 1182 467
rect 1193 462 1390 467
rect 1577 462 1606 467
rect 1713 462 1742 467
rect 1761 462 2006 467
rect 2169 462 2262 467
rect 993 457 1086 462
rect 1385 457 1558 462
rect 1601 457 1718 462
rect 2257 457 2262 462
rect 2377 462 2406 467
rect 2449 462 2558 467
rect 2377 457 2382 462
rect 657 452 750 457
rect 801 452 998 457
rect 1081 452 1366 457
rect 1553 447 1558 457
rect 2257 452 2382 457
rect 353 442 422 447
rect 561 442 646 447
rect 713 442 822 447
rect 913 442 1134 447
rect 1177 442 1214 447
rect 1345 442 1422 447
rect 1505 442 1542 447
rect 1553 442 1638 447
rect 1665 442 1718 447
rect 1761 442 1958 447
rect 1977 442 2022 447
rect 2033 442 2126 447
rect 2145 442 2238 447
rect 641 437 718 442
rect 817 437 918 442
rect 1345 437 1350 442
rect 1761 437 1766 442
rect 481 432 590 437
rect 737 432 798 437
rect 793 427 798 432
rect 937 432 1350 437
rect 1369 432 1438 437
rect 1489 432 1766 437
rect 1953 437 1958 442
rect 2145 437 2150 442
rect 1953 432 2150 437
rect 2233 437 2238 442
rect 2233 432 2262 437
rect 2313 432 2534 437
rect 2617 432 2662 437
rect 937 427 942 432
rect 97 422 214 427
rect 313 422 358 427
rect 401 422 534 427
rect 353 417 358 422
rect 529 417 534 422
rect 625 422 718 427
rect 793 422 942 427
rect 1017 422 1214 427
rect 1401 422 1446 427
rect 1473 422 1526 427
rect 1585 422 1646 427
rect 1697 422 1758 427
rect 625 417 630 422
rect 249 412 342 417
rect 353 412 430 417
rect 529 412 630 417
rect 713 417 718 422
rect 1889 417 1894 427
rect 2057 422 2150 427
rect 2161 422 2342 427
rect 713 412 774 417
rect 1009 412 1070 417
rect 1169 412 1270 417
rect 1289 412 1366 417
rect 1649 412 1870 417
rect 1889 412 1934 417
rect 1961 412 1998 417
rect 1089 407 1174 412
rect 1289 407 1294 412
rect 257 402 734 407
rect 753 402 806 407
rect 825 402 958 407
rect 977 402 1094 407
rect 1193 402 1294 407
rect 1361 407 1366 412
rect 2161 407 2166 422
rect 2233 412 2350 417
rect 1361 402 2166 407
rect 2337 402 2414 407
rect 753 397 758 402
rect 825 397 830 402
rect 265 392 422 397
rect 569 392 598 397
rect 689 392 758 397
rect 777 392 830 397
rect 953 397 958 402
rect 953 392 1342 397
rect 1401 392 1486 397
rect 1521 392 1566 397
rect 1601 392 1686 397
rect 1737 392 1838 397
rect 1897 392 1942 397
rect 441 387 534 392
rect 593 387 694 392
rect 321 382 446 387
rect 529 382 558 387
rect 713 382 830 387
rect 1057 382 1262 387
rect 1345 382 1398 387
rect 1553 382 1654 387
rect 1913 382 2302 387
rect 849 377 974 382
rect 1753 377 1854 382
rect 177 372 246 377
rect 289 372 526 377
rect 537 372 662 377
rect 697 372 854 377
rect 969 372 998 377
rect 1009 372 1542 377
rect 1665 372 1758 377
rect 1849 372 1878 377
rect 177 367 182 372
rect 65 362 182 367
rect 241 367 246 372
rect 241 362 318 367
rect 425 362 486 367
rect 193 352 222 357
rect 305 352 334 357
rect 217 347 310 352
rect 657 347 662 372
rect 1009 367 1014 372
rect 1537 367 1670 372
rect 769 362 1014 367
rect 1105 362 1190 367
rect 1769 362 1814 367
rect 1889 362 1958 367
rect 2097 362 2182 367
rect 2601 362 2662 367
rect 1185 357 1190 362
rect 1249 357 1478 362
rect 681 352 742 357
rect 849 352 998 357
rect 1105 352 1166 357
rect 1185 352 1254 357
rect 1473 352 2118 357
rect 2129 352 2350 357
rect 2529 352 2622 357
rect 2113 347 2118 352
rect 345 342 382 347
rect 521 342 590 347
rect 657 342 686 347
rect 753 342 1198 347
rect 1265 342 1342 347
rect 1385 342 1462 347
rect 1545 342 1574 347
rect 1657 342 1686 347
rect 521 337 526 342
rect 281 332 350 337
rect 497 332 526 337
rect 585 337 590 342
rect 681 337 758 342
rect 1569 337 1662 342
rect 1793 337 1798 347
rect 1817 342 1902 347
rect 1921 342 1950 347
rect 2113 342 2206 347
rect 585 332 614 337
rect 865 332 1206 337
rect 1689 332 1798 337
rect 2201 337 2206 342
rect 2329 342 2358 347
rect 2329 337 2334 342
rect 2201 332 2334 337
rect 2425 332 2470 337
rect 385 322 478 327
rect 721 322 910 327
rect 953 322 1022 327
rect 1129 322 1190 327
rect 1225 322 1278 327
rect 1305 322 1358 327
rect 1377 322 1638 327
rect 1873 322 1910 327
rect 1969 322 2094 327
rect 2129 322 2182 327
rect 385 317 390 322
rect 361 312 390 317
rect 473 317 478 322
rect 1377 317 1382 322
rect 473 312 1382 317
rect 1633 317 1638 322
rect 1737 317 1854 322
rect 1969 317 1974 322
rect 1633 312 1742 317
rect 1849 312 1974 317
rect 2089 317 2094 322
rect 2089 312 2326 317
rect 313 302 502 307
rect 825 302 894 307
rect 945 302 1022 307
rect 1137 302 1222 307
rect 1233 302 1622 307
rect 1753 302 1886 307
rect 1905 302 1950 307
rect 2137 302 2174 307
rect 2281 302 2374 307
rect 689 297 806 302
rect 1233 297 1238 302
rect 97 292 174 297
rect 425 292 454 297
rect 449 287 454 292
rect 513 292 694 297
rect 801 292 1238 297
rect 1249 292 1518 297
rect 1737 292 2038 297
rect 2057 292 2134 297
rect 2385 292 2646 297
rect 513 287 518 292
rect 2033 287 2038 292
rect 2385 287 2390 292
rect 449 282 518 287
rect 705 282 918 287
rect 1017 282 1166 287
rect 1409 282 1470 287
rect 1561 282 1918 287
rect 2033 282 2078 287
rect 2145 282 2390 287
rect 1185 277 1294 282
rect 2073 277 2150 282
rect 609 272 1190 277
rect 1289 272 1582 277
rect 1745 272 2054 277
rect 1577 267 1750 272
rect 521 262 838 267
rect 929 262 1118 267
rect 1193 262 1278 267
rect 1473 262 1558 267
rect 1825 262 1854 267
rect 2065 262 2150 267
rect 2329 262 2574 267
rect 1297 257 1454 262
rect 1849 257 2070 262
rect 2329 257 2334 262
rect 441 252 574 257
rect 745 252 1302 257
rect 1449 252 1582 257
rect 1633 252 1694 257
rect 2145 252 2334 257
rect 2569 257 2574 262
rect 2569 252 2598 257
rect 593 247 726 252
rect 473 242 598 247
rect 721 242 1510 247
rect 1841 242 1958 247
rect 1977 242 2094 247
rect 1841 237 1846 242
rect 217 232 318 237
rect 529 232 590 237
rect 617 232 798 237
rect 817 232 1262 237
rect 1361 232 1846 237
rect 1953 237 1958 242
rect 1953 232 2038 237
rect 2105 232 2614 237
rect 369 222 670 227
rect 689 217 758 222
rect 817 217 822 232
rect 1257 227 1366 232
rect 2033 227 2110 232
rect 913 222 1214 227
rect 1385 222 1414 227
rect 1465 222 1542 227
rect 1761 222 2014 227
rect 2217 222 2246 227
rect 2313 222 2398 227
rect 1561 217 1742 222
rect 401 212 694 217
rect 753 212 822 217
rect 841 212 1566 217
rect 1737 212 1782 217
rect 2025 212 2150 217
rect 2177 212 2454 217
rect 2473 212 2574 217
rect 1777 207 2030 212
rect 2473 207 2478 212
rect 353 202 454 207
rect 681 202 742 207
rect 817 202 934 207
rect 953 202 1110 207
rect 1409 202 1438 207
rect 1489 202 1550 207
rect 1569 202 1758 207
rect 2089 202 2254 207
rect 2273 202 2478 207
rect 2569 207 2574 212
rect 2569 202 2598 207
rect 521 197 662 202
rect 817 197 822 202
rect 1569 197 1574 202
rect 2273 197 2278 202
rect 329 192 358 197
rect 465 192 526 197
rect 657 192 822 197
rect 833 192 926 197
rect 985 192 1046 197
rect 1209 192 1326 197
rect 1481 192 1502 197
rect 1521 192 1574 197
rect 1593 192 1670 197
rect 1777 192 2078 197
rect 2153 192 2278 197
rect 2369 192 2438 197
rect 2457 192 2558 197
rect 353 187 470 192
rect 1521 187 1526 192
rect 537 182 694 187
rect 1145 182 1278 187
rect 1441 182 1526 187
rect 1297 177 1366 182
rect 1777 177 1782 192
rect 2073 187 2158 192
rect 2177 182 2438 187
rect 393 172 494 177
rect 537 172 558 177
rect 665 172 830 177
rect 897 172 974 177
rect 1153 172 1302 177
rect 1361 172 1782 177
rect 2137 172 2230 177
rect 505 162 558 167
rect 785 162 862 167
rect 937 162 998 167
rect 1161 162 1246 167
rect 1257 162 1350 167
rect 1801 162 1918 167
rect 1369 157 1518 162
rect 1801 157 1806 162
rect 169 152 326 157
rect 377 152 1374 157
rect 1513 152 1806 157
rect 1913 157 1918 162
rect 1961 162 2118 167
rect 2281 162 2366 167
rect 2385 162 2502 167
rect 1961 157 1966 162
rect 1913 152 1966 157
rect 2113 157 2118 162
rect 2385 157 2390 162
rect 2113 152 2390 157
rect 2409 152 2566 157
rect 321 137 326 152
rect 345 142 446 147
rect 481 142 1070 147
rect 1257 142 1414 147
rect 1433 142 1502 147
rect 2017 142 2094 147
rect 2353 142 2558 147
rect 1065 137 1262 142
rect 1409 137 1414 142
rect 2017 137 2022 142
rect 2089 137 2278 142
rect 321 132 678 137
rect 1409 132 1438 137
rect 1513 132 2022 137
rect 2273 132 2518 137
rect 673 127 678 132
rect 761 127 1046 132
rect 1433 127 1518 132
rect 441 122 470 127
rect 633 122 662 127
rect 673 122 766 127
rect 1041 122 1094 127
rect 1217 122 1326 127
rect 2033 122 2246 127
rect 2257 122 2294 127
rect 465 117 574 122
rect 633 117 638 122
rect 297 112 382 117
rect 569 112 638 117
rect 785 112 1046 117
rect 1089 107 1094 122
rect 1113 112 1198 117
rect 1345 112 1462 117
rect 1793 112 1870 117
rect 1953 112 2086 117
rect 2097 112 2166 117
rect 1345 107 1350 112
rect 521 102 550 107
rect 545 97 550 102
rect 881 102 934 107
rect 1089 102 1110 107
rect 881 97 886 102
rect 545 92 886 97
rect 929 97 934 102
rect 1105 97 1110 102
rect 1209 102 1350 107
rect 1457 107 1462 112
rect 1457 102 2030 107
rect 1209 97 1214 102
rect 2025 97 2030 102
rect 2097 97 2102 112
rect 2161 107 2166 112
rect 2289 112 2398 117
rect 2289 107 2294 112
rect 2393 107 2398 112
rect 2457 112 2622 117
rect 2457 107 2462 112
rect 2113 102 2142 107
rect 2161 102 2294 107
rect 2313 102 2374 107
rect 2393 102 2462 107
rect 929 92 1078 97
rect 1105 92 1214 97
rect 1305 92 1358 97
rect 1073 77 1078 92
rect 1305 77 1310 92
rect 1353 87 1358 92
rect 1417 92 1446 97
rect 2025 92 2102 97
rect 1417 87 1422 92
rect 1353 82 1422 87
rect 2137 87 2142 102
rect 2313 87 2318 102
rect 2137 82 2318 87
rect 1073 72 1310 77
use AND2X2  AND2X2_0
timestamp 1710841341
transform 1 0 744 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1710841341
transform 1 0 680 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1710841341
transform 1 0 880 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1710841341
transform 1 0 696 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1710841341
transform 1 0 520 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1710841341
transform 1 0 2392 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1710841341
transform 1 0 2320 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1710841341
transform 1 0 1696 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1710841341
transform 1 0 1800 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1710841341
transform 1 0 2376 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1710841341
transform 1 0 960 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1710841341
transform 1 0 2160 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1710841341
transform 1 0 1536 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1710841341
transform 1 0 304 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1710841341
transform 1 0 2224 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1710841341
transform 1 0 1464 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1710841341
transform 1 0 1512 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1710841341
transform 1 0 1192 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1710841341
transform 1 0 1224 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1710841341
transform 1 0 544 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_20
timestamp 1710841341
transform 1 0 600 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1710841341
transform 1 0 672 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1710841341
transform 1 0 664 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_23
timestamp 1710841341
transform 1 0 440 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1710841341
transform 1 0 480 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_25
timestamp 1710841341
transform 1 0 408 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_26
timestamp 1710841341
transform 1 0 592 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_27
timestamp 1710841341
transform 1 0 584 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_28
timestamp 1710841341
transform 1 0 568 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_29
timestamp 1710841341
transform 1 0 792 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_30
timestamp 1710841341
transform 1 0 888 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_31
timestamp 1710841341
transform 1 0 1192 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_32
timestamp 1710841341
transform 1 0 480 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_33
timestamp 1710841341
transform 1 0 520 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_34
timestamp 1710841341
transform 1 0 1512 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_35
timestamp 1710841341
transform 1 0 1400 0 -1 370
box -8 -3 40 105
use AND2X2  AND2X2_36
timestamp 1710841341
transform 1 0 1408 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_37
timestamp 1710841341
transform 1 0 1552 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_38
timestamp 1710841341
transform 1 0 1656 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_39
timestamp 1710841341
transform 1 0 1504 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_40
timestamp 1710841341
transform 1 0 1704 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_41
timestamp 1710841341
transform 1 0 1728 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_42
timestamp 1710841341
transform 1 0 1728 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_43
timestamp 1710841341
transform 1 0 2496 0 -1 1170
box -8 -3 40 105
use AND2X2  AND2X2_44
timestamp 1710841341
transform 1 0 2416 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_45
timestamp 1710841341
transform 1 0 2192 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_46
timestamp 1710841341
transform 1 0 2360 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_47
timestamp 1710841341
transform 1 0 2344 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_48
timestamp 1710841341
transform 1 0 1896 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_49
timestamp 1710841341
transform 1 0 2088 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_50
timestamp 1710841341
transform 1 0 1896 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_51
timestamp 1710841341
transform 1 0 2040 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_52
timestamp 1710841341
transform 1 0 1984 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_53
timestamp 1710841341
transform 1 0 2272 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_54
timestamp 1710841341
transform 1 0 2200 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_55
timestamp 1710841341
transform 1 0 1552 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_56
timestamp 1710841341
transform 1 0 424 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_57
timestamp 1710841341
transform 1 0 160 0 1 2370
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1710841341
transform 1 0 240 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1710841341
transform 1 0 264 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1710841341
transform 1 0 200 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1710841341
transform 1 0 352 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1710841341
transform 1 0 584 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1710841341
transform 1 0 400 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1710841341
transform 1 0 496 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1710841341
transform 1 0 440 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1710841341
transform 1 0 744 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1710841341
transform 1 0 760 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1710841341
transform 1 0 1040 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1710841341
transform 1 0 1096 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1710841341
transform 1 0 288 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1710841341
transform 1 0 352 0 -1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1710841341
transform 1 0 792 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1710841341
transform 1 0 440 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1710841341
transform 1 0 1016 0 -1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1710841341
transform 1 0 856 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1710841341
transform 1 0 800 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1710841341
transform 1 0 1168 0 -1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1710841341
transform 1 0 1240 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1710841341
transform 1 0 1080 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1710841341
transform 1 0 1568 0 -1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1710841341
transform 1 0 1360 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1710841341
transform 1 0 1744 0 -1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1710841341
transform 1 0 1976 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1710841341
transform 1 0 1912 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_27
timestamp 1710841341
transform 1 0 1872 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_28
timestamp 1710841341
transform 1 0 1944 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_29
timestamp 1710841341
transform 1 0 2400 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_30
timestamp 1710841341
transform 1 0 2392 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_31
timestamp 1710841341
transform 1 0 2448 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_32
timestamp 1710841341
transform 1 0 2144 0 -1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_33
timestamp 1710841341
transform 1 0 2352 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_34
timestamp 1710841341
transform 1 0 2472 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_35
timestamp 1710841341
transform 1 0 2144 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_36
timestamp 1710841341
transform 1 0 2408 0 -1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_37
timestamp 1710841341
transform 1 0 2584 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_38
timestamp 1710841341
transform 1 0 2080 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_39
timestamp 1710841341
transform 1 0 2528 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_40
timestamp 1710841341
transform 1 0 2536 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_41
timestamp 1710841341
transform 1 0 2024 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_42
timestamp 1710841341
transform 1 0 2520 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_43
timestamp 1710841341
transform 1 0 800 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_44
timestamp 1710841341
transform 1 0 2632 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_45
timestamp 1710841341
transform 1 0 1008 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_46
timestamp 1710841341
transform 1 0 1880 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_47
timestamp 1710841341
transform 1 0 864 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_48
timestamp 1710841341
transform 1 0 1904 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_49
timestamp 1710841341
transform 1 0 2632 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_50
timestamp 1710841341
transform 1 0 2632 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_51
timestamp 1710841341
transform 1 0 2136 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_52
timestamp 1710841341
transform 1 0 2568 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_53
timestamp 1710841341
transform 1 0 2360 0 1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_54
timestamp 1710841341
transform 1 0 2408 0 -1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_55
timestamp 1710841341
transform 1 0 2008 0 1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_56
timestamp 1710841341
transform 1 0 2040 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_57
timestamp 1710841341
transform 1 0 2080 0 -1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_58
timestamp 1710841341
transform 1 0 1728 0 1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_59
timestamp 1710841341
transform 1 0 1584 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_60
timestamp 1710841341
transform 1 0 1560 0 1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_61
timestamp 1710841341
transform 1 0 1368 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_62
timestamp 1710841341
transform 1 0 1184 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_63
timestamp 1710841341
transform 1 0 944 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_64
timestamp 1710841341
transform 1 0 848 0 -1 1970
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1710841341
transform 1 0 272 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1710841341
transform 1 0 120 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1710841341
transform 1 0 288 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1710841341
transform 1 0 88 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1710841341
transform 1 0 240 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1710841341
transform 1 0 88 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1710841341
transform 1 0 448 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1710841341
transform 1 0 496 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1710841341
transform 1 0 848 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1710841341
transform 1 0 800 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1710841341
transform 1 0 952 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1710841341
transform 1 0 848 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1710841341
transform 1 0 400 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1710841341
transform 1 0 672 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1710841341
transform 1 0 728 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1710841341
transform 1 0 1416 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1710841341
transform 1 0 1464 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1710841341
transform 1 0 1896 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1710841341
transform 1 0 2208 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1710841341
transform 1 0 1568 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1710841341
transform 1 0 2304 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1710841341
transform 1 0 2184 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1710841341
transform 1 0 2256 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1710841341
transform 1 0 2144 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1710841341
transform 1 0 2176 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1710841341
transform 1 0 2024 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1710841341
transform 1 0 2032 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1710841341
transform 1 0 2224 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1710841341
transform 1 0 784 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1710841341
transform 1 0 1856 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1710841341
transform 1 0 1664 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1710841341
transform 1 0 1576 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1710841341
transform 1 0 1552 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1710841341
transform 1 0 1232 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1710841341
transform 1 0 1296 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1710841341
transform 1 0 1488 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1710841341
transform 1 0 1168 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1710841341
transform 1 0 1176 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1710841341
transform 1 0 1448 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1710841341
transform 1 0 1064 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1710841341
transform 1 0 1000 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1710841341
transform 1 0 1408 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1710841341
transform 1 0 808 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1710841341
transform 1 0 696 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1710841341
transform 1 0 184 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1710841341
transform 1 0 184 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1710841341
transform 1 0 152 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1710841341
transform 1 0 160 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1710841341
transform 1 0 160 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1710841341
transform 1 0 72 0 1 2170
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1710841341
transform 1 0 1344 0 -1 770
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1710841341
transform 1 0 1360 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1710841341
transform 1 0 1216 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1710841341
transform 1 0 1296 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1710841341
transform 1 0 1296 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1710841341
transform 1 0 1368 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1710841341
transform 1 0 2136 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1710841341
transform 1 0 1992 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1710841341
transform 1 0 1160 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1710841341
transform 1 0 1184 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1710841341
transform 1 0 1152 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1710841341
transform 1 0 744 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1710841341
transform 1 0 1456 0 1 1170
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1710841341
transform 1 0 408 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1710841341
transform 1 0 560 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1710841341
transform 1 0 536 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1710841341
transform 1 0 656 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1710841341
transform 1 0 256 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1710841341
transform 1 0 360 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1710841341
transform 1 0 256 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1710841341
transform 1 0 328 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1710841341
transform 1 0 576 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1710841341
transform 1 0 296 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1710841341
transform 1 0 392 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1710841341
transform 1 0 440 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1710841341
transform 1 0 456 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1710841341
transform 1 0 552 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1710841341
transform 1 0 72 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1710841341
transform 1 0 120 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1710841341
transform 1 0 360 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1710841341
transform 1 0 400 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1710841341
transform 1 0 480 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1710841341
transform 1 0 528 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1710841341
transform 1 0 656 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1710841341
transform 1 0 128 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1710841341
transform 1 0 112 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1710841341
transform 1 0 88 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1710841341
transform 1 0 280 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1710841341
transform 1 0 328 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1710841341
transform 1 0 648 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1710841341
transform 1 0 976 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1710841341
transform 1 0 160 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1710841341
transform 1 0 240 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1710841341
transform 1 0 728 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1710841341
transform 1 0 1056 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1710841341
transform 1 0 1624 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1710841341
transform 1 0 1832 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1710841341
transform 1 0 1992 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1710841341
transform 1 0 1840 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1710841341
transform 1 0 2440 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1710841341
transform 1 0 2408 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1710841341
transform 1 0 2472 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1710841341
transform 1 0 2576 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1710841341
transform 1 0 2576 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1710841341
transform 1 0 2576 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1710841341
transform 1 0 2576 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1710841341
transform 1 0 1920 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1710841341
transform 1 0 2576 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1710841341
transform 1 0 2576 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1710841341
transform 1 0 2408 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1710841341
transform 1 0 2056 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1710841341
transform 1 0 1616 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1710841341
transform 1 0 1432 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1710841341
transform 1 0 1096 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1710841341
transform 1 0 984 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1710841341
transform 1 0 816 0 1 2370
box -8 -3 104 105
use FILL  FILL_0
timestamp 1710841341
transform 1 0 2664 0 1 2370
box -8 -3 16 105
use FILL  FILL_1
timestamp 1710841341
transform 1 0 2656 0 1 2370
box -8 -3 16 105
use FILL  FILL_2
timestamp 1710841341
transform 1 0 2648 0 1 2370
box -8 -3 16 105
use FILL  FILL_3
timestamp 1710841341
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use FILL  FILL_4
timestamp 1710841341
transform 1 0 2592 0 1 2370
box -8 -3 16 105
use FILL  FILL_5
timestamp 1710841341
transform 1 0 2584 0 1 2370
box -8 -3 16 105
use FILL  FILL_6
timestamp 1710841341
transform 1 0 2576 0 1 2370
box -8 -3 16 105
use FILL  FILL_7
timestamp 1710841341
transform 1 0 2568 0 1 2370
box -8 -3 16 105
use FILL  FILL_8
timestamp 1710841341
transform 1 0 2512 0 1 2370
box -8 -3 16 105
use FILL  FILL_9
timestamp 1710841341
transform 1 0 2504 0 1 2370
box -8 -3 16 105
use FILL  FILL_10
timestamp 1710841341
transform 1 0 2400 0 1 2370
box -8 -3 16 105
use FILL  FILL_11
timestamp 1710841341
transform 1 0 2392 0 1 2370
box -8 -3 16 105
use FILL  FILL_12
timestamp 1710841341
transform 1 0 2352 0 1 2370
box -8 -3 16 105
use FILL  FILL_13
timestamp 1710841341
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use FILL  FILL_14
timestamp 1710841341
transform 1 0 2312 0 1 2370
box -8 -3 16 105
use FILL  FILL_15
timestamp 1710841341
transform 1 0 2304 0 1 2370
box -8 -3 16 105
use FILL  FILL_16
timestamp 1710841341
transform 1 0 2272 0 1 2370
box -8 -3 16 105
use FILL  FILL_17
timestamp 1710841341
transform 1 0 2264 0 1 2370
box -8 -3 16 105
use FILL  FILL_18
timestamp 1710841341
transform 1 0 2256 0 1 2370
box -8 -3 16 105
use FILL  FILL_19
timestamp 1710841341
transform 1 0 2208 0 1 2370
box -8 -3 16 105
use FILL  FILL_20
timestamp 1710841341
transform 1 0 2200 0 1 2370
box -8 -3 16 105
use FILL  FILL_21
timestamp 1710841341
transform 1 0 2168 0 1 2370
box -8 -3 16 105
use FILL  FILL_22
timestamp 1710841341
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_23
timestamp 1710841341
transform 1 0 2152 0 1 2370
box -8 -3 16 105
use FILL  FILL_24
timestamp 1710841341
transform 1 0 2048 0 1 2370
box -8 -3 16 105
use FILL  FILL_25
timestamp 1710841341
transform 1 0 2040 0 1 2370
box -8 -3 16 105
use FILL  FILL_26
timestamp 1710841341
transform 1 0 1976 0 1 2370
box -8 -3 16 105
use FILL  FILL_27
timestamp 1710841341
transform 1 0 1968 0 1 2370
box -8 -3 16 105
use FILL  FILL_28
timestamp 1710841341
transform 1 0 1960 0 1 2370
box -8 -3 16 105
use FILL  FILL_29
timestamp 1710841341
transform 1 0 1952 0 1 2370
box -8 -3 16 105
use FILL  FILL_30
timestamp 1710841341
transform 1 0 1920 0 1 2370
box -8 -3 16 105
use FILL  FILL_31
timestamp 1710841341
transform 1 0 1912 0 1 2370
box -8 -3 16 105
use FILL  FILL_32
timestamp 1710841341
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use FILL  FILL_33
timestamp 1710841341
transform 1 0 1856 0 1 2370
box -8 -3 16 105
use FILL  FILL_34
timestamp 1710841341
transform 1 0 1848 0 1 2370
box -8 -3 16 105
use FILL  FILL_35
timestamp 1710841341
transform 1 0 1816 0 1 2370
box -8 -3 16 105
use FILL  FILL_36
timestamp 1710841341
transform 1 0 1808 0 1 2370
box -8 -3 16 105
use FILL  FILL_37
timestamp 1710841341
transform 1 0 1776 0 1 2370
box -8 -3 16 105
use FILL  FILL_38
timestamp 1710841341
transform 1 0 1768 0 1 2370
box -8 -3 16 105
use FILL  FILL_39
timestamp 1710841341
transform 1 0 1760 0 1 2370
box -8 -3 16 105
use FILL  FILL_40
timestamp 1710841341
transform 1 0 1720 0 1 2370
box -8 -3 16 105
use FILL  FILL_41
timestamp 1710841341
transform 1 0 1712 0 1 2370
box -8 -3 16 105
use FILL  FILL_42
timestamp 1710841341
transform 1 0 1608 0 1 2370
box -8 -3 16 105
use FILL  FILL_43
timestamp 1710841341
transform 1 0 1600 0 1 2370
box -8 -3 16 105
use FILL  FILL_44
timestamp 1710841341
transform 1 0 1592 0 1 2370
box -8 -3 16 105
use FILL  FILL_45
timestamp 1710841341
transform 1 0 1552 0 1 2370
box -8 -3 16 105
use FILL  FILL_46
timestamp 1710841341
transform 1 0 1544 0 1 2370
box -8 -3 16 105
use FILL  FILL_47
timestamp 1710841341
transform 1 0 1536 0 1 2370
box -8 -3 16 105
use FILL  FILL_48
timestamp 1710841341
transform 1 0 1528 0 1 2370
box -8 -3 16 105
use FILL  FILL_49
timestamp 1710841341
transform 1 0 1424 0 1 2370
box -8 -3 16 105
use FILL  FILL_50
timestamp 1710841341
transform 1 0 1416 0 1 2370
box -8 -3 16 105
use FILL  FILL_51
timestamp 1710841341
transform 1 0 1376 0 1 2370
box -8 -3 16 105
use FILL  FILL_52
timestamp 1710841341
transform 1 0 1368 0 1 2370
box -8 -3 16 105
use FILL  FILL_53
timestamp 1710841341
transform 1 0 1360 0 1 2370
box -8 -3 16 105
use FILL  FILL_54
timestamp 1710841341
transform 1 0 1320 0 1 2370
box -8 -3 16 105
use FILL  FILL_55
timestamp 1710841341
transform 1 0 1312 0 1 2370
box -8 -3 16 105
use FILL  FILL_56
timestamp 1710841341
transform 1 0 1304 0 1 2370
box -8 -3 16 105
use FILL  FILL_57
timestamp 1710841341
transform 1 0 1296 0 1 2370
box -8 -3 16 105
use FILL  FILL_58
timestamp 1710841341
transform 1 0 1256 0 1 2370
box -8 -3 16 105
use FILL  FILL_59
timestamp 1710841341
transform 1 0 1248 0 1 2370
box -8 -3 16 105
use FILL  FILL_60
timestamp 1710841341
transform 1 0 1240 0 1 2370
box -8 -3 16 105
use FILL  FILL_61
timestamp 1710841341
transform 1 0 1200 0 1 2370
box -8 -3 16 105
use FILL  FILL_62
timestamp 1710841341
transform 1 0 1192 0 1 2370
box -8 -3 16 105
use FILL  FILL_63
timestamp 1710841341
transform 1 0 976 0 1 2370
box -8 -3 16 105
use FILL  FILL_64
timestamp 1710841341
transform 1 0 968 0 1 2370
box -8 -3 16 105
use FILL  FILL_65
timestamp 1710841341
transform 1 0 960 0 1 2370
box -8 -3 16 105
use FILL  FILL_66
timestamp 1710841341
transform 1 0 920 0 1 2370
box -8 -3 16 105
use FILL  FILL_67
timestamp 1710841341
transform 1 0 912 0 1 2370
box -8 -3 16 105
use FILL  FILL_68
timestamp 1710841341
transform 1 0 808 0 1 2370
box -8 -3 16 105
use FILL  FILL_69
timestamp 1710841341
transform 1 0 800 0 1 2370
box -8 -3 16 105
use FILL  FILL_70
timestamp 1710841341
transform 1 0 752 0 1 2370
box -8 -3 16 105
use FILL  FILL_71
timestamp 1710841341
transform 1 0 624 0 1 2370
box -8 -3 16 105
use FILL  FILL_72
timestamp 1710841341
transform 1 0 520 0 1 2370
box -8 -3 16 105
use FILL  FILL_73
timestamp 1710841341
transform 1 0 400 0 1 2370
box -8 -3 16 105
use FILL  FILL_74
timestamp 1710841341
transform 1 0 392 0 1 2370
box -8 -3 16 105
use FILL  FILL_75
timestamp 1710841341
transform 1 0 384 0 1 2370
box -8 -3 16 105
use FILL  FILL_76
timestamp 1710841341
transform 1 0 344 0 1 2370
box -8 -3 16 105
use FILL  FILL_77
timestamp 1710841341
transform 1 0 336 0 1 2370
box -8 -3 16 105
use FILL  FILL_78
timestamp 1710841341
transform 1 0 328 0 1 2370
box -8 -3 16 105
use FILL  FILL_79
timestamp 1710841341
transform 1 0 320 0 1 2370
box -8 -3 16 105
use FILL  FILL_80
timestamp 1710841341
transform 1 0 264 0 1 2370
box -8 -3 16 105
use FILL  FILL_81
timestamp 1710841341
transform 1 0 224 0 1 2370
box -8 -3 16 105
use FILL  FILL_82
timestamp 1710841341
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_83
timestamp 1710841341
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_84
timestamp 1710841341
transform 1 0 128 0 1 2370
box -8 -3 16 105
use FILL  FILL_85
timestamp 1710841341
transform 1 0 120 0 1 2370
box -8 -3 16 105
use FILL  FILL_86
timestamp 1710841341
transform 1 0 112 0 1 2370
box -8 -3 16 105
use FILL  FILL_87
timestamp 1710841341
transform 1 0 2664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_88
timestamp 1710841341
transform 1 0 2656 0 -1 2370
box -8 -3 16 105
use FILL  FILL_89
timestamp 1710841341
transform 1 0 2624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_90
timestamp 1710841341
transform 1 0 2616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_91
timestamp 1710841341
transform 1 0 2608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_92
timestamp 1710841341
transform 1 0 2600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_93
timestamp 1710841341
transform 1 0 2552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_94
timestamp 1710841341
transform 1 0 2544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_95
timestamp 1710841341
transform 1 0 2536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_96
timestamp 1710841341
transform 1 0 2528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_97
timestamp 1710841341
transform 1 0 2488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_98
timestamp 1710841341
transform 1 0 2480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_99
timestamp 1710841341
transform 1 0 2472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_100
timestamp 1710841341
transform 1 0 2464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_101
timestamp 1710841341
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_102
timestamp 1710841341
transform 1 0 2448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_103
timestamp 1710841341
transform 1 0 2440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_104
timestamp 1710841341
transform 1 0 2400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_105
timestamp 1710841341
transform 1 0 2392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_106
timestamp 1710841341
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_107
timestamp 1710841341
transform 1 0 2376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_108
timestamp 1710841341
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_109
timestamp 1710841341
transform 1 0 2320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_110
timestamp 1710841341
transform 1 0 2312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_111
timestamp 1710841341
transform 1 0 2304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_112
timestamp 1710841341
transform 1 0 2280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_113
timestamp 1710841341
transform 1 0 2240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_114
timestamp 1710841341
transform 1 0 2232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_115
timestamp 1710841341
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_116
timestamp 1710841341
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_117
timestamp 1710841341
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_118
timestamp 1710841341
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_119
timestamp 1710841341
transform 1 0 2136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_120
timestamp 1710841341
transform 1 0 2128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_121
timestamp 1710841341
transform 1 0 2120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_122
timestamp 1710841341
transform 1 0 2112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_123
timestamp 1710841341
transform 1 0 2072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_124
timestamp 1710841341
transform 1 0 2064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_125
timestamp 1710841341
transform 1 0 2056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_126
timestamp 1710841341
transform 1 0 2048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_127
timestamp 1710841341
transform 1 0 2000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_128
timestamp 1710841341
transform 1 0 1992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_129
timestamp 1710841341
transform 1 0 1984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_130
timestamp 1710841341
transform 1 0 1976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_131
timestamp 1710841341
transform 1 0 1936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_132
timestamp 1710841341
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_133
timestamp 1710841341
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_134
timestamp 1710841341
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_135
timestamp 1710841341
transform 1 0 1888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_136
timestamp 1710841341
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_137
timestamp 1710841341
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_138
timestamp 1710841341
transform 1 0 1808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_139
timestamp 1710841341
transform 1 0 1800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_140
timestamp 1710841341
transform 1 0 1792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_141
timestamp 1710841341
transform 1 0 1784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_142
timestamp 1710841341
transform 1 0 1752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_143
timestamp 1710841341
transform 1 0 1720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_144
timestamp 1710841341
transform 1 0 1712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_145
timestamp 1710841341
transform 1 0 1704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_146
timestamp 1710841341
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_147
timestamp 1710841341
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_148
timestamp 1710841341
transform 1 0 1640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_149
timestamp 1710841341
transform 1 0 1632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_150
timestamp 1710841341
transform 1 0 1624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_151
timestamp 1710841341
transform 1 0 1600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_152
timestamp 1710841341
transform 1 0 1592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_153
timestamp 1710841341
transform 1 0 1544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_154
timestamp 1710841341
transform 1 0 1536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_155
timestamp 1710841341
transform 1 0 1528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_156
timestamp 1710841341
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_157
timestamp 1710841341
transform 1 0 1472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_158
timestamp 1710841341
transform 1 0 1464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_159
timestamp 1710841341
transform 1 0 1456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_160
timestamp 1710841341
transform 1 0 1448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_161
timestamp 1710841341
transform 1 0 1408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_162
timestamp 1710841341
transform 1 0 1368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_163
timestamp 1710841341
transform 1 0 1360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_164
timestamp 1710841341
transform 1 0 1352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_165
timestamp 1710841341
transform 1 0 1344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_166
timestamp 1710841341
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_167
timestamp 1710841341
transform 1 0 1296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_168
timestamp 1710841341
transform 1 0 1288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_169
timestamp 1710841341
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_170
timestamp 1710841341
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_171
timestamp 1710841341
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_172
timestamp 1710841341
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_173
timestamp 1710841341
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_174
timestamp 1710841341
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_175
timestamp 1710841341
transform 1 0 1136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_176
timestamp 1710841341
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_177
timestamp 1710841341
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_178
timestamp 1710841341
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_179
timestamp 1710841341
transform 1 0 1072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_180
timestamp 1710841341
transform 1 0 1064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_181
timestamp 1710841341
transform 1 0 1056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_182
timestamp 1710841341
transform 1 0 1048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_183
timestamp 1710841341
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_184
timestamp 1710841341
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_185
timestamp 1710841341
transform 1 0 992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_186
timestamp 1710841341
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_187
timestamp 1710841341
transform 1 0 944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_188
timestamp 1710841341
transform 1 0 936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_189
timestamp 1710841341
transform 1 0 928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_190
timestamp 1710841341
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_191
timestamp 1710841341
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_192
timestamp 1710841341
transform 1 0 872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_193
timestamp 1710841341
transform 1 0 832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_194
timestamp 1710841341
transform 1 0 824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_195
timestamp 1710841341
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_196
timestamp 1710841341
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_197
timestamp 1710841341
transform 1 0 752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_198
timestamp 1710841341
transform 1 0 552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_199
timestamp 1710841341
transform 1 0 544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_200
timestamp 1710841341
transform 1 0 536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_201
timestamp 1710841341
transform 1 0 472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_202
timestamp 1710841341
transform 1 0 464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_203
timestamp 1710841341
transform 1 0 456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_204
timestamp 1710841341
transform 1 0 432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_205
timestamp 1710841341
transform 1 0 392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_206
timestamp 1710841341
transform 1 0 384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_207
timestamp 1710841341
transform 1 0 376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_208
timestamp 1710841341
transform 1 0 336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_209
timestamp 1710841341
transform 1 0 312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_210
timestamp 1710841341
transform 1 0 304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_211
timestamp 1710841341
transform 1 0 296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_212
timestamp 1710841341
transform 1 0 272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_213
timestamp 1710841341
transform 1 0 264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_214
timestamp 1710841341
transform 1 0 224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_215
timestamp 1710841341
transform 1 0 216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_216
timestamp 1710841341
transform 1 0 208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_217
timestamp 1710841341
transform 1 0 200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_218
timestamp 1710841341
transform 1 0 192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_219
timestamp 1710841341
transform 1 0 160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_220
timestamp 1710841341
transform 1 0 152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_221
timestamp 1710841341
transform 1 0 144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_222
timestamp 1710841341
transform 1 0 136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_223
timestamp 1710841341
transform 1 0 128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_224
timestamp 1710841341
transform 1 0 104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_225
timestamp 1710841341
transform 1 0 96 0 -1 2370
box -8 -3 16 105
use FILL  FILL_226
timestamp 1710841341
transform 1 0 88 0 -1 2370
box -8 -3 16 105
use FILL  FILL_227
timestamp 1710841341
transform 1 0 80 0 -1 2370
box -8 -3 16 105
use FILL  FILL_228
timestamp 1710841341
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_229
timestamp 1710841341
transform 1 0 2664 0 1 2170
box -8 -3 16 105
use FILL  FILL_230
timestamp 1710841341
transform 1 0 2656 0 1 2170
box -8 -3 16 105
use FILL  FILL_231
timestamp 1710841341
transform 1 0 2648 0 1 2170
box -8 -3 16 105
use FILL  FILL_232
timestamp 1710841341
transform 1 0 2640 0 1 2170
box -8 -3 16 105
use FILL  FILL_233
timestamp 1710841341
transform 1 0 2632 0 1 2170
box -8 -3 16 105
use FILL  FILL_234
timestamp 1710841341
transform 1 0 2592 0 1 2170
box -8 -3 16 105
use FILL  FILL_235
timestamp 1710841341
transform 1 0 2584 0 1 2170
box -8 -3 16 105
use FILL  FILL_236
timestamp 1710841341
transform 1 0 2544 0 1 2170
box -8 -3 16 105
use FILL  FILL_237
timestamp 1710841341
transform 1 0 2536 0 1 2170
box -8 -3 16 105
use FILL  FILL_238
timestamp 1710841341
transform 1 0 2528 0 1 2170
box -8 -3 16 105
use FILL  FILL_239
timestamp 1710841341
transform 1 0 2488 0 1 2170
box -8 -3 16 105
use FILL  FILL_240
timestamp 1710841341
transform 1 0 2456 0 1 2170
box -8 -3 16 105
use FILL  FILL_241
timestamp 1710841341
transform 1 0 2448 0 1 2170
box -8 -3 16 105
use FILL  FILL_242
timestamp 1710841341
transform 1 0 2440 0 1 2170
box -8 -3 16 105
use FILL  FILL_243
timestamp 1710841341
transform 1 0 2408 0 1 2170
box -8 -3 16 105
use FILL  FILL_244
timestamp 1710841341
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_245
timestamp 1710841341
transform 1 0 2376 0 1 2170
box -8 -3 16 105
use FILL  FILL_246
timestamp 1710841341
transform 1 0 2368 0 1 2170
box -8 -3 16 105
use FILL  FILL_247
timestamp 1710841341
transform 1 0 2336 0 1 2170
box -8 -3 16 105
use FILL  FILL_248
timestamp 1710841341
transform 1 0 2312 0 1 2170
box -8 -3 16 105
use FILL  FILL_249
timestamp 1710841341
transform 1 0 2304 0 1 2170
box -8 -3 16 105
use FILL  FILL_250
timestamp 1710841341
transform 1 0 2296 0 1 2170
box -8 -3 16 105
use FILL  FILL_251
timestamp 1710841341
transform 1 0 2288 0 1 2170
box -8 -3 16 105
use FILL  FILL_252
timestamp 1710841341
transform 1 0 2256 0 1 2170
box -8 -3 16 105
use FILL  FILL_253
timestamp 1710841341
transform 1 0 2216 0 1 2170
box -8 -3 16 105
use FILL  FILL_254
timestamp 1710841341
transform 1 0 2208 0 1 2170
box -8 -3 16 105
use FILL  FILL_255
timestamp 1710841341
transform 1 0 2200 0 1 2170
box -8 -3 16 105
use FILL  FILL_256
timestamp 1710841341
transform 1 0 2192 0 1 2170
box -8 -3 16 105
use FILL  FILL_257
timestamp 1710841341
transform 1 0 2152 0 1 2170
box -8 -3 16 105
use FILL  FILL_258
timestamp 1710841341
transform 1 0 2144 0 1 2170
box -8 -3 16 105
use FILL  FILL_259
timestamp 1710841341
transform 1 0 2112 0 1 2170
box -8 -3 16 105
use FILL  FILL_260
timestamp 1710841341
transform 1 0 2088 0 1 2170
box -8 -3 16 105
use FILL  FILL_261
timestamp 1710841341
transform 1 0 2080 0 1 2170
box -8 -3 16 105
use FILL  FILL_262
timestamp 1710841341
transform 1 0 2072 0 1 2170
box -8 -3 16 105
use FILL  FILL_263
timestamp 1710841341
transform 1 0 2064 0 1 2170
box -8 -3 16 105
use FILL  FILL_264
timestamp 1710841341
transform 1 0 2056 0 1 2170
box -8 -3 16 105
use FILL  FILL_265
timestamp 1710841341
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use FILL  FILL_266
timestamp 1710841341
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_267
timestamp 1710841341
transform 1 0 1992 0 1 2170
box -8 -3 16 105
use FILL  FILL_268
timestamp 1710841341
transform 1 0 1952 0 1 2170
box -8 -3 16 105
use FILL  FILL_269
timestamp 1710841341
transform 1 0 1944 0 1 2170
box -8 -3 16 105
use FILL  FILL_270
timestamp 1710841341
transform 1 0 1912 0 1 2170
box -8 -3 16 105
use FILL  FILL_271
timestamp 1710841341
transform 1 0 1904 0 1 2170
box -8 -3 16 105
use FILL  FILL_272
timestamp 1710841341
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use FILL  FILL_273
timestamp 1710841341
transform 1 0 1856 0 1 2170
box -8 -3 16 105
use FILL  FILL_274
timestamp 1710841341
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use FILL  FILL_275
timestamp 1710841341
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_276
timestamp 1710841341
transform 1 0 1808 0 1 2170
box -8 -3 16 105
use FILL  FILL_277
timestamp 1710841341
transform 1 0 1800 0 1 2170
box -8 -3 16 105
use FILL  FILL_278
timestamp 1710841341
transform 1 0 1792 0 1 2170
box -8 -3 16 105
use FILL  FILL_279
timestamp 1710841341
transform 1 0 1744 0 1 2170
box -8 -3 16 105
use FILL  FILL_280
timestamp 1710841341
transform 1 0 1736 0 1 2170
box -8 -3 16 105
use FILL  FILL_281
timestamp 1710841341
transform 1 0 1728 0 1 2170
box -8 -3 16 105
use FILL  FILL_282
timestamp 1710841341
transform 1 0 1720 0 1 2170
box -8 -3 16 105
use FILL  FILL_283
timestamp 1710841341
transform 1 0 1680 0 1 2170
box -8 -3 16 105
use FILL  FILL_284
timestamp 1710841341
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use FILL  FILL_285
timestamp 1710841341
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use FILL  FILL_286
timestamp 1710841341
transform 1 0 1624 0 1 2170
box -8 -3 16 105
use FILL  FILL_287
timestamp 1710841341
transform 1 0 1616 0 1 2170
box -8 -3 16 105
use FILL  FILL_288
timestamp 1710841341
transform 1 0 1608 0 1 2170
box -8 -3 16 105
use FILL  FILL_289
timestamp 1710841341
transform 1 0 1568 0 1 2170
box -8 -3 16 105
use FILL  FILL_290
timestamp 1710841341
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use FILL  FILL_291
timestamp 1710841341
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_292
timestamp 1710841341
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use FILL  FILL_293
timestamp 1710841341
transform 1 0 1504 0 1 2170
box -8 -3 16 105
use FILL  FILL_294
timestamp 1710841341
transform 1 0 1496 0 1 2170
box -8 -3 16 105
use FILL  FILL_295
timestamp 1710841341
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_296
timestamp 1710841341
transform 1 0 1440 0 1 2170
box -8 -3 16 105
use FILL  FILL_297
timestamp 1710841341
transform 1 0 1432 0 1 2170
box -8 -3 16 105
use FILL  FILL_298
timestamp 1710841341
transform 1 0 1424 0 1 2170
box -8 -3 16 105
use FILL  FILL_299
timestamp 1710841341
transform 1 0 1416 0 1 2170
box -8 -3 16 105
use FILL  FILL_300
timestamp 1710841341
transform 1 0 1408 0 1 2170
box -8 -3 16 105
use FILL  FILL_301
timestamp 1710841341
transform 1 0 1360 0 1 2170
box -8 -3 16 105
use FILL  FILL_302
timestamp 1710841341
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_303
timestamp 1710841341
transform 1 0 1344 0 1 2170
box -8 -3 16 105
use FILL  FILL_304
timestamp 1710841341
transform 1 0 1336 0 1 2170
box -8 -3 16 105
use FILL  FILL_305
timestamp 1710841341
transform 1 0 1296 0 1 2170
box -8 -3 16 105
use FILL  FILL_306
timestamp 1710841341
transform 1 0 1288 0 1 2170
box -8 -3 16 105
use FILL  FILL_307
timestamp 1710841341
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use FILL  FILL_308
timestamp 1710841341
transform 1 0 1240 0 1 2170
box -8 -3 16 105
use FILL  FILL_309
timestamp 1710841341
transform 1 0 1232 0 1 2170
box -8 -3 16 105
use FILL  FILL_310
timestamp 1710841341
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_311
timestamp 1710841341
transform 1 0 1184 0 1 2170
box -8 -3 16 105
use FILL  FILL_312
timestamp 1710841341
transform 1 0 1176 0 1 2170
box -8 -3 16 105
use FILL  FILL_313
timestamp 1710841341
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_314
timestamp 1710841341
transform 1 0 1128 0 1 2170
box -8 -3 16 105
use FILL  FILL_315
timestamp 1710841341
transform 1 0 1120 0 1 2170
box -8 -3 16 105
use FILL  FILL_316
timestamp 1710841341
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_317
timestamp 1710841341
transform 1 0 1072 0 1 2170
box -8 -3 16 105
use FILL  FILL_318
timestamp 1710841341
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_319
timestamp 1710841341
transform 1 0 1040 0 1 2170
box -8 -3 16 105
use FILL  FILL_320
timestamp 1710841341
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use FILL  FILL_321
timestamp 1710841341
transform 1 0 992 0 1 2170
box -8 -3 16 105
use FILL  FILL_322
timestamp 1710841341
transform 1 0 984 0 1 2170
box -8 -3 16 105
use FILL  FILL_323
timestamp 1710841341
transform 1 0 976 0 1 2170
box -8 -3 16 105
use FILL  FILL_324
timestamp 1710841341
transform 1 0 968 0 1 2170
box -8 -3 16 105
use FILL  FILL_325
timestamp 1710841341
transform 1 0 928 0 1 2170
box -8 -3 16 105
use FILL  FILL_326
timestamp 1710841341
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_327
timestamp 1710841341
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_328
timestamp 1710841341
transform 1 0 872 0 1 2170
box -8 -3 16 105
use FILL  FILL_329
timestamp 1710841341
transform 1 0 864 0 1 2170
box -8 -3 16 105
use FILL  FILL_330
timestamp 1710841341
transform 1 0 856 0 1 2170
box -8 -3 16 105
use FILL  FILL_331
timestamp 1710841341
transform 1 0 848 0 1 2170
box -8 -3 16 105
use FILL  FILL_332
timestamp 1710841341
transform 1 0 840 0 1 2170
box -8 -3 16 105
use FILL  FILL_333
timestamp 1710841341
transform 1 0 784 0 1 2170
box -8 -3 16 105
use FILL  FILL_334
timestamp 1710841341
transform 1 0 776 0 1 2170
box -8 -3 16 105
use FILL  FILL_335
timestamp 1710841341
transform 1 0 768 0 1 2170
box -8 -3 16 105
use FILL  FILL_336
timestamp 1710841341
transform 1 0 760 0 1 2170
box -8 -3 16 105
use FILL  FILL_337
timestamp 1710841341
transform 1 0 736 0 1 2170
box -8 -3 16 105
use FILL  FILL_338
timestamp 1710841341
transform 1 0 728 0 1 2170
box -8 -3 16 105
use FILL  FILL_339
timestamp 1710841341
transform 1 0 720 0 1 2170
box -8 -3 16 105
use FILL  FILL_340
timestamp 1710841341
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_341
timestamp 1710841341
transform 1 0 672 0 1 2170
box -8 -3 16 105
use FILL  FILL_342
timestamp 1710841341
transform 1 0 664 0 1 2170
box -8 -3 16 105
use FILL  FILL_343
timestamp 1710841341
transform 1 0 656 0 1 2170
box -8 -3 16 105
use FILL  FILL_344
timestamp 1710841341
transform 1 0 648 0 1 2170
box -8 -3 16 105
use FILL  FILL_345
timestamp 1710841341
transform 1 0 640 0 1 2170
box -8 -3 16 105
use FILL  FILL_346
timestamp 1710841341
transform 1 0 632 0 1 2170
box -8 -3 16 105
use FILL  FILL_347
timestamp 1710841341
transform 1 0 528 0 1 2170
box -8 -3 16 105
use FILL  FILL_348
timestamp 1710841341
transform 1 0 472 0 1 2170
box -8 -3 16 105
use FILL  FILL_349
timestamp 1710841341
transform 1 0 464 0 1 2170
box -8 -3 16 105
use FILL  FILL_350
timestamp 1710841341
transform 1 0 456 0 1 2170
box -8 -3 16 105
use FILL  FILL_351
timestamp 1710841341
transform 1 0 408 0 1 2170
box -8 -3 16 105
use FILL  FILL_352
timestamp 1710841341
transform 1 0 400 0 1 2170
box -8 -3 16 105
use FILL  FILL_353
timestamp 1710841341
transform 1 0 344 0 1 2170
box -8 -3 16 105
use FILL  FILL_354
timestamp 1710841341
transform 1 0 336 0 1 2170
box -8 -3 16 105
use FILL  FILL_355
timestamp 1710841341
transform 1 0 296 0 1 2170
box -8 -3 16 105
use FILL  FILL_356
timestamp 1710841341
transform 1 0 288 0 1 2170
box -8 -3 16 105
use FILL  FILL_357
timestamp 1710841341
transform 1 0 232 0 1 2170
box -8 -3 16 105
use FILL  FILL_358
timestamp 1710841341
transform 1 0 144 0 1 2170
box -8 -3 16 105
use FILL  FILL_359
timestamp 1710841341
transform 1 0 136 0 1 2170
box -8 -3 16 105
use FILL  FILL_360
timestamp 1710841341
transform 1 0 128 0 1 2170
box -8 -3 16 105
use FILL  FILL_361
timestamp 1710841341
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_362
timestamp 1710841341
transform 1 0 2624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_363
timestamp 1710841341
transform 1 0 2616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_364
timestamp 1710841341
transform 1 0 2608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_365
timestamp 1710841341
transform 1 0 2584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_366
timestamp 1710841341
transform 1 0 2576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_367
timestamp 1710841341
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_368
timestamp 1710841341
transform 1 0 2512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_369
timestamp 1710841341
transform 1 0 2504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_370
timestamp 1710841341
transform 1 0 2496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_371
timestamp 1710841341
transform 1 0 2488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_372
timestamp 1710841341
transform 1 0 2440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_373
timestamp 1710841341
transform 1 0 2432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_374
timestamp 1710841341
transform 1 0 2424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_375
timestamp 1710841341
transform 1 0 2368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_376
timestamp 1710841341
transform 1 0 2360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_377
timestamp 1710841341
transform 1 0 2352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_378
timestamp 1710841341
transform 1 0 2320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_379
timestamp 1710841341
transform 1 0 2312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_380
timestamp 1710841341
transform 1 0 2264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_381
timestamp 1710841341
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_382
timestamp 1710841341
transform 1 0 2248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_383
timestamp 1710841341
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_384
timestamp 1710841341
transform 1 0 2208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_385
timestamp 1710841341
transform 1 0 2200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_386
timestamp 1710841341
transform 1 0 2160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_387
timestamp 1710841341
transform 1 0 2136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_388
timestamp 1710841341
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_389
timestamp 1710841341
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_390
timestamp 1710841341
transform 1 0 2072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_391
timestamp 1710841341
transform 1 0 2064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_392
timestamp 1710841341
transform 1 0 2032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_393
timestamp 1710841341
transform 1 0 2024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_394
timestamp 1710841341
transform 1 0 1992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_395
timestamp 1710841341
transform 1 0 1968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_396
timestamp 1710841341
transform 1 0 1960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_397
timestamp 1710841341
transform 1 0 1920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_398
timestamp 1710841341
transform 1 0 1912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_399
timestamp 1710841341
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_400
timestamp 1710841341
transform 1 0 1896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_401
timestamp 1710841341
transform 1 0 1848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_402
timestamp 1710841341
transform 1 0 1840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_403
timestamp 1710841341
transform 1 0 1808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_404
timestamp 1710841341
transform 1 0 1800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_405
timestamp 1710841341
transform 1 0 1792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_406
timestamp 1710841341
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_407
timestamp 1710841341
transform 1 0 1728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_408
timestamp 1710841341
transform 1 0 1720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_409
timestamp 1710841341
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_410
timestamp 1710841341
transform 1 0 1672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_411
timestamp 1710841341
transform 1 0 1632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_412
timestamp 1710841341
transform 1 0 1624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_413
timestamp 1710841341
transform 1 0 1616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_414
timestamp 1710841341
transform 1 0 1576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_415
timestamp 1710841341
transform 1 0 1568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_416
timestamp 1710841341
transform 1 0 1560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_417
timestamp 1710841341
transform 1 0 1512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_418
timestamp 1710841341
transform 1 0 1504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_419
timestamp 1710841341
transform 1 0 1496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_420
timestamp 1710841341
transform 1 0 1448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_421
timestamp 1710841341
transform 1 0 1400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_422
timestamp 1710841341
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_423
timestamp 1710841341
transform 1 0 1384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_424
timestamp 1710841341
transform 1 0 1344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_425
timestamp 1710841341
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_426
timestamp 1710841341
transform 1 0 1288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_427
timestamp 1710841341
transform 1 0 1280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_428
timestamp 1710841341
transform 1 0 1272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_429
timestamp 1710841341
transform 1 0 1224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_430
timestamp 1710841341
transform 1 0 1216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_431
timestamp 1710841341
transform 1 0 1208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_432
timestamp 1710841341
transform 1 0 1160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_433
timestamp 1710841341
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_434
timestamp 1710841341
transform 1 0 1120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_435
timestamp 1710841341
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_436
timestamp 1710841341
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_437
timestamp 1710841341
transform 1 0 1096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_438
timestamp 1710841341
transform 1 0 1088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_439
timestamp 1710841341
transform 1 0 1032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_440
timestamp 1710841341
transform 1 0 1024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_441
timestamp 1710841341
transform 1 0 1016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_442
timestamp 1710841341
transform 1 0 952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_443
timestamp 1710841341
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_444
timestamp 1710841341
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_445
timestamp 1710841341
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_446
timestamp 1710841341
transform 1 0 864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_447
timestamp 1710841341
transform 1 0 856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_448
timestamp 1710841341
transform 1 0 848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_449
timestamp 1710841341
transform 1 0 792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_450
timestamp 1710841341
transform 1 0 784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_451
timestamp 1710841341
transform 1 0 744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_452
timestamp 1710841341
transform 1 0 736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_453
timestamp 1710841341
transform 1 0 688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_454
timestamp 1710841341
transform 1 0 680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_455
timestamp 1710841341
transform 1 0 672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_456
timestamp 1710841341
transform 1 0 472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_457
timestamp 1710841341
transform 1 0 400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_458
timestamp 1710841341
transform 1 0 392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_459
timestamp 1710841341
transform 1 0 320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_460
timestamp 1710841341
transform 1 0 312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_461
timestamp 1710841341
transform 1 0 232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_462
timestamp 1710841341
transform 1 0 152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_463
timestamp 1710841341
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_464
timestamp 1710841341
transform 1 0 136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_465
timestamp 1710841341
transform 1 0 128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_466
timestamp 1710841341
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_467
timestamp 1710841341
transform 1 0 2568 0 1 1970
box -8 -3 16 105
use FILL  FILL_468
timestamp 1710841341
transform 1 0 2560 0 1 1970
box -8 -3 16 105
use FILL  FILL_469
timestamp 1710841341
transform 1 0 2528 0 1 1970
box -8 -3 16 105
use FILL  FILL_470
timestamp 1710841341
transform 1 0 2488 0 1 1970
box -8 -3 16 105
use FILL  FILL_471
timestamp 1710841341
transform 1 0 2480 0 1 1970
box -8 -3 16 105
use FILL  FILL_472
timestamp 1710841341
transform 1 0 2472 0 1 1970
box -8 -3 16 105
use FILL  FILL_473
timestamp 1710841341
transform 1 0 2464 0 1 1970
box -8 -3 16 105
use FILL  FILL_474
timestamp 1710841341
transform 1 0 2456 0 1 1970
box -8 -3 16 105
use FILL  FILL_475
timestamp 1710841341
transform 1 0 2408 0 1 1970
box -8 -3 16 105
use FILL  FILL_476
timestamp 1710841341
transform 1 0 2400 0 1 1970
box -8 -3 16 105
use FILL  FILL_477
timestamp 1710841341
transform 1 0 2392 0 1 1970
box -8 -3 16 105
use FILL  FILL_478
timestamp 1710841341
transform 1 0 2384 0 1 1970
box -8 -3 16 105
use FILL  FILL_479
timestamp 1710841341
transform 1 0 2376 0 1 1970
box -8 -3 16 105
use FILL  FILL_480
timestamp 1710841341
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use FILL  FILL_481
timestamp 1710841341
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_482
timestamp 1710841341
transform 1 0 2304 0 1 1970
box -8 -3 16 105
use FILL  FILL_483
timestamp 1710841341
transform 1 0 2280 0 1 1970
box -8 -3 16 105
use FILL  FILL_484
timestamp 1710841341
transform 1 0 2272 0 1 1970
box -8 -3 16 105
use FILL  FILL_485
timestamp 1710841341
transform 1 0 2240 0 1 1970
box -8 -3 16 105
use FILL  FILL_486
timestamp 1710841341
transform 1 0 2216 0 1 1970
box -8 -3 16 105
use FILL  FILL_487
timestamp 1710841341
transform 1 0 2208 0 1 1970
box -8 -3 16 105
use FILL  FILL_488
timestamp 1710841341
transform 1 0 2168 0 1 1970
box -8 -3 16 105
use FILL  FILL_489
timestamp 1710841341
transform 1 0 2160 0 1 1970
box -8 -3 16 105
use FILL  FILL_490
timestamp 1710841341
transform 1 0 2152 0 1 1970
box -8 -3 16 105
use FILL  FILL_491
timestamp 1710841341
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use FILL  FILL_492
timestamp 1710841341
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_493
timestamp 1710841341
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use FILL  FILL_494
timestamp 1710841341
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use FILL  FILL_495
timestamp 1710841341
transform 1 0 2032 0 1 1970
box -8 -3 16 105
use FILL  FILL_496
timestamp 1710841341
transform 1 0 2024 0 1 1970
box -8 -3 16 105
use FILL  FILL_497
timestamp 1710841341
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_498
timestamp 1710841341
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_499
timestamp 1710841341
transform 1 0 1984 0 1 1970
box -8 -3 16 105
use FILL  FILL_500
timestamp 1710841341
transform 1 0 1936 0 1 1970
box -8 -3 16 105
use FILL  FILL_501
timestamp 1710841341
transform 1 0 1928 0 1 1970
box -8 -3 16 105
use FILL  FILL_502
timestamp 1710841341
transform 1 0 1920 0 1 1970
box -8 -3 16 105
use FILL  FILL_503
timestamp 1710841341
transform 1 0 1896 0 1 1970
box -8 -3 16 105
use FILL  FILL_504
timestamp 1710841341
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use FILL  FILL_505
timestamp 1710841341
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_506
timestamp 1710841341
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_507
timestamp 1710841341
transform 1 0 1800 0 1 1970
box -8 -3 16 105
use FILL  FILL_508
timestamp 1710841341
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_509
timestamp 1710841341
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use FILL  FILL_510
timestamp 1710841341
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use FILL  FILL_511
timestamp 1710841341
transform 1 0 1752 0 1 1970
box -8 -3 16 105
use FILL  FILL_512
timestamp 1710841341
transform 1 0 1704 0 1 1970
box -8 -3 16 105
use FILL  FILL_513
timestamp 1710841341
transform 1 0 1696 0 1 1970
box -8 -3 16 105
use FILL  FILL_514
timestamp 1710841341
transform 1 0 1688 0 1 1970
box -8 -3 16 105
use FILL  FILL_515
timestamp 1710841341
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use FILL  FILL_516
timestamp 1710841341
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use FILL  FILL_517
timestamp 1710841341
transform 1 0 1624 0 1 1970
box -8 -3 16 105
use FILL  FILL_518
timestamp 1710841341
transform 1 0 1616 0 1 1970
box -8 -3 16 105
use FILL  FILL_519
timestamp 1710841341
transform 1 0 1608 0 1 1970
box -8 -3 16 105
use FILL  FILL_520
timestamp 1710841341
transform 1 0 1568 0 1 1970
box -8 -3 16 105
use FILL  FILL_521
timestamp 1710841341
transform 1 0 1528 0 1 1970
box -8 -3 16 105
use FILL  FILL_522
timestamp 1710841341
transform 1 0 1520 0 1 1970
box -8 -3 16 105
use FILL  FILL_523
timestamp 1710841341
transform 1 0 1512 0 1 1970
box -8 -3 16 105
use FILL  FILL_524
timestamp 1710841341
transform 1 0 1464 0 1 1970
box -8 -3 16 105
use FILL  FILL_525
timestamp 1710841341
transform 1 0 1456 0 1 1970
box -8 -3 16 105
use FILL  FILL_526
timestamp 1710841341
transform 1 0 1448 0 1 1970
box -8 -3 16 105
use FILL  FILL_527
timestamp 1710841341
transform 1 0 1440 0 1 1970
box -8 -3 16 105
use FILL  FILL_528
timestamp 1710841341
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_529
timestamp 1710841341
transform 1 0 1400 0 1 1970
box -8 -3 16 105
use FILL  FILL_530
timestamp 1710841341
transform 1 0 1368 0 1 1970
box -8 -3 16 105
use FILL  FILL_531
timestamp 1710841341
transform 1 0 1360 0 1 1970
box -8 -3 16 105
use FILL  FILL_532
timestamp 1710841341
transform 1 0 1336 0 1 1970
box -8 -3 16 105
use FILL  FILL_533
timestamp 1710841341
transform 1 0 1328 0 1 1970
box -8 -3 16 105
use FILL  FILL_534
timestamp 1710841341
transform 1 0 1296 0 1 1970
box -8 -3 16 105
use FILL  FILL_535
timestamp 1710841341
transform 1 0 1288 0 1 1970
box -8 -3 16 105
use FILL  FILL_536
timestamp 1710841341
transform 1 0 1280 0 1 1970
box -8 -3 16 105
use FILL  FILL_537
timestamp 1710841341
transform 1 0 1240 0 1 1970
box -8 -3 16 105
use FILL  FILL_538
timestamp 1710841341
transform 1 0 1232 0 1 1970
box -8 -3 16 105
use FILL  FILL_539
timestamp 1710841341
transform 1 0 1224 0 1 1970
box -8 -3 16 105
use FILL  FILL_540
timestamp 1710841341
transform 1 0 1216 0 1 1970
box -8 -3 16 105
use FILL  FILL_541
timestamp 1710841341
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_542
timestamp 1710841341
transform 1 0 1160 0 1 1970
box -8 -3 16 105
use FILL  FILL_543
timestamp 1710841341
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_544
timestamp 1710841341
transform 1 0 1112 0 1 1970
box -8 -3 16 105
use FILL  FILL_545
timestamp 1710841341
transform 1 0 1104 0 1 1970
box -8 -3 16 105
use FILL  FILL_546
timestamp 1710841341
transform 1 0 1056 0 1 1970
box -8 -3 16 105
use FILL  FILL_547
timestamp 1710841341
transform 1 0 1048 0 1 1970
box -8 -3 16 105
use FILL  FILL_548
timestamp 1710841341
transform 1 0 1040 0 1 1970
box -8 -3 16 105
use FILL  FILL_549
timestamp 1710841341
transform 1 0 992 0 1 1970
box -8 -3 16 105
use FILL  FILL_550
timestamp 1710841341
transform 1 0 984 0 1 1970
box -8 -3 16 105
use FILL  FILL_551
timestamp 1710841341
transform 1 0 976 0 1 1970
box -8 -3 16 105
use FILL  FILL_552
timestamp 1710841341
transform 1 0 968 0 1 1970
box -8 -3 16 105
use FILL  FILL_553
timestamp 1710841341
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_554
timestamp 1710841341
transform 1 0 912 0 1 1970
box -8 -3 16 105
use FILL  FILL_555
timestamp 1710841341
transform 1 0 872 0 1 1970
box -8 -3 16 105
use FILL  FILL_556
timestamp 1710841341
transform 1 0 864 0 1 1970
box -8 -3 16 105
use FILL  FILL_557
timestamp 1710841341
transform 1 0 856 0 1 1970
box -8 -3 16 105
use FILL  FILL_558
timestamp 1710841341
transform 1 0 848 0 1 1970
box -8 -3 16 105
use FILL  FILL_559
timestamp 1710841341
transform 1 0 800 0 1 1970
box -8 -3 16 105
use FILL  FILL_560
timestamp 1710841341
transform 1 0 792 0 1 1970
box -8 -3 16 105
use FILL  FILL_561
timestamp 1710841341
transform 1 0 744 0 1 1970
box -8 -3 16 105
use FILL  FILL_562
timestamp 1710841341
transform 1 0 736 0 1 1970
box -8 -3 16 105
use FILL  FILL_563
timestamp 1710841341
transform 1 0 728 0 1 1970
box -8 -3 16 105
use FILL  FILL_564
timestamp 1710841341
transform 1 0 656 0 1 1970
box -8 -3 16 105
use FILL  FILL_565
timestamp 1710841341
transform 1 0 648 0 1 1970
box -8 -3 16 105
use FILL  FILL_566
timestamp 1710841341
transform 1 0 608 0 1 1970
box -8 -3 16 105
use FILL  FILL_567
timestamp 1710841341
transform 1 0 600 0 1 1970
box -8 -3 16 105
use FILL  FILL_568
timestamp 1710841341
transform 1 0 592 0 1 1970
box -8 -3 16 105
use FILL  FILL_569
timestamp 1710841341
transform 1 0 568 0 1 1970
box -8 -3 16 105
use FILL  FILL_570
timestamp 1710841341
transform 1 0 560 0 1 1970
box -8 -3 16 105
use FILL  FILL_571
timestamp 1710841341
transform 1 0 504 0 1 1970
box -8 -3 16 105
use FILL  FILL_572
timestamp 1710841341
transform 1 0 496 0 1 1970
box -8 -3 16 105
use FILL  FILL_573
timestamp 1710841341
transform 1 0 392 0 1 1970
box -8 -3 16 105
use FILL  FILL_574
timestamp 1710841341
transform 1 0 384 0 1 1970
box -8 -3 16 105
use FILL  FILL_575
timestamp 1710841341
transform 1 0 376 0 1 1970
box -8 -3 16 105
use FILL  FILL_576
timestamp 1710841341
transform 1 0 368 0 1 1970
box -8 -3 16 105
use FILL  FILL_577
timestamp 1710841341
transform 1 0 312 0 1 1970
box -8 -3 16 105
use FILL  FILL_578
timestamp 1710841341
transform 1 0 304 0 1 1970
box -8 -3 16 105
use FILL  FILL_579
timestamp 1710841341
transform 1 0 296 0 1 1970
box -8 -3 16 105
use FILL  FILL_580
timestamp 1710841341
transform 1 0 232 0 1 1970
box -8 -3 16 105
use FILL  FILL_581
timestamp 1710841341
transform 1 0 224 0 1 1970
box -8 -3 16 105
use FILL  FILL_582
timestamp 1710841341
transform 1 0 216 0 1 1970
box -8 -3 16 105
use FILL  FILL_583
timestamp 1710841341
transform 1 0 152 0 1 1970
box -8 -3 16 105
use FILL  FILL_584
timestamp 1710841341
transform 1 0 2664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_585
timestamp 1710841341
transform 1 0 2656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_586
timestamp 1710841341
transform 1 0 2648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_587
timestamp 1710841341
transform 1 0 2640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_588
timestamp 1710841341
transform 1 0 2632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_589
timestamp 1710841341
transform 1 0 2624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_590
timestamp 1710841341
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_591
timestamp 1710841341
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_592
timestamp 1710841341
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_593
timestamp 1710841341
transform 1 0 2560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_594
timestamp 1710841341
transform 1 0 2552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_595
timestamp 1710841341
transform 1 0 2544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_596
timestamp 1710841341
transform 1 0 2536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_597
timestamp 1710841341
transform 1 0 2512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_598
timestamp 1710841341
transform 1 0 2504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_599
timestamp 1710841341
transform 1 0 2464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_600
timestamp 1710841341
transform 1 0 2456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_601
timestamp 1710841341
transform 1 0 2448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_602
timestamp 1710841341
transform 1 0 2440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_603
timestamp 1710841341
transform 1 0 2408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_604
timestamp 1710841341
transform 1 0 2400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_605
timestamp 1710841341
transform 1 0 2392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_606
timestamp 1710841341
transform 1 0 2384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_607
timestamp 1710841341
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_608
timestamp 1710841341
transform 1 0 2328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_609
timestamp 1710841341
transform 1 0 2320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_610
timestamp 1710841341
transform 1 0 2312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_611
timestamp 1710841341
transform 1 0 2288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_612
timestamp 1710841341
transform 1 0 2280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_613
timestamp 1710841341
transform 1 0 2232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_614
timestamp 1710841341
transform 1 0 2224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_615
timestamp 1710841341
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_616
timestamp 1710841341
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_617
timestamp 1710841341
transform 1 0 2184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_618
timestamp 1710841341
transform 1 0 2176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_619
timestamp 1710841341
transform 1 0 2168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_620
timestamp 1710841341
transform 1 0 2128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_621
timestamp 1710841341
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_622
timestamp 1710841341
transform 1 0 2112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_623
timestamp 1710841341
transform 1 0 2104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_624
timestamp 1710841341
transform 1 0 2096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_625
timestamp 1710841341
transform 1 0 2072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_626
timestamp 1710841341
transform 1 0 2032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_627
timestamp 1710841341
transform 1 0 2024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_628
timestamp 1710841341
transform 1 0 2016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_629
timestamp 1710841341
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_630
timestamp 1710841341
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_631
timestamp 1710841341
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_632
timestamp 1710841341
transform 1 0 1856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_633
timestamp 1710841341
transform 1 0 1824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_634
timestamp 1710841341
transform 1 0 1816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_635
timestamp 1710841341
transform 1 0 1768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_636
timestamp 1710841341
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_637
timestamp 1710841341
transform 1 0 1752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_638
timestamp 1710841341
transform 1 0 1744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_639
timestamp 1710841341
transform 1 0 1696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_640
timestamp 1710841341
transform 1 0 1688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_641
timestamp 1710841341
transform 1 0 1680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_642
timestamp 1710841341
transform 1 0 1640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_643
timestamp 1710841341
transform 1 0 1632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_644
timestamp 1710841341
transform 1 0 1624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_645
timestamp 1710841341
transform 1 0 1592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_646
timestamp 1710841341
transform 1 0 1584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_647
timestamp 1710841341
transform 1 0 1544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_648
timestamp 1710841341
transform 1 0 1504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_649
timestamp 1710841341
transform 1 0 1496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_650
timestamp 1710841341
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_651
timestamp 1710841341
transform 1 0 1464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_652
timestamp 1710841341
transform 1 0 1432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_653
timestamp 1710841341
transform 1 0 1424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_654
timestamp 1710841341
transform 1 0 1416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_655
timestamp 1710841341
transform 1 0 1376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_656
timestamp 1710841341
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_657
timestamp 1710841341
transform 1 0 1328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_658
timestamp 1710841341
transform 1 0 1320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_659
timestamp 1710841341
transform 1 0 1312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_660
timestamp 1710841341
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_661
timestamp 1710841341
transform 1 0 1240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_662
timestamp 1710841341
transform 1 0 1232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_663
timestamp 1710841341
transform 1 0 1224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_664
timestamp 1710841341
transform 1 0 1184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_665
timestamp 1710841341
transform 1 0 1176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_666
timestamp 1710841341
transform 1 0 1136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_667
timestamp 1710841341
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_668
timestamp 1710841341
transform 1 0 1088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_669
timestamp 1710841341
transform 1 0 1080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_670
timestamp 1710841341
transform 1 0 1072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_671
timestamp 1710841341
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_672
timestamp 1710841341
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_673
timestamp 1710841341
transform 1 0 984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_674
timestamp 1710841341
transform 1 0 976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_675
timestamp 1710841341
transform 1 0 968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_676
timestamp 1710841341
transform 1 0 928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_677
timestamp 1710841341
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_678
timestamp 1710841341
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_679
timestamp 1710841341
transform 1 0 880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_680
timestamp 1710841341
transform 1 0 840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_681
timestamp 1710841341
transform 1 0 832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_682
timestamp 1710841341
transform 1 0 792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_683
timestamp 1710841341
transform 1 0 784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_684
timestamp 1710841341
transform 1 0 776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_685
timestamp 1710841341
transform 1 0 712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_686
timestamp 1710841341
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_687
timestamp 1710841341
transform 1 0 648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_688
timestamp 1710841341
transform 1 0 320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_689
timestamp 1710841341
transform 1 0 312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_690
timestamp 1710841341
transform 1 0 304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_691
timestamp 1710841341
transform 1 0 248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_692
timestamp 1710841341
transform 1 0 2568 0 1 1770
box -8 -3 16 105
use FILL  FILL_693
timestamp 1710841341
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_694
timestamp 1710841341
transform 1 0 2496 0 1 1770
box -8 -3 16 105
use FILL  FILL_695
timestamp 1710841341
transform 1 0 2456 0 1 1770
box -8 -3 16 105
use FILL  FILL_696
timestamp 1710841341
transform 1 0 2416 0 1 1770
box -8 -3 16 105
use FILL  FILL_697
timestamp 1710841341
transform 1 0 2408 0 1 1770
box -8 -3 16 105
use FILL  FILL_698
timestamp 1710841341
transform 1 0 2400 0 1 1770
box -8 -3 16 105
use FILL  FILL_699
timestamp 1710841341
transform 1 0 2352 0 1 1770
box -8 -3 16 105
use FILL  FILL_700
timestamp 1710841341
transform 1 0 2280 0 1 1770
box -8 -3 16 105
use FILL  FILL_701
timestamp 1710841341
transform 1 0 2272 0 1 1770
box -8 -3 16 105
use FILL  FILL_702
timestamp 1710841341
transform 1 0 2264 0 1 1770
box -8 -3 16 105
use FILL  FILL_703
timestamp 1710841341
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_704
timestamp 1710841341
transform 1 0 2184 0 1 1770
box -8 -3 16 105
use FILL  FILL_705
timestamp 1710841341
transform 1 0 2128 0 1 1770
box -8 -3 16 105
use FILL  FILL_706
timestamp 1710841341
transform 1 0 2120 0 1 1770
box -8 -3 16 105
use FILL  FILL_707
timestamp 1710841341
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use FILL  FILL_708
timestamp 1710841341
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_709
timestamp 1710841341
transform 1 0 2016 0 1 1770
box -8 -3 16 105
use FILL  FILL_710
timestamp 1710841341
transform 1 0 2008 0 1 1770
box -8 -3 16 105
use FILL  FILL_711
timestamp 1710841341
transform 1 0 1960 0 1 1770
box -8 -3 16 105
use FILL  FILL_712
timestamp 1710841341
transform 1 0 1952 0 1 1770
box -8 -3 16 105
use FILL  FILL_713
timestamp 1710841341
transform 1 0 1944 0 1 1770
box -8 -3 16 105
use FILL  FILL_714
timestamp 1710841341
transform 1 0 1936 0 1 1770
box -8 -3 16 105
use FILL  FILL_715
timestamp 1710841341
transform 1 0 1896 0 1 1770
box -8 -3 16 105
use FILL  FILL_716
timestamp 1710841341
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_717
timestamp 1710841341
transform 1 0 1840 0 1 1770
box -8 -3 16 105
use FILL  FILL_718
timestamp 1710841341
transform 1 0 1832 0 1 1770
box -8 -3 16 105
use FILL  FILL_719
timestamp 1710841341
transform 1 0 1824 0 1 1770
box -8 -3 16 105
use FILL  FILL_720
timestamp 1710841341
transform 1 0 1776 0 1 1770
box -8 -3 16 105
use FILL  FILL_721
timestamp 1710841341
transform 1 0 1768 0 1 1770
box -8 -3 16 105
use FILL  FILL_722
timestamp 1710841341
transform 1 0 1760 0 1 1770
box -8 -3 16 105
use FILL  FILL_723
timestamp 1710841341
transform 1 0 1720 0 1 1770
box -8 -3 16 105
use FILL  FILL_724
timestamp 1710841341
transform 1 0 1712 0 1 1770
box -8 -3 16 105
use FILL  FILL_725
timestamp 1710841341
transform 1 0 1704 0 1 1770
box -8 -3 16 105
use FILL  FILL_726
timestamp 1710841341
transform 1 0 1656 0 1 1770
box -8 -3 16 105
use FILL  FILL_727
timestamp 1710841341
transform 1 0 1632 0 1 1770
box -8 -3 16 105
use FILL  FILL_728
timestamp 1710841341
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use FILL  FILL_729
timestamp 1710841341
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_730
timestamp 1710841341
transform 1 0 1568 0 1 1770
box -8 -3 16 105
use FILL  FILL_731
timestamp 1710841341
transform 1 0 1560 0 1 1770
box -8 -3 16 105
use FILL  FILL_732
timestamp 1710841341
transform 1 0 1520 0 1 1770
box -8 -3 16 105
use FILL  FILL_733
timestamp 1710841341
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_734
timestamp 1710841341
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_735
timestamp 1710841341
transform 1 0 1496 0 1 1770
box -8 -3 16 105
use FILL  FILL_736
timestamp 1710841341
transform 1 0 1448 0 1 1770
box -8 -3 16 105
use FILL  FILL_737
timestamp 1710841341
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use FILL  FILL_738
timestamp 1710841341
transform 1 0 1408 0 1 1770
box -8 -3 16 105
use FILL  FILL_739
timestamp 1710841341
transform 1 0 1400 0 1 1770
box -8 -3 16 105
use FILL  FILL_740
timestamp 1710841341
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use FILL  FILL_741
timestamp 1710841341
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use FILL  FILL_742
timestamp 1710841341
transform 1 0 1312 0 1 1770
box -8 -3 16 105
use FILL  FILL_743
timestamp 1710841341
transform 1 0 1304 0 1 1770
box -8 -3 16 105
use FILL  FILL_744
timestamp 1710841341
transform 1 0 1296 0 1 1770
box -8 -3 16 105
use FILL  FILL_745
timestamp 1710841341
transform 1 0 1248 0 1 1770
box -8 -3 16 105
use FILL  FILL_746
timestamp 1710841341
transform 1 0 1240 0 1 1770
box -8 -3 16 105
use FILL  FILL_747
timestamp 1710841341
transform 1 0 1216 0 1 1770
box -8 -3 16 105
use FILL  FILL_748
timestamp 1710841341
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_749
timestamp 1710841341
transform 1 0 1168 0 1 1770
box -8 -3 16 105
use FILL  FILL_750
timestamp 1710841341
transform 1 0 1160 0 1 1770
box -8 -3 16 105
use FILL  FILL_751
timestamp 1710841341
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use FILL  FILL_752
timestamp 1710841341
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_753
timestamp 1710841341
transform 1 0 1080 0 1 1770
box -8 -3 16 105
use FILL  FILL_754
timestamp 1710841341
transform 1 0 1072 0 1 1770
box -8 -3 16 105
use FILL  FILL_755
timestamp 1710841341
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_756
timestamp 1710841341
transform 1 0 1032 0 1 1770
box -8 -3 16 105
use FILL  FILL_757
timestamp 1710841341
transform 1 0 992 0 1 1770
box -8 -3 16 105
use FILL  FILL_758
timestamp 1710841341
transform 1 0 984 0 1 1770
box -8 -3 16 105
use FILL  FILL_759
timestamp 1710841341
transform 1 0 976 0 1 1770
box -8 -3 16 105
use FILL  FILL_760
timestamp 1710841341
transform 1 0 936 0 1 1770
box -8 -3 16 105
use FILL  FILL_761
timestamp 1710841341
transform 1 0 928 0 1 1770
box -8 -3 16 105
use FILL  FILL_762
timestamp 1710841341
transform 1 0 880 0 1 1770
box -8 -3 16 105
use FILL  FILL_763
timestamp 1710841341
transform 1 0 872 0 1 1770
box -8 -3 16 105
use FILL  FILL_764
timestamp 1710841341
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_765
timestamp 1710841341
transform 1 0 856 0 1 1770
box -8 -3 16 105
use FILL  FILL_766
timestamp 1710841341
transform 1 0 824 0 1 1770
box -8 -3 16 105
use FILL  FILL_767
timestamp 1710841341
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_768
timestamp 1710841341
transform 1 0 792 0 1 1770
box -8 -3 16 105
use FILL  FILL_769
timestamp 1710841341
transform 1 0 736 0 1 1770
box -8 -3 16 105
use FILL  FILL_770
timestamp 1710841341
transform 1 0 728 0 1 1770
box -8 -3 16 105
use FILL  FILL_771
timestamp 1710841341
transform 1 0 720 0 1 1770
box -8 -3 16 105
use FILL  FILL_772
timestamp 1710841341
transform 1 0 680 0 1 1770
box -8 -3 16 105
use FILL  FILL_773
timestamp 1710841341
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_774
timestamp 1710841341
transform 1 0 632 0 1 1770
box -8 -3 16 105
use FILL  FILL_775
timestamp 1710841341
transform 1 0 624 0 1 1770
box -8 -3 16 105
use FILL  FILL_776
timestamp 1710841341
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_777
timestamp 1710841341
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_778
timestamp 1710841341
transform 1 0 568 0 1 1770
box -8 -3 16 105
use FILL  FILL_779
timestamp 1710841341
transform 1 0 512 0 1 1770
box -8 -3 16 105
use FILL  FILL_780
timestamp 1710841341
transform 1 0 504 0 1 1770
box -8 -3 16 105
use FILL  FILL_781
timestamp 1710841341
transform 1 0 496 0 1 1770
box -8 -3 16 105
use FILL  FILL_782
timestamp 1710841341
transform 1 0 464 0 1 1770
box -8 -3 16 105
use FILL  FILL_783
timestamp 1710841341
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_784
timestamp 1710841341
transform 1 0 352 0 1 1770
box -8 -3 16 105
use FILL  FILL_785
timestamp 1710841341
transform 1 0 248 0 1 1770
box -8 -3 16 105
use FILL  FILL_786
timestamp 1710841341
transform 1 0 240 0 1 1770
box -8 -3 16 105
use FILL  FILL_787
timestamp 1710841341
transform 1 0 232 0 1 1770
box -8 -3 16 105
use FILL  FILL_788
timestamp 1710841341
transform 1 0 224 0 1 1770
box -8 -3 16 105
use FILL  FILL_789
timestamp 1710841341
transform 1 0 216 0 1 1770
box -8 -3 16 105
use FILL  FILL_790
timestamp 1710841341
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_791
timestamp 1710841341
transform 1 0 200 0 1 1770
box -8 -3 16 105
use FILL  FILL_792
timestamp 1710841341
transform 1 0 192 0 1 1770
box -8 -3 16 105
use FILL  FILL_793
timestamp 1710841341
transform 1 0 184 0 1 1770
box -8 -3 16 105
use FILL  FILL_794
timestamp 1710841341
transform 1 0 176 0 1 1770
box -8 -3 16 105
use FILL  FILL_795
timestamp 1710841341
transform 1 0 168 0 1 1770
box -8 -3 16 105
use FILL  FILL_796
timestamp 1710841341
transform 1 0 160 0 1 1770
box -8 -3 16 105
use FILL  FILL_797
timestamp 1710841341
transform 1 0 152 0 1 1770
box -8 -3 16 105
use FILL  FILL_798
timestamp 1710841341
transform 1 0 144 0 1 1770
box -8 -3 16 105
use FILL  FILL_799
timestamp 1710841341
transform 1 0 136 0 1 1770
box -8 -3 16 105
use FILL  FILL_800
timestamp 1710841341
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_801
timestamp 1710841341
transform 1 0 120 0 1 1770
box -8 -3 16 105
use FILL  FILL_802
timestamp 1710841341
transform 1 0 112 0 1 1770
box -8 -3 16 105
use FILL  FILL_803
timestamp 1710841341
transform 1 0 104 0 1 1770
box -8 -3 16 105
use FILL  FILL_804
timestamp 1710841341
transform 1 0 96 0 1 1770
box -8 -3 16 105
use FILL  FILL_805
timestamp 1710841341
transform 1 0 88 0 1 1770
box -8 -3 16 105
use FILL  FILL_806
timestamp 1710841341
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_807
timestamp 1710841341
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_808
timestamp 1710841341
transform 1 0 2664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_809
timestamp 1710841341
transform 1 0 2624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_810
timestamp 1710841341
transform 1 0 2616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_811
timestamp 1710841341
transform 1 0 2608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_812
timestamp 1710841341
transform 1 0 2576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_813
timestamp 1710841341
transform 1 0 2552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_814
timestamp 1710841341
transform 1 0 2544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_815
timestamp 1710841341
transform 1 0 2496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_816
timestamp 1710841341
transform 1 0 2488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_817
timestamp 1710841341
transform 1 0 2480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_818
timestamp 1710841341
transform 1 0 2448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_819
timestamp 1710841341
transform 1 0 2424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_820
timestamp 1710841341
transform 1 0 2416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_821
timestamp 1710841341
transform 1 0 2376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_822
timestamp 1710841341
transform 1 0 2368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_823
timestamp 1710841341
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_824
timestamp 1710841341
transform 1 0 2312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_825
timestamp 1710841341
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_826
timestamp 1710841341
transform 1 0 2264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_827
timestamp 1710841341
transform 1 0 2216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_828
timestamp 1710841341
transform 1 0 2208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_829
timestamp 1710841341
transform 1 0 2200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_830
timestamp 1710841341
transform 1 0 2160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_831
timestamp 1710841341
transform 1 0 2152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_832
timestamp 1710841341
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_833
timestamp 1710841341
transform 1 0 2104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_834
timestamp 1710841341
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_835
timestamp 1710841341
transform 1 0 2040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_836
timestamp 1710841341
transform 1 0 2032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_837
timestamp 1710841341
transform 1 0 2024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_838
timestamp 1710841341
transform 1 0 2016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_839
timestamp 1710841341
transform 1 0 1952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_840
timestamp 1710841341
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_841
timestamp 1710841341
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_842
timestamp 1710841341
transform 1 0 1896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_843
timestamp 1710841341
transform 1 0 1888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_844
timestamp 1710841341
transform 1 0 1848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_845
timestamp 1710841341
transform 1 0 1840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_846
timestamp 1710841341
transform 1 0 1832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_847
timestamp 1710841341
transform 1 0 1824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_848
timestamp 1710841341
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_849
timestamp 1710841341
transform 1 0 1760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_850
timestamp 1710841341
transform 1 0 1752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_851
timestamp 1710841341
transform 1 0 1744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_852
timestamp 1710841341
transform 1 0 1736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_853
timestamp 1710841341
transform 1 0 1680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_854
timestamp 1710841341
transform 1 0 1672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_855
timestamp 1710841341
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_856
timestamp 1710841341
transform 1 0 1656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_857
timestamp 1710841341
transform 1 0 1616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_858
timestamp 1710841341
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_859
timestamp 1710841341
transform 1 0 1576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_860
timestamp 1710841341
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_861
timestamp 1710841341
transform 1 0 1560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_862
timestamp 1710841341
transform 1 0 1528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_863
timestamp 1710841341
transform 1 0 1504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_864
timestamp 1710841341
transform 1 0 1496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_865
timestamp 1710841341
transform 1 0 1464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_866
timestamp 1710841341
transform 1 0 1456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_867
timestamp 1710841341
transform 1 0 1448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_868
timestamp 1710841341
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_869
timestamp 1710841341
transform 1 0 1400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_870
timestamp 1710841341
transform 1 0 1392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_871
timestamp 1710841341
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_872
timestamp 1710841341
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_873
timestamp 1710841341
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_874
timestamp 1710841341
transform 1 0 1304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_875
timestamp 1710841341
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_876
timestamp 1710841341
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_877
timestamp 1710841341
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_878
timestamp 1710841341
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_879
timestamp 1710841341
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_880
timestamp 1710841341
transform 1 0 1128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_881
timestamp 1710841341
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_882
timestamp 1710841341
transform 1 0 1088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_883
timestamp 1710841341
transform 1 0 1080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_884
timestamp 1710841341
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_885
timestamp 1710841341
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_886
timestamp 1710841341
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_887
timestamp 1710841341
transform 1 0 952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_888
timestamp 1710841341
transform 1 0 944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_889
timestamp 1710841341
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_890
timestamp 1710841341
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_891
timestamp 1710841341
transform 1 0 888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_892
timestamp 1710841341
transform 1 0 880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_893
timestamp 1710841341
transform 1 0 840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_894
timestamp 1710841341
transform 1 0 832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_895
timestamp 1710841341
transform 1 0 824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_896
timestamp 1710841341
transform 1 0 776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_897
timestamp 1710841341
transform 1 0 768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_898
timestamp 1710841341
transform 1 0 760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_899
timestamp 1710841341
transform 1 0 752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_900
timestamp 1710841341
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_901
timestamp 1710841341
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_902
timestamp 1710841341
transform 1 0 680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_903
timestamp 1710841341
transform 1 0 640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_904
timestamp 1710841341
transform 1 0 632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_905
timestamp 1710841341
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_906
timestamp 1710841341
transform 1 0 584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_907
timestamp 1710841341
transform 1 0 576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_908
timestamp 1710841341
transform 1 0 536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_909
timestamp 1710841341
transform 1 0 432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_910
timestamp 1710841341
transform 1 0 424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_911
timestamp 1710841341
transform 1 0 416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_912
timestamp 1710841341
transform 1 0 408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_913
timestamp 1710841341
transform 1 0 400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_914
timestamp 1710841341
transform 1 0 392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_915
timestamp 1710841341
transform 1 0 368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_916
timestamp 1710841341
transform 1 0 328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_917
timestamp 1710841341
transform 1 0 320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_918
timestamp 1710841341
transform 1 0 312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_919
timestamp 1710841341
transform 1 0 304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_920
timestamp 1710841341
transform 1 0 296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_921
timestamp 1710841341
transform 1 0 232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_922
timestamp 1710841341
transform 1 0 224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_923
timestamp 1710841341
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_924
timestamp 1710841341
transform 1 0 2568 0 1 1570
box -8 -3 16 105
use FILL  FILL_925
timestamp 1710841341
transform 1 0 2560 0 1 1570
box -8 -3 16 105
use FILL  FILL_926
timestamp 1710841341
transform 1 0 2552 0 1 1570
box -8 -3 16 105
use FILL  FILL_927
timestamp 1710841341
transform 1 0 2528 0 1 1570
box -8 -3 16 105
use FILL  FILL_928
timestamp 1710841341
transform 1 0 2520 0 1 1570
box -8 -3 16 105
use FILL  FILL_929
timestamp 1710841341
transform 1 0 2472 0 1 1570
box -8 -3 16 105
use FILL  FILL_930
timestamp 1710841341
transform 1 0 2464 0 1 1570
box -8 -3 16 105
use FILL  FILL_931
timestamp 1710841341
transform 1 0 2456 0 1 1570
box -8 -3 16 105
use FILL  FILL_932
timestamp 1710841341
transform 1 0 2448 0 1 1570
box -8 -3 16 105
use FILL  FILL_933
timestamp 1710841341
transform 1 0 2424 0 1 1570
box -8 -3 16 105
use FILL  FILL_934
timestamp 1710841341
transform 1 0 2400 0 1 1570
box -8 -3 16 105
use FILL  FILL_935
timestamp 1710841341
transform 1 0 2392 0 1 1570
box -8 -3 16 105
use FILL  FILL_936
timestamp 1710841341
transform 1 0 2384 0 1 1570
box -8 -3 16 105
use FILL  FILL_937
timestamp 1710841341
transform 1 0 2376 0 1 1570
box -8 -3 16 105
use FILL  FILL_938
timestamp 1710841341
transform 1 0 2336 0 1 1570
box -8 -3 16 105
use FILL  FILL_939
timestamp 1710841341
transform 1 0 2328 0 1 1570
box -8 -3 16 105
use FILL  FILL_940
timestamp 1710841341
transform 1 0 2320 0 1 1570
box -8 -3 16 105
use FILL  FILL_941
timestamp 1710841341
transform 1 0 2312 0 1 1570
box -8 -3 16 105
use FILL  FILL_942
timestamp 1710841341
transform 1 0 2280 0 1 1570
box -8 -3 16 105
use FILL  FILL_943
timestamp 1710841341
transform 1 0 2256 0 1 1570
box -8 -3 16 105
use FILL  FILL_944
timestamp 1710841341
transform 1 0 2248 0 1 1570
box -8 -3 16 105
use FILL  FILL_945
timestamp 1710841341
transform 1 0 2240 0 1 1570
box -8 -3 16 105
use FILL  FILL_946
timestamp 1710841341
transform 1 0 2208 0 1 1570
box -8 -3 16 105
use FILL  FILL_947
timestamp 1710841341
transform 1 0 2200 0 1 1570
box -8 -3 16 105
use FILL  FILL_948
timestamp 1710841341
transform 1 0 2192 0 1 1570
box -8 -3 16 105
use FILL  FILL_949
timestamp 1710841341
transform 1 0 2184 0 1 1570
box -8 -3 16 105
use FILL  FILL_950
timestamp 1710841341
transform 1 0 2144 0 1 1570
box -8 -3 16 105
use FILL  FILL_951
timestamp 1710841341
transform 1 0 2136 0 1 1570
box -8 -3 16 105
use FILL  FILL_952
timestamp 1710841341
transform 1 0 2128 0 1 1570
box -8 -3 16 105
use FILL  FILL_953
timestamp 1710841341
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_954
timestamp 1710841341
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_955
timestamp 1710841341
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_956
timestamp 1710841341
transform 1 0 2032 0 1 1570
box -8 -3 16 105
use FILL  FILL_957
timestamp 1710841341
transform 1 0 2024 0 1 1570
box -8 -3 16 105
use FILL  FILL_958
timestamp 1710841341
transform 1 0 1976 0 1 1570
box -8 -3 16 105
use FILL  FILL_959
timestamp 1710841341
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use FILL  FILL_960
timestamp 1710841341
transform 1 0 1960 0 1 1570
box -8 -3 16 105
use FILL  FILL_961
timestamp 1710841341
transform 1 0 1952 0 1 1570
box -8 -3 16 105
use FILL  FILL_962
timestamp 1710841341
transform 1 0 1912 0 1 1570
box -8 -3 16 105
use FILL  FILL_963
timestamp 1710841341
transform 1 0 1904 0 1 1570
box -8 -3 16 105
use FILL  FILL_964
timestamp 1710841341
transform 1 0 1896 0 1 1570
box -8 -3 16 105
use FILL  FILL_965
timestamp 1710841341
transform 1 0 1848 0 1 1570
box -8 -3 16 105
use FILL  FILL_966
timestamp 1710841341
transform 1 0 1840 0 1 1570
box -8 -3 16 105
use FILL  FILL_967
timestamp 1710841341
transform 1 0 1832 0 1 1570
box -8 -3 16 105
use FILL  FILL_968
timestamp 1710841341
transform 1 0 1824 0 1 1570
box -8 -3 16 105
use FILL  FILL_969
timestamp 1710841341
transform 1 0 1784 0 1 1570
box -8 -3 16 105
use FILL  FILL_970
timestamp 1710841341
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use FILL  FILL_971
timestamp 1710841341
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_972
timestamp 1710841341
transform 1 0 1736 0 1 1570
box -8 -3 16 105
use FILL  FILL_973
timestamp 1710841341
transform 1 0 1728 0 1 1570
box -8 -3 16 105
use FILL  FILL_974
timestamp 1710841341
transform 1 0 1688 0 1 1570
box -8 -3 16 105
use FILL  FILL_975
timestamp 1710841341
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use FILL  FILL_976
timestamp 1710841341
transform 1 0 1672 0 1 1570
box -8 -3 16 105
use FILL  FILL_977
timestamp 1710841341
transform 1 0 1664 0 1 1570
box -8 -3 16 105
use FILL  FILL_978
timestamp 1710841341
transform 1 0 1632 0 1 1570
box -8 -3 16 105
use FILL  FILL_979
timestamp 1710841341
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use FILL  FILL_980
timestamp 1710841341
transform 1 0 1616 0 1 1570
box -8 -3 16 105
use FILL  FILL_981
timestamp 1710841341
transform 1 0 1584 0 1 1570
box -8 -3 16 105
use FILL  FILL_982
timestamp 1710841341
transform 1 0 1576 0 1 1570
box -8 -3 16 105
use FILL  FILL_983
timestamp 1710841341
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use FILL  FILL_984
timestamp 1710841341
transform 1 0 1536 0 1 1570
box -8 -3 16 105
use FILL  FILL_985
timestamp 1710841341
transform 1 0 1528 0 1 1570
box -8 -3 16 105
use FILL  FILL_986
timestamp 1710841341
transform 1 0 1520 0 1 1570
box -8 -3 16 105
use FILL  FILL_987
timestamp 1710841341
transform 1 0 1496 0 1 1570
box -8 -3 16 105
use FILL  FILL_988
timestamp 1710841341
transform 1 0 1488 0 1 1570
box -8 -3 16 105
use FILL  FILL_989
timestamp 1710841341
transform 1 0 1448 0 1 1570
box -8 -3 16 105
use FILL  FILL_990
timestamp 1710841341
transform 1 0 1440 0 1 1570
box -8 -3 16 105
use FILL  FILL_991
timestamp 1710841341
transform 1 0 1432 0 1 1570
box -8 -3 16 105
use FILL  FILL_992
timestamp 1710841341
transform 1 0 1424 0 1 1570
box -8 -3 16 105
use FILL  FILL_993
timestamp 1710841341
transform 1 0 1416 0 1 1570
box -8 -3 16 105
use FILL  FILL_994
timestamp 1710841341
transform 1 0 1376 0 1 1570
box -8 -3 16 105
use FILL  FILL_995
timestamp 1710841341
transform 1 0 1368 0 1 1570
box -8 -3 16 105
use FILL  FILL_996
timestamp 1710841341
transform 1 0 1360 0 1 1570
box -8 -3 16 105
use FILL  FILL_997
timestamp 1710841341
transform 1 0 1320 0 1 1570
box -8 -3 16 105
use FILL  FILL_998
timestamp 1710841341
transform 1 0 1312 0 1 1570
box -8 -3 16 105
use FILL  FILL_999
timestamp 1710841341
transform 1 0 1304 0 1 1570
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1710841341
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1710841341
transform 1 0 1288 0 1 1570
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1710841341
transform 1 0 1256 0 1 1570
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1710841341
transform 1 0 1248 0 1 1570
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1710841341
transform 1 0 1240 0 1 1570
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1710841341
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1710841341
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1710841341
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1710841341
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1710841341
transform 1 0 1160 0 1 1570
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1710841341
transform 1 0 1152 0 1 1570
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1710841341
transform 1 0 1128 0 1 1570
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1710841341
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1710841341
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1710841341
transform 1 0 1104 0 1 1570
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1710841341
transform 1 0 1064 0 1 1570
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1710841341
transform 1 0 1056 0 1 1570
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1710841341
transform 1 0 1048 0 1 1570
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1710841341
transform 1 0 1040 0 1 1570
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1710841341
transform 1 0 1000 0 1 1570
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1710841341
transform 1 0 992 0 1 1570
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1710841341
transform 1 0 984 0 1 1570
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1710841341
transform 1 0 976 0 1 1570
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1710841341
transform 1 0 968 0 1 1570
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1710841341
transform 1 0 960 0 1 1570
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1710841341
transform 1 0 920 0 1 1570
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1710841341
transform 1 0 912 0 1 1570
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1710841341
transform 1 0 904 0 1 1570
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1710841341
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1710841341
transform 1 0 856 0 1 1570
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1710841341
transform 1 0 848 0 1 1570
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1710841341
transform 1 0 840 0 1 1570
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1710841341
transform 1 0 832 0 1 1570
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1710841341
transform 1 0 776 0 1 1570
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1710841341
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1710841341
transform 1 0 760 0 1 1570
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1710841341
transform 1 0 720 0 1 1570
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1710841341
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1710841341
transform 1 0 704 0 1 1570
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1710841341
transform 1 0 672 0 1 1570
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1710841341
transform 1 0 664 0 1 1570
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1710841341
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1710841341
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1710841341
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1710841341
transform 1 0 568 0 1 1570
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1710841341
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1710841341
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1710841341
transform 1 0 488 0 1 1570
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1710841341
transform 1 0 288 0 1 1570
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1710841341
transform 1 0 280 0 1 1570
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1710841341
transform 1 0 224 0 1 1570
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1710841341
transform 1 0 2664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1710841341
transform 1 0 2624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1710841341
transform 1 0 2616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1710841341
transform 1 0 2608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1710841341
transform 1 0 2600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1710841341
transform 1 0 2552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1710841341
transform 1 0 2544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1710841341
transform 1 0 2520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1710841341
transform 1 0 2512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1710841341
transform 1 0 2480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1710841341
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1710841341
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1710841341
transform 1 0 2416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1710841341
transform 1 0 2408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1710841341
transform 1 0 2336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1710841341
transform 1 0 2328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1710841341
transform 1 0 2320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1710841341
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1710841341
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1710841341
transform 1 0 2264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1710841341
transform 1 0 2208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1710841341
transform 1 0 2200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1710841341
transform 1 0 2192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1710841341
transform 1 0 2184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1710841341
transform 1 0 2144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1710841341
transform 1 0 2136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1710841341
transform 1 0 2080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1710841341
transform 1 0 2072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1710841341
transform 1 0 2024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1710841341
transform 1 0 2016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1710841341
transform 1 0 2008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1710841341
transform 1 0 1968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1710841341
transform 1 0 1960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1710841341
transform 1 0 1928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1710841341
transform 1 0 1920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1710841341
transform 1 0 1888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1710841341
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1710841341
transform 1 0 1872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1710841341
transform 1 0 1832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1710841341
transform 1 0 1824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1710841341
transform 1 0 1816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1710841341
transform 1 0 1792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1710841341
transform 1 0 1760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1710841341
transform 1 0 1752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1710841341
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1710841341
transform 1 0 1712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1710841341
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1710841341
transform 1 0 1696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1710841341
transform 1 0 1664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1710841341
transform 1 0 1656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1710841341
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1710841341
transform 1 0 1616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1710841341
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1710841341
transform 1 0 1576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1710841341
transform 1 0 1568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1710841341
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1710841341
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1710841341
transform 1 0 1520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1710841341
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1710841341
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1710841341
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1710841341
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1710841341
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1710841341
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1710841341
transform 1 0 1416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1710841341
transform 1 0 1408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1710841341
transform 1 0 1368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1710841341
transform 1 0 1360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1710841341
transform 1 0 1336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1710841341
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1710841341
transform 1 0 1320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1710841341
transform 1 0 1288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1710841341
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1710841341
transform 1 0 1248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1710841341
transform 1 0 1240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1710841341
transform 1 0 1232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1710841341
transform 1 0 1224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1710841341
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1710841341
transform 1 0 1168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1710841341
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1710841341
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1710841341
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1710841341
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1710841341
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1710841341
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1710841341
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1710841341
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1710841341
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1710841341
transform 1 0 1008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1710841341
transform 1 0 1000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1710841341
transform 1 0 968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1710841341
transform 1 0 960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1710841341
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1710841341
transform 1 0 904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1710841341
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1710841341
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1710841341
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1710841341
transform 1 0 848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1710841341
transform 1 0 840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1710841341
transform 1 0 808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1710841341
transform 1 0 800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1710841341
transform 1 0 792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1710841341
transform 1 0 784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1710841341
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1710841341
transform 1 0 736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1710841341
transform 1 0 712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1710841341
transform 1 0 704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1710841341
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1710841341
transform 1 0 640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1710841341
transform 1 0 632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1710841341
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1710841341
transform 1 0 536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1710841341
transform 1 0 528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1710841341
transform 1 0 520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1710841341
transform 1 0 512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1710841341
transform 1 0 464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1710841341
transform 1 0 456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1710841341
transform 1 0 352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1710841341
transform 1 0 248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1710841341
transform 1 0 216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1710841341
transform 1 0 112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1710841341
transform 1 0 104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1710841341
transform 1 0 96 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1710841341
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1710841341
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1710841341
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1710841341
transform 1 0 2568 0 1 1370
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1710841341
transform 1 0 2512 0 1 1370
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1710841341
transform 1 0 2504 0 1 1370
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1710841341
transform 1 0 2432 0 1 1370
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1710841341
transform 1 0 2424 0 1 1370
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1710841341
transform 1 0 2416 0 1 1370
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1710841341
transform 1 0 2336 0 1 1370
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1710841341
transform 1 0 2328 0 1 1370
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1710841341
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1710841341
transform 1 0 2272 0 1 1370
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1710841341
transform 1 0 2264 0 1 1370
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1710841341
transform 1 0 2232 0 1 1370
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1710841341
transform 1 0 2224 0 1 1370
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1710841341
transform 1 0 2184 0 1 1370
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1710841341
transform 1 0 2176 0 1 1370
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1710841341
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1710841341
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1710841341
transform 1 0 2120 0 1 1370
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1710841341
transform 1 0 2080 0 1 1370
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1710841341
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1710841341
transform 1 0 2064 0 1 1370
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1710841341
transform 1 0 2016 0 1 1370
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1710841341
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1710841341
transform 1 0 1984 0 1 1370
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1710841341
transform 1 0 1976 0 1 1370
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1710841341
transform 1 0 1936 0 1 1370
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1710841341
transform 1 0 1928 0 1 1370
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1710841341
transform 1 0 1888 0 1 1370
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1710841341
transform 1 0 1848 0 1 1370
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1710841341
transform 1 0 1840 0 1 1370
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1710841341
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1710841341
transform 1 0 1792 0 1 1370
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1710841341
transform 1 0 1784 0 1 1370
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1710841341
transform 1 0 1776 0 1 1370
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1710841341
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1710841341
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1710841341
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1710841341
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1710841341
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1710841341
transform 1 0 1656 0 1 1370
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1710841341
transform 1 0 1648 0 1 1370
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1710841341
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1710841341
transform 1 0 1608 0 1 1370
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1710841341
transform 1 0 1584 0 1 1370
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1710841341
transform 1 0 1576 0 1 1370
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1710841341
transform 1 0 1552 0 1 1370
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1710841341
transform 1 0 1544 0 1 1370
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1710841341
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1710841341
transform 1 0 1496 0 1 1370
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1710841341
transform 1 0 1456 0 1 1370
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1710841341
transform 1 0 1448 0 1 1370
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1710841341
transform 1 0 1440 0 1 1370
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1710841341
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1710841341
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1710841341
transform 1 0 1384 0 1 1370
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1710841341
transform 1 0 1376 0 1 1370
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1710841341
transform 1 0 1336 0 1 1370
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1710841341
transform 1 0 1328 0 1 1370
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1710841341
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1710841341
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1710841341
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1710841341
transform 1 0 1248 0 1 1370
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1710841341
transform 1 0 1240 0 1 1370
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1710841341
transform 1 0 1208 0 1 1370
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1710841341
transform 1 0 1200 0 1 1370
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1710841341
transform 1 0 1168 0 1 1370
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1710841341
transform 1 0 1160 0 1 1370
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1710841341
transform 1 0 1152 0 1 1370
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1710841341
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1710841341
transform 1 0 1112 0 1 1370
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1710841341
transform 1 0 1104 0 1 1370
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1710841341
transform 1 0 1096 0 1 1370
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1710841341
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1710841341
transform 1 0 1040 0 1 1370
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1710841341
transform 1 0 1032 0 1 1370
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1710841341
transform 1 0 1024 0 1 1370
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1710841341
transform 1 0 1016 0 1 1370
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1710841341
transform 1 0 1008 0 1 1370
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1710841341
transform 1 0 1000 0 1 1370
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1710841341
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1710841341
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1710841341
transform 1 0 944 0 1 1370
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1710841341
transform 1 0 936 0 1 1370
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1710841341
transform 1 0 928 0 1 1370
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1710841341
transform 1 0 920 0 1 1370
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1710841341
transform 1 0 880 0 1 1370
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1710841341
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1710841341
transform 1 0 864 0 1 1370
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1710841341
transform 1 0 832 0 1 1370
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1710841341
transform 1 0 824 0 1 1370
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1710841341
transform 1 0 816 0 1 1370
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1710841341
transform 1 0 808 0 1 1370
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1710841341
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1710841341
transform 1 0 752 0 1 1370
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1710841341
transform 1 0 744 0 1 1370
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1710841341
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1710841341
transform 1 0 728 0 1 1370
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1710841341
transform 1 0 688 0 1 1370
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1710841341
transform 1 0 680 0 1 1370
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1710841341
transform 1 0 656 0 1 1370
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1710841341
transform 1 0 648 0 1 1370
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1710841341
transform 1 0 640 0 1 1370
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1710841341
transform 1 0 608 0 1 1370
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1710841341
transform 1 0 600 0 1 1370
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1710841341
transform 1 0 568 0 1 1370
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1710841341
transform 1 0 560 0 1 1370
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1710841341
transform 1 0 552 0 1 1370
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1710841341
transform 1 0 528 0 1 1370
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1710841341
transform 1 0 496 0 1 1370
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1710841341
transform 1 0 488 0 1 1370
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1710841341
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1710841341
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1710841341
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1710841341
transform 1 0 416 0 1 1370
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1710841341
transform 1 0 408 0 1 1370
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1710841341
transform 1 0 400 0 1 1370
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1710841341
transform 1 0 392 0 1 1370
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1710841341
transform 1 0 296 0 1 1370
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1710841341
transform 1 0 288 0 1 1370
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1710841341
transform 1 0 280 0 1 1370
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1710841341
transform 1 0 192 0 1 1370
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1710841341
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1710841341
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1710841341
transform 1 0 168 0 1 1370
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1710841341
transform 1 0 2664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1710841341
transform 1 0 2656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1710841341
transform 1 0 2648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1710841341
transform 1 0 2640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1710841341
transform 1 0 2632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1710841341
transform 1 0 2624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1710841341
transform 1 0 2600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1710841341
transform 1 0 2592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1710841341
transform 1 0 2584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1710841341
transform 1 0 2576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1710841341
transform 1 0 2568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1710841341
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1710841341
transform 1 0 2552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1710841341
transform 1 0 2544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1710841341
transform 1 0 2536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1710841341
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1710841341
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1710841341
transform 1 0 2480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1710841341
transform 1 0 2472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1710841341
transform 1 0 2464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1710841341
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1710841341
transform 1 0 2448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1710841341
transform 1 0 2440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1710841341
transform 1 0 2432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1710841341
transform 1 0 2424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1710841341
transform 1 0 2384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1710841341
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1710841341
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1710841341
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1710841341
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1710841341
transform 1 0 2344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1710841341
transform 1 0 2288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1710841341
transform 1 0 2280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1710841341
transform 1 0 2272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1710841341
transform 1 0 2264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1710841341
transform 1 0 2256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1710841341
transform 1 0 2216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1710841341
transform 1 0 2192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1710841341
transform 1 0 2184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1710841341
transform 1 0 2176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1710841341
transform 1 0 2168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1710841341
transform 1 0 2160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1710841341
transform 1 0 2104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1710841341
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1710841341
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1710841341
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1710841341
transform 1 0 2032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1710841341
transform 1 0 2024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1710841341
transform 1 0 2016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1710841341
transform 1 0 1984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1710841341
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1710841341
transform 1 0 1944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1710841341
transform 1 0 1936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1710841341
transform 1 0 1928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1710841341
transform 1 0 1888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1710841341
transform 1 0 1880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1710841341
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1710841341
transform 1 0 1832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1710841341
transform 1 0 1824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1710841341
transform 1 0 1816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1710841341
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1710841341
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1710841341
transform 1 0 1768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1710841341
transform 1 0 1728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1710841341
transform 1 0 1720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1710841341
transform 1 0 1712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1710841341
transform 1 0 1704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1710841341
transform 1 0 1696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1710841341
transform 1 0 1688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1710841341
transform 1 0 1648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1710841341
transform 1 0 1640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1710841341
transform 1 0 1632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1710841341
transform 1 0 1624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1710841341
transform 1 0 1600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1710841341
transform 1 0 1592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1710841341
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1710841341
transform 1 0 1576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1710841341
transform 1 0 1536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1710841341
transform 1 0 1528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1710841341
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1710841341
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1710841341
transform 1 0 1504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1710841341
transform 1 0 1480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1710841341
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1710841341
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1710841341
transform 1 0 1432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1710841341
transform 1 0 1424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1710841341
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1710841341
transform 1 0 1392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1710841341
transform 1 0 1360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1710841341
transform 1 0 1352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1710841341
transform 1 0 1344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1710841341
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1710841341
transform 1 0 1280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1710841341
transform 1 0 1272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1710841341
transform 1 0 1240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1710841341
transform 1 0 1232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1710841341
transform 1 0 1224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1710841341
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1710841341
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1710841341
transform 1 0 1176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1710841341
transform 1 0 1144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1710841341
transform 1 0 1136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1710841341
transform 1 0 1128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1710841341
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1710841341
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1710841341
transform 1 0 1080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1710841341
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1710841341
transform 1 0 1048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1710841341
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1710841341
transform 1 0 1016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1710841341
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1710841341
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1710841341
transform 1 0 968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1710841341
transform 1 0 960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1710841341
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1710841341
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1710841341
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1710841341
transform 1 0 872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1710841341
transform 1 0 864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1710841341
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1710841341
transform 1 0 824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1710841341
transform 1 0 816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1710841341
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1710841341
transform 1 0 752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1710841341
transform 1 0 744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1710841341
transform 1 0 736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1710841341
transform 1 0 728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1710841341
transform 1 0 720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1710841341
transform 1 0 680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1710841341
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1710841341
transform 1 0 632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1710841341
transform 1 0 624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1710841341
transform 1 0 616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1710841341
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1710841341
transform 1 0 568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1710841341
transform 1 0 560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1710841341
transform 1 0 512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1710841341
transform 1 0 472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1710841341
transform 1 0 432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1710841341
transform 1 0 384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1710841341
transform 1 0 376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1710841341
transform 1 0 368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1710841341
transform 1 0 336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1710841341
transform 1 0 328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1710841341
transform 1 0 304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1710841341
transform 1 0 296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1710841341
transform 1 0 256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1710841341
transform 1 0 232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1710841341
transform 1 0 224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1710841341
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1710841341
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1710841341
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1710841341
transform 1 0 2568 0 1 1170
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1710841341
transform 1 0 2504 0 1 1170
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1710841341
transform 1 0 2496 0 1 1170
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1710841341
transform 1 0 2488 0 1 1170
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1710841341
transform 1 0 2408 0 1 1170
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1710841341
transform 1 0 2400 0 1 1170
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1710841341
transform 1 0 2392 0 1 1170
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1710841341
transform 1 0 2328 0 1 1170
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1710841341
transform 1 0 2320 0 1 1170
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1710841341
transform 1 0 2312 0 1 1170
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1710841341
transform 1 0 2272 0 1 1170
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1710841341
transform 1 0 2264 0 1 1170
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1710841341
transform 1 0 2232 0 1 1170
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1710841341
transform 1 0 2224 0 1 1170
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1710841341
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1710841341
transform 1 0 2136 0 1 1170
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1710841341
transform 1 0 2128 0 1 1170
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1710841341
transform 1 0 2120 0 1 1170
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1710841341
transform 1 0 2112 0 1 1170
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1710841341
transform 1 0 2072 0 1 1170
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1710841341
transform 1 0 2064 0 1 1170
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1710841341
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1710841341
transform 1 0 2016 0 1 1170
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1710841341
transform 1 0 2008 0 1 1170
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1710841341
transform 1 0 2000 0 1 1170
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1710841341
transform 1 0 1992 0 1 1170
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1710841341
transform 1 0 1960 0 1 1170
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1710841341
transform 1 0 1936 0 1 1170
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1710841341
transform 1 0 1928 0 1 1170
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1710841341
transform 1 0 1920 0 1 1170
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1710841341
transform 1 0 1888 0 1 1170
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1710841341
transform 1 0 1880 0 1 1170
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1710841341
transform 1 0 1872 0 1 1170
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1710841341
transform 1 0 1840 0 1 1170
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1710841341
transform 1 0 1832 0 1 1170
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1710841341
transform 1 0 1824 0 1 1170
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1710841341
transform 1 0 1816 0 1 1170
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1710841341
transform 1 0 1768 0 1 1170
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1710841341
transform 1 0 1760 0 1 1170
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1710841341
transform 1 0 1752 0 1 1170
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1710841341
transform 1 0 1744 0 1 1170
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1710841341
transform 1 0 1736 0 1 1170
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1710841341
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1710841341
transform 1 0 1688 0 1 1170
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1710841341
transform 1 0 1680 0 1 1170
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1710841341
transform 1 0 1672 0 1 1170
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1710841341
transform 1 0 1664 0 1 1170
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1710841341
transform 1 0 1632 0 1 1170
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1710841341
transform 1 0 1624 0 1 1170
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1710841341
transform 1 0 1616 0 1 1170
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1710841341
transform 1 0 1608 0 1 1170
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1710841341
transform 1 0 1600 0 1 1170
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1710841341
transform 1 0 1560 0 1 1170
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1710841341
transform 1 0 1552 0 1 1170
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1710841341
transform 1 0 1544 0 1 1170
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1710841341
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1710841341
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1710841341
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1710841341
transform 1 0 1488 0 1 1170
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1710841341
transform 1 0 1480 0 1 1170
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1710841341
transform 1 0 1448 0 1 1170
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1710841341
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1710841341
transform 1 0 1432 0 1 1170
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1710841341
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1710841341
transform 1 0 1416 0 1 1170
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1710841341
transform 1 0 1376 0 1 1170
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1710841341
transform 1 0 1368 0 1 1170
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1710841341
transform 1 0 1360 0 1 1170
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1710841341
transform 1 0 1352 0 1 1170
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1710841341
transform 1 0 1344 0 1 1170
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1710841341
transform 1 0 1336 0 1 1170
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1710841341
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1710841341
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1710841341
transform 1 0 1288 0 1 1170
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1710841341
transform 1 0 1280 0 1 1170
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1710841341
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1710841341
transform 1 0 1240 0 1 1170
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1710841341
transform 1 0 1232 0 1 1170
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1710841341
transform 1 0 1224 0 1 1170
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1710841341
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1710841341
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1710841341
transform 1 0 1176 0 1 1170
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1710841341
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1710841341
transform 1 0 1160 0 1 1170
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1710841341
transform 1 0 1128 0 1 1170
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1710841341
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1710841341
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1710841341
transform 1 0 1080 0 1 1170
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1710841341
transform 1 0 1072 0 1 1170
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1710841341
transform 1 0 1064 0 1 1170
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1710841341
transform 1 0 1056 0 1 1170
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1710841341
transform 1 0 1024 0 1 1170
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1710841341
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1710841341
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1710841341
transform 1 0 1000 0 1 1170
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1710841341
transform 1 0 992 0 1 1170
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1710841341
transform 1 0 960 0 1 1170
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1710841341
transform 1 0 952 0 1 1170
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1710841341
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1710841341
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1710841341
transform 1 0 904 0 1 1170
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1710841341
transform 1 0 896 0 1 1170
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1710841341
transform 1 0 888 0 1 1170
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1710841341
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1710841341
transform 1 0 832 0 1 1170
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1710841341
transform 1 0 824 0 1 1170
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1710841341
transform 1 0 816 0 1 1170
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1710841341
transform 1 0 808 0 1 1170
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1710841341
transform 1 0 768 0 1 1170
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1710841341
transform 1 0 760 0 1 1170
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1710841341
transform 1 0 736 0 1 1170
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1710841341
transform 1 0 728 0 1 1170
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1710841341
transform 1 0 720 0 1 1170
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1710841341
transform 1 0 680 0 1 1170
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1710841341
transform 1 0 672 0 1 1170
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1710841341
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1710841341
transform 1 0 640 0 1 1170
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1710841341
transform 1 0 632 0 1 1170
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1710841341
transform 1 0 624 0 1 1170
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1710841341
transform 1 0 560 0 1 1170
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1710841341
transform 1 0 552 0 1 1170
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1710841341
transform 1 0 544 0 1 1170
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1710841341
transform 1 0 536 0 1 1170
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1710841341
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1710841341
transform 1 0 480 0 1 1170
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1710841341
transform 1 0 472 0 1 1170
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1710841341
transform 1 0 464 0 1 1170
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1710841341
transform 1 0 456 0 1 1170
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1710841341
transform 1 0 400 0 1 1170
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1710841341
transform 1 0 392 0 1 1170
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1710841341
transform 1 0 384 0 1 1170
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1710841341
transform 1 0 344 0 1 1170
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1710841341
transform 1 0 336 0 1 1170
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1710841341
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1710841341
transform 1 0 320 0 1 1170
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1710841341
transform 1 0 312 0 1 1170
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1710841341
transform 1 0 264 0 1 1170
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1710841341
transform 1 0 256 0 1 1170
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1710841341
transform 1 0 248 0 1 1170
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1710841341
transform 1 0 240 0 1 1170
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1710841341
transform 1 0 232 0 1 1170
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1710841341
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1710841341
transform 1 0 184 0 1 1170
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1710841341
transform 1 0 176 0 1 1170
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1710841341
transform 1 0 168 0 1 1170
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1710841341
transform 1 0 160 0 1 1170
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1710841341
transform 1 0 152 0 1 1170
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1710841341
transform 1 0 144 0 1 1170
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1710841341
transform 1 0 136 0 1 1170
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1710841341
transform 1 0 96 0 1 1170
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1710841341
transform 1 0 88 0 1 1170
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1710841341
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1710841341
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1710841341
transform 1 0 2664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1710841341
transform 1 0 2640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1710841341
transform 1 0 2608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1710841341
transform 1 0 2600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1710841341
transform 1 0 2560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1710841341
transform 1 0 2552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1710841341
transform 1 0 2544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1710841341
transform 1 0 2488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1710841341
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1710841341
transform 1 0 2472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1710841341
transform 1 0 2448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1710841341
transform 1 0 2408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1710841341
transform 1 0 2400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1710841341
transform 1 0 2392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1710841341
transform 1 0 2360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1710841341
transform 1 0 2352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1710841341
transform 1 0 2312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1710841341
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1710841341
transform 1 0 2296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1710841341
transform 1 0 2248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1710841341
transform 1 0 2240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1710841341
transform 1 0 2232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1710841341
transform 1 0 2224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1710841341
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1710841341
transform 1 0 2168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1710841341
transform 1 0 2160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1710841341
transform 1 0 2152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1710841341
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1710841341
transform 1 0 2088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1710841341
transform 1 0 2080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1710841341
transform 1 0 2072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1710841341
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1710841341
transform 1 0 2056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1710841341
transform 1 0 2016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1710841341
transform 1 0 1992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1710841341
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1710841341
transform 1 0 1976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1710841341
transform 1 0 1968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1710841341
transform 1 0 1936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1710841341
transform 1 0 1928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1710841341
transform 1 0 1920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1710841341
transform 1 0 1888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1710841341
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1710841341
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1710841341
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1710841341
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1710841341
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1710841341
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1710841341
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1710841341
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1710841341
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1710841341
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1710841341
transform 1 0 1736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1710841341
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1710841341
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1710841341
transform 1 0 1688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1710841341
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1710841341
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1710841341
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1710841341
transform 1 0 1632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1710841341
transform 1 0 1624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1710841341
transform 1 0 1616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1710841341
transform 1 0 1576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1710841341
transform 1 0 1568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1710841341
transform 1 0 1560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1710841341
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1710841341
transform 1 0 1520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1710841341
transform 1 0 1512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1710841341
transform 1 0 1504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1710841341
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1710841341
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1710841341
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1710841341
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1710841341
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1710841341
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1710841341
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1710841341
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1710841341
transform 1 0 1392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1710841341
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1710841341
transform 1 0 1352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1710841341
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1710841341
transform 1 0 1336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1710841341
transform 1 0 1312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1710841341
transform 1 0 1304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1710841341
transform 1 0 1296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1710841341
transform 1 0 1288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1710841341
transform 1 0 1256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1710841341
transform 1 0 1248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1710841341
transform 1 0 1240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1710841341
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1710841341
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1710841341
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1710841341
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1710841341
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1710841341
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1710841341
transform 1 0 1136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1710841341
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1710841341
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1710841341
transform 1 0 1112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1710841341
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1710841341
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1710841341
transform 1 0 1064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1710841341
transform 1 0 1056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1710841341
transform 1 0 1048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1710841341
transform 1 0 1016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1710841341
transform 1 0 1008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1710841341
transform 1 0 1000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1710841341
transform 1 0 968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1710841341
transform 1 0 960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1710841341
transform 1 0 952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1710841341
transform 1 0 944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1710841341
transform 1 0 936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1710841341
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1710841341
transform 1 0 888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1710841341
transform 1 0 880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1710841341
transform 1 0 872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1710841341
transform 1 0 832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1710841341
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1710841341
transform 1 0 816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1710841341
transform 1 0 808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1710841341
transform 1 0 800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1710841341
transform 1 0 792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1710841341
transform 1 0 752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1710841341
transform 1 0 744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1710841341
transform 1 0 736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1710841341
transform 1 0 728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1710841341
transform 1 0 720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1710841341
transform 1 0 680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1710841341
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1710841341
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1710841341
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1710841341
transform 1 0 616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1710841341
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1710841341
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1710841341
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1710841341
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1710841341
transform 1 0 536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1710841341
transform 1 0 528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1710841341
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1710841341
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1710841341
transform 1 0 488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1710841341
transform 1 0 440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1710841341
transform 1 0 432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1710841341
transform 1 0 408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1710841341
transform 1 0 400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1710841341
transform 1 0 336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1710841341
transform 1 0 328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1710841341
transform 1 0 320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1710841341
transform 1 0 280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1710841341
transform 1 0 240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1710841341
transform 1 0 232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1710841341
transform 1 0 224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1710841341
transform 1 0 160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1710841341
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1710841341
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1710841341
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1710841341
transform 1 0 2624 0 1 970
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1710841341
transform 1 0 2616 0 1 970
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1710841341
transform 1 0 2576 0 1 970
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1710841341
transform 1 0 2568 0 1 970
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1710841341
transform 1 0 2560 0 1 970
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1710841341
transform 1 0 2512 0 1 970
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1710841341
transform 1 0 2504 0 1 970
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1710841341
transform 1 0 2456 0 1 970
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1710841341
transform 1 0 2448 0 1 970
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1710841341
transform 1 0 2440 0 1 970
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1710841341
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1710841341
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1710841341
transform 1 0 2360 0 1 970
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1710841341
transform 1 0 2320 0 1 970
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1710841341
transform 1 0 2312 0 1 970
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1710841341
transform 1 0 2304 0 1 970
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1710841341
transform 1 0 2264 0 1 970
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1710841341
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1710841341
transform 1 0 2224 0 1 970
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1710841341
transform 1 0 2176 0 1 970
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1710841341
transform 1 0 2168 0 1 970
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1710841341
transform 1 0 2128 0 1 970
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1710841341
transform 1 0 2120 0 1 970
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1710841341
transform 1 0 2112 0 1 970
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1710841341
transform 1 0 2072 0 1 970
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1710841341
transform 1 0 2064 0 1 970
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1710841341
transform 1 0 2016 0 1 970
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1710841341
transform 1 0 2008 0 1 970
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1710841341
transform 1 0 2000 0 1 970
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1710841341
transform 1 0 1992 0 1 970
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1710841341
transform 1 0 1936 0 1 970
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1710841341
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1710841341
transform 1 0 1920 0 1 970
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1710841341
transform 1 0 1912 0 1 970
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1710841341
transform 1 0 1904 0 1 970
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1710841341
transform 1 0 1896 0 1 970
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1710841341
transform 1 0 1848 0 1 970
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1710841341
transform 1 0 1840 0 1 970
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1710841341
transform 1 0 1832 0 1 970
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1710841341
transform 1 0 1824 0 1 970
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1710841341
transform 1 0 1776 0 1 970
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1710841341
transform 1 0 1768 0 1 970
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1710841341
transform 1 0 1760 0 1 970
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1710841341
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1710841341
transform 1 0 1680 0 1 970
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1710841341
transform 1 0 1672 0 1 970
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1710841341
transform 1 0 1640 0 1 970
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1710841341
transform 1 0 1632 0 1 970
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1710841341
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1710841341
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1710841341
transform 1 0 1584 0 1 970
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1710841341
transform 1 0 1576 0 1 970
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1710841341
transform 1 0 1568 0 1 970
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1710841341
transform 1 0 1560 0 1 970
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1710841341
transform 1 0 1552 0 1 970
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1710841341
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1710841341
transform 1 0 1512 0 1 970
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1710841341
transform 1 0 1504 0 1 970
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1710841341
transform 1 0 1496 0 1 970
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1710841341
transform 1 0 1488 0 1 970
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1710841341
transform 1 0 1456 0 1 970
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1710841341
transform 1 0 1448 0 1 970
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1710841341
transform 1 0 1440 0 1 970
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1710841341
transform 1 0 1432 0 1 970
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1710841341
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1710841341
transform 1 0 1392 0 1 970
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1710841341
transform 1 0 1384 0 1 970
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1710841341
transform 1 0 1376 0 1 970
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1710841341
transform 1 0 1368 0 1 970
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1710841341
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1710841341
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1710841341
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1710841341
transform 1 0 1288 0 1 970
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1710841341
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1710841341
transform 1 0 1272 0 1 970
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1710841341
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1710841341
transform 1 0 1256 0 1 970
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1710841341
transform 1 0 1224 0 1 970
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1710841341
transform 1 0 1216 0 1 970
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1710841341
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1710841341
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1710841341
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1710841341
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1710841341
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1710841341
transform 1 0 1088 0 1 970
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1710841341
transform 1 0 1080 0 1 970
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1710841341
transform 1 0 1072 0 1 970
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1710841341
transform 1 0 1064 0 1 970
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1710841341
transform 1 0 1024 0 1 970
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1710841341
transform 1 0 1016 0 1 970
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1710841341
transform 1 0 1008 0 1 970
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1710841341
transform 1 0 1000 0 1 970
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1710841341
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1710841341
transform 1 0 944 0 1 970
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1710841341
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1710841341
transform 1 0 928 0 1 970
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1710841341
transform 1 0 920 0 1 970
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1710841341
transform 1 0 912 0 1 970
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1710841341
transform 1 0 872 0 1 970
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1710841341
transform 1 0 864 0 1 970
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1710841341
transform 1 0 856 0 1 970
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1710841341
transform 1 0 848 0 1 970
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1710841341
transform 1 0 840 0 1 970
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1710841341
transform 1 0 792 0 1 970
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1710841341
transform 1 0 784 0 1 970
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1710841341
transform 1 0 776 0 1 970
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1710841341
transform 1 0 768 0 1 970
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1710841341
transform 1 0 760 0 1 970
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1710841341
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1710841341
transform 1 0 688 0 1 970
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1710841341
transform 1 0 680 0 1 970
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1710841341
transform 1 0 672 0 1 970
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1710841341
transform 1 0 664 0 1 970
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1710841341
transform 1 0 624 0 1 970
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1710841341
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1710841341
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1710841341
transform 1 0 568 0 1 970
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1710841341
transform 1 0 504 0 1 970
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1710841341
transform 1 0 496 0 1 970
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1710841341
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1710841341
transform 1 0 480 0 1 970
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1710841341
transform 1 0 472 0 1 970
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1710841341
transform 1 0 432 0 1 970
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1710841341
transform 1 0 392 0 1 970
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1710841341
transform 1 0 384 0 1 970
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1710841341
transform 1 0 376 0 1 970
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1710841341
transform 1 0 272 0 1 970
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1710841341
transform 1 0 264 0 1 970
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1710841341
transform 1 0 224 0 1 970
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1710841341
transform 1 0 216 0 1 970
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1710841341
transform 1 0 192 0 1 970
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1710841341
transform 1 0 184 0 1 970
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1710841341
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1710841341
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1710841341
transform 1 0 160 0 1 970
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1710841341
transform 1 0 152 0 1 970
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1710841341
transform 1 0 144 0 1 970
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1710841341
transform 1 0 136 0 1 970
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1710841341
transform 1 0 128 0 1 970
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1710841341
transform 1 0 120 0 1 970
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1710841341
transform 1 0 112 0 1 970
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1710841341
transform 1 0 104 0 1 970
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1710841341
transform 1 0 96 0 1 970
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1710841341
transform 1 0 88 0 1 970
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1710841341
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1710841341
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1710841341
transform 1 0 2664 0 -1 970
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1710841341
transform 1 0 2632 0 -1 970
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1710841341
transform 1 0 2624 0 -1 970
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1710841341
transform 1 0 2616 0 -1 970
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1710841341
transform 1 0 2592 0 -1 970
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1710841341
transform 1 0 2584 0 -1 970
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1710841341
transform 1 0 2544 0 -1 970
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1710841341
transform 1 0 2536 0 -1 970
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1710841341
transform 1 0 2432 0 -1 970
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1710841341
transform 1 0 2424 0 -1 970
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1710841341
transform 1 0 2384 0 -1 970
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1710841341
transform 1 0 2352 0 -1 970
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1710841341
transform 1 0 2344 0 -1 970
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1710841341
transform 1 0 2336 0 -1 970
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1710841341
transform 1 0 2328 0 -1 970
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1710841341
transform 1 0 2288 0 -1 970
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1710841341
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1710841341
transform 1 0 2256 0 -1 970
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1710841341
transform 1 0 2248 0 -1 970
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1710841341
transform 1 0 2200 0 -1 970
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1710841341
transform 1 0 2192 0 -1 970
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1710841341
transform 1 0 2184 0 -1 970
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1710841341
transform 1 0 2176 0 -1 970
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1710841341
transform 1 0 2136 0 -1 970
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1710841341
transform 1 0 2104 0 -1 970
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1710841341
transform 1 0 2096 0 -1 970
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1710841341
transform 1 0 2088 0 -1 970
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1710841341
transform 1 0 2080 0 -1 970
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1710841341
transform 1 0 2072 0 -1 970
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1710841341
transform 1 0 2024 0 -1 970
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1710841341
transform 1 0 2016 0 -1 970
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1710841341
transform 1 0 2008 0 -1 970
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1710841341
transform 1 0 1984 0 -1 970
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1710841341
transform 1 0 1952 0 -1 970
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1710841341
transform 1 0 1944 0 -1 970
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1710841341
transform 1 0 1936 0 -1 970
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1710841341
transform 1 0 1928 0 -1 970
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1710841341
transform 1 0 1880 0 -1 970
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1710841341
transform 1 0 1872 0 -1 970
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1710841341
transform 1 0 1864 0 -1 970
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1710841341
transform 1 0 1856 0 -1 970
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1710841341
transform 1 0 1808 0 -1 970
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1710841341
transform 1 0 1800 0 -1 970
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1710841341
transform 1 0 1792 0 -1 970
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1710841341
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1710841341
transform 1 0 1744 0 -1 970
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1710841341
transform 1 0 1736 0 -1 970
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1710841341
transform 1 0 1728 0 -1 970
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1710841341
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1710841341
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1710841341
transform 1 0 1672 0 -1 970
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1710841341
transform 1 0 1664 0 -1 970
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1710841341
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1710841341
transform 1 0 1616 0 -1 970
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1710841341
transform 1 0 1608 0 -1 970
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1710841341
transform 1 0 1600 0 -1 970
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1710841341
transform 1 0 1560 0 -1 970
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1710841341
transform 1 0 1552 0 -1 970
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1710841341
transform 1 0 1544 0 -1 970
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1710841341
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1710841341
transform 1 0 1512 0 -1 970
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1710841341
transform 1 0 1504 0 -1 970
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1710841341
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1710841341
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1710841341
transform 1 0 1448 0 -1 970
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1710841341
transform 1 0 1408 0 -1 970
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1710841341
transform 1 0 1400 0 -1 970
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1710841341
transform 1 0 1392 0 -1 970
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1710841341
transform 1 0 1384 0 -1 970
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1710841341
transform 1 0 1336 0 -1 970
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1710841341
transform 1 0 1328 0 -1 970
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1710841341
transform 1 0 1320 0 -1 970
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1710841341
transform 1 0 1272 0 -1 970
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1710841341
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1710841341
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1710841341
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1710841341
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1710841341
transform 1 0 1184 0 -1 970
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1710841341
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1710841341
transform 1 0 1168 0 -1 970
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1710841341
transform 1 0 1128 0 -1 970
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1710841341
transform 1 0 1120 0 -1 970
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1710841341
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1710841341
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1710841341
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1710841341
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1710841341
transform 1 0 1016 0 -1 970
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1710841341
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1710841341
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1710841341
transform 1 0 976 0 -1 970
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1710841341
transform 1 0 968 0 -1 970
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1710841341
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1710841341
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1710841341
transform 1 0 880 0 -1 970
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1710841341
transform 1 0 872 0 -1 970
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1710841341
transform 1 0 840 0 -1 970
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1710841341
transform 1 0 832 0 -1 970
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1710841341
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1710841341
transform 1 0 784 0 -1 970
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1710841341
transform 1 0 776 0 -1 970
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1710841341
transform 1 0 736 0 -1 970
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1710841341
transform 1 0 728 0 -1 970
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1710841341
transform 1 0 720 0 -1 970
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1710841341
transform 1 0 712 0 -1 970
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1710841341
transform 1 0 656 0 -1 970
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1710841341
transform 1 0 648 0 -1 970
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1710841341
transform 1 0 640 0 -1 970
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1710841341
transform 1 0 632 0 -1 970
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1710841341
transform 1 0 592 0 -1 970
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1710841341
transform 1 0 552 0 -1 970
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1710841341
transform 1 0 544 0 -1 970
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1710841341
transform 1 0 536 0 -1 970
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1710841341
transform 1 0 528 0 -1 970
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1710841341
transform 1 0 520 0 -1 970
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1710841341
transform 1 0 464 0 -1 970
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1710841341
transform 1 0 456 0 -1 970
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1710841341
transform 1 0 448 0 -1 970
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1710841341
transform 1 0 440 0 -1 970
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1710841341
transform 1 0 432 0 -1 970
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1710841341
transform 1 0 384 0 -1 970
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1710841341
transform 1 0 376 0 -1 970
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1710841341
transform 1 0 368 0 -1 970
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1710841341
transform 1 0 360 0 -1 970
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1710841341
transform 1 0 328 0 -1 970
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1710841341
transform 1 0 320 0 -1 970
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1710841341
transform 1 0 312 0 -1 970
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1710841341
transform 1 0 304 0 -1 970
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1710841341
transform 1 0 296 0 -1 970
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1710841341
transform 1 0 288 0 -1 970
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1710841341
transform 1 0 280 0 -1 970
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1710841341
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1710841341
transform 1 0 224 0 -1 970
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1710841341
transform 1 0 216 0 -1 970
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1710841341
transform 1 0 208 0 -1 970
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1710841341
transform 1 0 104 0 -1 970
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1710841341
transform 1 0 96 0 -1 970
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1710841341
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1710841341
transform 1 0 2664 0 1 770
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1710841341
transform 1 0 2656 0 1 770
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1710841341
transform 1 0 2608 0 1 770
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1710841341
transform 1 0 2600 0 1 770
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1710841341
transform 1 0 2592 0 1 770
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1710841341
transform 1 0 2584 0 1 770
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1710841341
transform 1 0 2552 0 1 770
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1710841341
transform 1 0 2544 0 1 770
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1710841341
transform 1 0 2504 0 1 770
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1710841341
transform 1 0 2496 0 1 770
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1710841341
transform 1 0 2488 0 1 770
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1710841341
transform 1 0 2480 0 1 770
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1710841341
transform 1 0 2448 0 1 770
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1710841341
transform 1 0 2440 0 1 770
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1710841341
transform 1 0 2432 0 1 770
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1710841341
transform 1 0 2392 0 1 770
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1710841341
transform 1 0 2384 0 1 770
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1710841341
transform 1 0 2376 0 1 770
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1710841341
transform 1 0 2368 0 1 770
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1710841341
transform 1 0 2344 0 1 770
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1710841341
transform 1 0 2336 0 1 770
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1710841341
transform 1 0 2312 0 1 770
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1710841341
transform 1 0 2304 0 1 770
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1710841341
transform 1 0 2296 0 1 770
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1710841341
transform 1 0 2256 0 1 770
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1710841341
transform 1 0 2248 0 1 770
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1710841341
transform 1 0 2240 0 1 770
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1710841341
transform 1 0 2208 0 1 770
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1710841341
transform 1 0 2200 0 1 770
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1710841341
transform 1 0 2192 0 1 770
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1710841341
transform 1 0 2152 0 1 770
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1710841341
transform 1 0 2144 0 1 770
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1710841341
transform 1 0 2104 0 1 770
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1710841341
transform 1 0 2096 0 1 770
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1710841341
transform 1 0 2088 0 1 770
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1710841341
transform 1 0 2080 0 1 770
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1710841341
transform 1 0 2032 0 1 770
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1710841341
transform 1 0 2024 0 1 770
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1710841341
transform 1 0 2016 0 1 770
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1710841341
transform 1 0 2008 0 1 770
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1710841341
transform 1 0 1968 0 1 770
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1710841341
transform 1 0 1960 0 1 770
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1710841341
transform 1 0 1928 0 1 770
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1710841341
transform 1 0 1920 0 1 770
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1710841341
transform 1 0 1912 0 1 770
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1710841341
transform 1 0 1904 0 1 770
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1710841341
transform 1 0 1864 0 1 770
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1710841341
transform 1 0 1856 0 1 770
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1710841341
transform 1 0 1848 0 1 770
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1710841341
transform 1 0 1840 0 1 770
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1710841341
transform 1 0 1808 0 1 770
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1710841341
transform 1 0 1800 0 1 770
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1710841341
transform 1 0 1776 0 1 770
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1710841341
transform 1 0 1768 0 1 770
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1710841341
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1710841341
transform 1 0 1720 0 1 770
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1710841341
transform 1 0 1712 0 1 770
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1710841341
transform 1 0 1704 0 1 770
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1710841341
transform 1 0 1696 0 1 770
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1710841341
transform 1 0 1672 0 1 770
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1710841341
transform 1 0 1664 0 1 770
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1710841341
transform 1 0 1656 0 1 770
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1710841341
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1710841341
transform 1 0 1608 0 1 770
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1710841341
transform 1 0 1600 0 1 770
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1710841341
transform 1 0 1592 0 1 770
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1710841341
transform 1 0 1584 0 1 770
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1710841341
transform 1 0 1560 0 1 770
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1710841341
transform 1 0 1552 0 1 770
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1710841341
transform 1 0 1520 0 1 770
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1710841341
transform 1 0 1512 0 1 770
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1710841341
transform 1 0 1504 0 1 770
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1710841341
transform 1 0 1480 0 1 770
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1710841341
transform 1 0 1472 0 1 770
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1710841341
transform 1 0 1464 0 1 770
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1710841341
transform 1 0 1456 0 1 770
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1710841341
transform 1 0 1408 0 1 770
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1710841341
transform 1 0 1400 0 1 770
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1710841341
transform 1 0 1392 0 1 770
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1710841341
transform 1 0 1384 0 1 770
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1710841341
transform 1 0 1376 0 1 770
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1710841341
transform 1 0 1368 0 1 770
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1710841341
transform 1 0 1336 0 1 770
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1710841341
transform 1 0 1328 0 1 770
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1710841341
transform 1 0 1320 0 1 770
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1710841341
transform 1 0 1288 0 1 770
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1710841341
transform 1 0 1280 0 1 770
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1710841341
transform 1 0 1272 0 1 770
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1710841341
transform 1 0 1264 0 1 770
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1710841341
transform 1 0 1232 0 1 770
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1710841341
transform 1 0 1208 0 1 770
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1710841341
transform 1 0 1200 0 1 770
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1710841341
transform 1 0 1192 0 1 770
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1710841341
transform 1 0 1184 0 1 770
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1710841341
transform 1 0 1144 0 1 770
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1710841341
transform 1 0 1136 0 1 770
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1710841341
transform 1 0 1112 0 1 770
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1710841341
transform 1 0 1104 0 1 770
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1710841341
transform 1 0 1096 0 1 770
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1710841341
transform 1 0 1056 0 1 770
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1710841341
transform 1 0 1048 0 1 770
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1710841341
transform 1 0 1040 0 1 770
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1710841341
transform 1 0 1000 0 1 770
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1710841341
transform 1 0 992 0 1 770
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1710841341
transform 1 0 984 0 1 770
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1710841341
transform 1 0 944 0 1 770
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1710841341
transform 1 0 936 0 1 770
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1710841341
transform 1 0 912 0 1 770
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1710841341
transform 1 0 904 0 1 770
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1710841341
transform 1 0 896 0 1 770
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1710841341
transform 1 0 888 0 1 770
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1710841341
transform 1 0 840 0 1 770
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1710841341
transform 1 0 832 0 1 770
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1710841341
transform 1 0 824 0 1 770
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1710841341
transform 1 0 792 0 1 770
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1710841341
transform 1 0 768 0 1 770
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1710841341
transform 1 0 760 0 1 770
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1710841341
transform 1 0 752 0 1 770
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1710841341
transform 1 0 720 0 1 770
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1710841341
transform 1 0 712 0 1 770
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1710841341
transform 1 0 680 0 1 770
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1710841341
transform 1 0 672 0 1 770
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1710841341
transform 1 0 664 0 1 770
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1710841341
transform 1 0 616 0 1 770
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1710841341
transform 1 0 576 0 1 770
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1710841341
transform 1 0 568 0 1 770
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1710841341
transform 1 0 504 0 1 770
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1710841341
transform 1 0 496 0 1 770
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1710841341
transform 1 0 488 0 1 770
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1710841341
transform 1 0 480 0 1 770
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1710841341
transform 1 0 448 0 1 770
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1710841341
transform 1 0 400 0 1 770
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1710841341
transform 1 0 392 0 1 770
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1710841341
transform 1 0 384 0 1 770
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1710841341
transform 1 0 336 0 1 770
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1710841341
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1710841341
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1710841341
transform 1 0 240 0 1 770
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1710841341
transform 1 0 232 0 1 770
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1710841341
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1710841341
transform 1 0 160 0 1 770
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1710841341
transform 1 0 152 0 1 770
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1710841341
transform 1 0 144 0 1 770
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1710841341
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1710841341
transform 1 0 2664 0 -1 770
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1710841341
transform 1 0 2632 0 -1 770
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1710841341
transform 1 0 2624 0 -1 770
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1710841341
transform 1 0 2616 0 -1 770
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1710841341
transform 1 0 2576 0 -1 770
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1710841341
transform 1 0 2568 0 -1 770
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1710841341
transform 1 0 2560 0 -1 770
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1710841341
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1710841341
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1710841341
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1710841341
transform 1 0 2464 0 -1 770
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1710841341
transform 1 0 2456 0 -1 770
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1710841341
transform 1 0 2448 0 -1 770
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1710841341
transform 1 0 2416 0 -1 770
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1710841341
transform 1 0 2408 0 -1 770
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1710841341
transform 1 0 2360 0 -1 770
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1710841341
transform 1 0 2352 0 -1 770
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1710841341
transform 1 0 2344 0 -1 770
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1710841341
transform 1 0 2288 0 -1 770
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1710841341
transform 1 0 2280 0 -1 770
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1710841341
transform 1 0 2272 0 -1 770
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1710841341
transform 1 0 2232 0 -1 770
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1710841341
transform 1 0 2224 0 -1 770
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1710841341
transform 1 0 2184 0 -1 770
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1710841341
transform 1 0 2176 0 -1 770
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1710841341
transform 1 0 2168 0 -1 770
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1710841341
transform 1 0 2120 0 -1 770
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1710841341
transform 1 0 2112 0 -1 770
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1710841341
transform 1 0 2104 0 -1 770
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1710841341
transform 1 0 2056 0 -1 770
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1710841341
transform 1 0 2032 0 -1 770
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1710841341
transform 1 0 2024 0 -1 770
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1710841341
transform 1 0 2016 0 -1 770
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1710841341
transform 1 0 1984 0 -1 770
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1710841341
transform 1 0 1976 0 -1 770
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1710841341
transform 1 0 1936 0 -1 770
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1710841341
transform 1 0 1832 0 -1 770
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1710841341
transform 1 0 1824 0 -1 770
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1710841341
transform 1 0 1776 0 -1 770
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1710841341
transform 1 0 1768 0 -1 770
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1710841341
transform 1 0 1760 0 -1 770
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1710841341
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1710841341
transform 1 0 1720 0 -1 770
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1710841341
transform 1 0 1688 0 -1 770
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1710841341
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1710841341
transform 1 0 1672 0 -1 770
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1710841341
transform 1 0 1664 0 -1 770
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1710841341
transform 1 0 1624 0 -1 770
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1710841341
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1710841341
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1710841341
transform 1 0 1560 0 -1 770
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1710841341
transform 1 0 1552 0 -1 770
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1710841341
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1710841341
transform 1 0 1536 0 -1 770
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1710841341
transform 1 0 1480 0 -1 770
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1710841341
transform 1 0 1472 0 -1 770
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1710841341
transform 1 0 1464 0 -1 770
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1710841341
transform 1 0 1432 0 -1 770
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1710841341
transform 1 0 1424 0 -1 770
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1710841341
transform 1 0 1416 0 -1 770
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1710841341
transform 1 0 1376 0 -1 770
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1710841341
transform 1 0 1368 0 -1 770
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1710841341
transform 1 0 1336 0 -1 770
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1710841341
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1710841341
transform 1 0 1304 0 -1 770
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1710841341
transform 1 0 1296 0 -1 770
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1710841341
transform 1 0 1264 0 -1 770
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1710841341
transform 1 0 1256 0 -1 770
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1710841341
transform 1 0 1248 0 -1 770
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1710841341
transform 1 0 1240 0 -1 770
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1710841341
transform 1 0 1192 0 -1 770
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1710841341
transform 1 0 1184 0 -1 770
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1710841341
transform 1 0 1176 0 -1 770
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1710841341
transform 1 0 1168 0 -1 770
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1710841341
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1710841341
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1710841341
transform 1 0 1096 0 -1 770
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1710841341
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1710841341
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1710841341
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1710841341
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1710841341
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1710841341
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1710841341
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1710841341
transform 1 0 976 0 -1 770
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1710841341
transform 1 0 968 0 -1 770
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1710841341
transform 1 0 936 0 -1 770
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1710841341
transform 1 0 928 0 -1 770
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1710841341
transform 1 0 920 0 -1 770
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1710841341
transform 1 0 888 0 -1 770
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1710841341
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1710841341
transform 1 0 856 0 -1 770
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1710841341
transform 1 0 848 0 -1 770
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1710841341
transform 1 0 840 0 -1 770
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1710841341
transform 1 0 800 0 -1 770
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1710841341
transform 1 0 792 0 -1 770
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1710841341
transform 1 0 784 0 -1 770
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1710841341
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1710841341
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1710841341
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1710841341
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1710841341
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1710841341
transform 1 0 664 0 -1 770
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1710841341
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1710841341
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1710841341
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1710841341
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1710841341
transform 1 0 592 0 -1 770
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1710841341
transform 1 0 584 0 -1 770
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1710841341
transform 1 0 552 0 -1 770
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1710841341
transform 1 0 544 0 -1 770
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1710841341
transform 1 0 536 0 -1 770
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1710841341
transform 1 0 528 0 -1 770
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1710841341
transform 1 0 488 0 -1 770
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1710841341
transform 1 0 480 0 -1 770
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1710841341
transform 1 0 472 0 -1 770
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1710841341
transform 1 0 432 0 -1 770
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1710841341
transform 1 0 424 0 -1 770
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1710841341
transform 1 0 320 0 -1 770
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1710841341
transform 1 0 312 0 -1 770
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1710841341
transform 1 0 304 0 -1 770
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1710841341
transform 1 0 296 0 -1 770
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1710841341
transform 1 0 256 0 -1 770
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1710841341
transform 1 0 248 0 -1 770
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1710841341
transform 1 0 240 0 -1 770
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1710841341
transform 1 0 232 0 -1 770
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1710841341
transform 1 0 192 0 -1 770
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1710841341
transform 1 0 152 0 -1 770
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1710841341
transform 1 0 144 0 -1 770
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1710841341
transform 1 0 136 0 -1 770
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1710841341
transform 1 0 128 0 -1 770
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1710841341
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1710841341
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1710841341
transform 1 0 2568 0 1 570
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1710841341
transform 1 0 2560 0 1 570
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1710841341
transform 1 0 2520 0 1 570
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1710841341
transform 1 0 2512 0 1 570
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1710841341
transform 1 0 2504 0 1 570
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1710841341
transform 1 0 2400 0 1 570
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1710841341
transform 1 0 2392 0 1 570
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1710841341
transform 1 0 2384 0 1 570
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1710841341
transform 1 0 2344 0 1 570
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1710841341
transform 1 0 2336 0 1 570
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1710841341
transform 1 0 2312 0 1 570
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1710841341
transform 1 0 2304 0 1 570
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1710841341
transform 1 0 2296 0 1 570
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1710841341
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1710841341
transform 1 0 2256 0 1 570
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1710841341
transform 1 0 2216 0 1 570
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1710841341
transform 1 0 2208 0 1 570
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1710841341
transform 1 0 2184 0 1 570
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1710841341
transform 1 0 2176 0 1 570
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1710841341
transform 1 0 2136 0 1 570
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1710841341
transform 1 0 2128 0 1 570
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1710841341
transform 1 0 2120 0 1 570
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1710841341
transform 1 0 2112 0 1 570
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1710841341
transform 1 0 2104 0 1 570
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1710841341
transform 1 0 2056 0 1 570
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1710841341
transform 1 0 2048 0 1 570
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1710841341
transform 1 0 2040 0 1 570
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1710841341
transform 1 0 2032 0 1 570
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1710841341
transform 1 0 2008 0 1 570
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1710841341
transform 1 0 1976 0 1 570
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1710841341
transform 1 0 1968 0 1 570
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1710841341
transform 1 0 1960 0 1 570
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1710841341
transform 1 0 1936 0 1 570
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1710841341
transform 1 0 1928 0 1 570
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1710841341
transform 1 0 1888 0 1 570
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1710841341
transform 1 0 1880 0 1 570
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1710841341
transform 1 0 1872 0 1 570
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1710841341
transform 1 0 1864 0 1 570
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1710841341
transform 1 0 1824 0 1 570
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1710841341
transform 1 0 1816 0 1 570
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1710841341
transform 1 0 1808 0 1 570
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1710841341
transform 1 0 1768 0 1 570
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1710841341
transform 1 0 1760 0 1 570
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1710841341
transform 1 0 1720 0 1 570
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1710841341
transform 1 0 1712 0 1 570
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1710841341
transform 1 0 1704 0 1 570
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1710841341
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1710841341
transform 1 0 1656 0 1 570
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1710841341
transform 1 0 1648 0 1 570
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1710841341
transform 1 0 1624 0 1 570
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1710841341
transform 1 0 1616 0 1 570
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1710841341
transform 1 0 1608 0 1 570
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1710841341
transform 1 0 1560 0 1 570
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1710841341
transform 1 0 1552 0 1 570
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1710841341
transform 1 0 1544 0 1 570
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1710841341
transform 1 0 1512 0 1 570
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1710841341
transform 1 0 1504 0 1 570
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1710841341
transform 1 0 1496 0 1 570
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1710841341
transform 1 0 1456 0 1 570
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1710841341
transform 1 0 1448 0 1 570
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1710841341
transform 1 0 1408 0 1 570
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1710841341
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1710841341
transform 1 0 1392 0 1 570
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1710841341
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1710841341
transform 1 0 1344 0 1 570
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1710841341
transform 1 0 1336 0 1 570
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1710841341
transform 1 0 1328 0 1 570
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1710841341
transform 1 0 1288 0 1 570
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1710841341
transform 1 0 1280 0 1 570
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1710841341
transform 1 0 1240 0 1 570
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1710841341
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1710841341
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1710841341
transform 1 0 1200 0 1 570
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1710841341
transform 1 0 1192 0 1 570
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1710841341
transform 1 0 1160 0 1 570
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1710841341
transform 1 0 1152 0 1 570
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1710841341
transform 1 0 1144 0 1 570
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1710841341
transform 1 0 1088 0 1 570
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1710841341
transform 1 0 1080 0 1 570
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1710841341
transform 1 0 1072 0 1 570
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1710841341
transform 1 0 968 0 1 570
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1710841341
transform 1 0 960 0 1 570
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1710841341
transform 1 0 912 0 1 570
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1710841341
transform 1 0 904 0 1 570
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1710841341
transform 1 0 896 0 1 570
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1710841341
transform 1 0 888 0 1 570
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1710841341
transform 1 0 840 0 1 570
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1710841341
transform 1 0 832 0 1 570
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1710841341
transform 1 0 824 0 1 570
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1710841341
transform 1 0 800 0 1 570
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1710841341
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1710841341
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1710841341
transform 1 0 744 0 1 570
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1710841341
transform 1 0 640 0 1 570
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1710841341
transform 1 0 632 0 1 570
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1710841341
transform 1 0 608 0 1 570
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1710841341
transform 1 0 568 0 1 570
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1710841341
transform 1 0 560 0 1 570
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1710841341
transform 1 0 552 0 1 570
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1710841341
transform 1 0 496 0 1 570
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1710841341
transform 1 0 488 0 1 570
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1710841341
transform 1 0 480 0 1 570
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1710841341
transform 1 0 472 0 1 570
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1710841341
transform 1 0 432 0 1 570
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1710841341
transform 1 0 424 0 1 570
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1710841341
transform 1 0 400 0 1 570
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1710841341
transform 1 0 392 0 1 570
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1710841341
transform 1 0 384 0 1 570
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1710841341
transform 1 0 360 0 1 570
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1710841341
transform 1 0 352 0 1 570
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1710841341
transform 1 0 320 0 1 570
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1710841341
transform 1 0 312 0 1 570
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1710841341
transform 1 0 304 0 1 570
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1710841341
transform 1 0 280 0 1 570
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1710841341
transform 1 0 272 0 1 570
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1710841341
transform 1 0 232 0 1 570
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1710841341
transform 1 0 224 0 1 570
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1710841341
transform 1 0 216 0 1 570
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1710841341
transform 1 0 208 0 1 570
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1710841341
transform 1 0 200 0 1 570
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1710841341
transform 1 0 152 0 1 570
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1710841341
transform 1 0 144 0 1 570
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1710841341
transform 1 0 136 0 1 570
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1710841341
transform 1 0 128 0 1 570
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1710841341
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1710841341
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1710841341
transform 1 0 2664 0 -1 570
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1710841341
transform 1 0 2656 0 -1 570
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1710841341
transform 1 0 2616 0 -1 570
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1710841341
transform 1 0 2608 0 -1 570
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1710841341
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1710841341
transform 1 0 2592 0 -1 570
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1710841341
transform 1 0 2584 0 -1 570
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1710841341
transform 1 0 2576 0 -1 570
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1710841341
transform 1 0 2544 0 -1 570
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1710841341
transform 1 0 2512 0 -1 570
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1710841341
transform 1 0 2504 0 -1 570
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1710841341
transform 1 0 2496 0 -1 570
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1710841341
transform 1 0 2488 0 -1 570
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1710841341
transform 1 0 2480 0 -1 570
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1710841341
transform 1 0 2472 0 -1 570
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1710841341
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1710841341
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1710841341
transform 1 0 2416 0 -1 570
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1710841341
transform 1 0 2408 0 -1 570
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1710841341
transform 1 0 2368 0 -1 570
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1710841341
transform 1 0 2360 0 -1 570
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1710841341
transform 1 0 2352 0 -1 570
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1710841341
transform 1 0 2344 0 -1 570
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1710841341
transform 1 0 2296 0 -1 570
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1710841341
transform 1 0 2288 0 -1 570
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1710841341
transform 1 0 2280 0 -1 570
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1710841341
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1710841341
transform 1 0 2232 0 -1 570
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1710841341
transform 1 0 2224 0 -1 570
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1710841341
transform 1 0 2184 0 -1 570
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1710841341
transform 1 0 2176 0 -1 570
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1710841341
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1710841341
transform 1 0 2128 0 -1 570
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1710841341
transform 1 0 2120 0 -1 570
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1710841341
transform 1 0 2112 0 -1 570
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1710841341
transform 1 0 2064 0 -1 570
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1710841341
transform 1 0 2056 0 -1 570
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1710841341
transform 1 0 2048 0 -1 570
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1710841341
transform 1 0 2008 0 -1 570
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1710841341
transform 1 0 2000 0 -1 570
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1710841341
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1710841341
transform 1 0 1952 0 -1 570
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1710841341
transform 1 0 1944 0 -1 570
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1710841341
transform 1 0 1936 0 -1 570
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1710841341
transform 1 0 1888 0 -1 570
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1710841341
transform 1 0 1880 0 -1 570
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1710841341
transform 1 0 1872 0 -1 570
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1710841341
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1710841341
transform 1 0 1792 0 -1 570
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1710841341
transform 1 0 1784 0 -1 570
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1710841341
transform 1 0 1776 0 -1 570
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1710841341
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1710841341
transform 1 0 1728 0 -1 570
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1710841341
transform 1 0 1688 0 -1 570
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1710841341
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1710841341
transform 1 0 1672 0 -1 570
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1710841341
transform 1 0 1648 0 -1 570
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1710841341
transform 1 0 1608 0 -1 570
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1710841341
transform 1 0 1600 0 -1 570
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1710841341
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1710841341
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1710841341
transform 1 0 1528 0 -1 570
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1710841341
transform 1 0 1520 0 -1 570
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1710841341
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1710841341
transform 1 0 1504 0 -1 570
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1710841341
transform 1 0 1456 0 -1 570
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1710841341
transform 1 0 1448 0 -1 570
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1710841341
transform 1 0 1440 0 -1 570
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1710841341
transform 1 0 1408 0 -1 570
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1710841341
transform 1 0 1400 0 -1 570
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1710841341
transform 1 0 1352 0 -1 570
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1710841341
transform 1 0 1344 0 -1 570
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1710841341
transform 1 0 1336 0 -1 570
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1710841341
transform 1 0 1312 0 -1 570
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1710841341
transform 1 0 1288 0 -1 570
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1710841341
transform 1 0 1256 0 -1 570
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1710841341
transform 1 0 1248 0 -1 570
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1710841341
transform 1 0 1240 0 -1 570
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1710841341
transform 1 0 1192 0 -1 570
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1710841341
transform 1 0 1160 0 -1 570
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1710841341
transform 1 0 1152 0 -1 570
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1710841341
transform 1 0 1144 0 -1 570
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1710841341
transform 1 0 1104 0 -1 570
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1710841341
transform 1 0 1096 0 -1 570
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1710841341
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1710841341
transform 1 0 1048 0 -1 570
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1710841341
transform 1 0 1024 0 -1 570
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1710841341
transform 1 0 1016 0 -1 570
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1710841341
transform 1 0 1008 0 -1 570
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1710841341
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1710841341
transform 1 0 952 0 -1 570
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1710841341
transform 1 0 928 0 -1 570
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1710841341
transform 1 0 920 0 -1 570
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1710841341
transform 1 0 896 0 -1 570
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1710841341
transform 1 0 888 0 -1 570
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1710841341
transform 1 0 840 0 -1 570
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1710841341
transform 1 0 832 0 -1 570
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1710841341
transform 1 0 784 0 -1 570
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1710841341
transform 1 0 776 0 -1 570
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1710841341
transform 1 0 768 0 -1 570
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1710841341
transform 1 0 720 0 -1 570
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1710841341
transform 1 0 712 0 -1 570
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1710841341
transform 1 0 704 0 -1 570
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1710841341
transform 1 0 664 0 -1 570
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1710841341
transform 1 0 656 0 -1 570
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1710841341
transform 1 0 648 0 -1 570
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1710841341
transform 1 0 640 0 -1 570
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1710841341
transform 1 0 584 0 -1 570
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1710841341
transform 1 0 576 0 -1 570
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1710841341
transform 1 0 568 0 -1 570
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1710841341
transform 1 0 560 0 -1 570
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1710841341
transform 1 0 512 0 -1 570
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1710841341
transform 1 0 472 0 -1 570
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1710841341
transform 1 0 464 0 -1 570
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1710841341
transform 1 0 432 0 -1 570
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1710841341
transform 1 0 424 0 -1 570
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1710841341
transform 1 0 384 0 -1 570
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1710841341
transform 1 0 376 0 -1 570
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1710841341
transform 1 0 368 0 -1 570
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1710841341
transform 1 0 328 0 -1 570
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1710841341
transform 1 0 320 0 -1 570
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1710841341
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1710841341
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1710841341
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1710841341
transform 1 0 240 0 -1 570
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1710841341
transform 1 0 232 0 -1 570
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1710841341
transform 1 0 192 0 -1 570
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1710841341
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1710841341
transform 1 0 176 0 -1 570
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1710841341
transform 1 0 168 0 -1 570
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1710841341
transform 1 0 136 0 -1 570
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1710841341
transform 1 0 128 0 -1 570
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1710841341
transform 1 0 120 0 -1 570
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1710841341
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1710841341
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1710841341
transform 1 0 2664 0 1 370
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1710841341
transform 1 0 2656 0 1 370
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1710841341
transform 1 0 2616 0 1 370
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1710841341
transform 1 0 2608 0 1 370
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1710841341
transform 1 0 2600 0 1 370
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1710841341
transform 1 0 2592 0 1 370
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1710841341
transform 1 0 2552 0 1 370
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1710841341
transform 1 0 2544 0 1 370
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1710841341
transform 1 0 2536 0 1 370
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1710841341
transform 1 0 2504 0 1 370
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1710841341
transform 1 0 2496 0 1 370
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1710841341
transform 1 0 2488 0 1 370
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1710841341
transform 1 0 2480 0 1 370
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1710841341
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1710841341
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1710841341
transform 1 0 2424 0 1 370
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1710841341
transform 1 0 2416 0 1 370
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1710841341
transform 1 0 2368 0 1 370
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1710841341
transform 1 0 2360 0 1 370
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1710841341
transform 1 0 2352 0 1 370
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1710841341
transform 1 0 2304 0 1 370
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1710841341
transform 1 0 2280 0 1 370
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1710841341
transform 1 0 2272 0 1 370
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1710841341
transform 1 0 2264 0 1 370
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1710841341
transform 1 0 2216 0 1 370
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1710841341
transform 1 0 2208 0 1 370
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1710841341
transform 1 0 2200 0 1 370
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1710841341
transform 1 0 2192 0 1 370
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1710841341
transform 1 0 2144 0 1 370
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1710841341
transform 1 0 2120 0 1 370
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1710841341
transform 1 0 2112 0 1 370
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1710841341
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1710841341
transform 1 0 2064 0 1 370
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1710841341
transform 1 0 2056 0 1 370
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1710841341
transform 1 0 2016 0 1 370
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1710841341
transform 1 0 2008 0 1 370
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1710841341
transform 1 0 1984 0 1 370
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1710841341
transform 1 0 1976 0 1 370
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1710841341
transform 1 0 1944 0 1 370
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1710841341
transform 1 0 1936 0 1 370
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1710841341
transform 1 0 1888 0 1 370
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1710841341
transform 1 0 1880 0 1 370
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1710841341
transform 1 0 1872 0 1 370
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1710841341
transform 1 0 1848 0 1 370
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1710841341
transform 1 0 1840 0 1 370
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1710841341
transform 1 0 1792 0 1 370
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1710841341
transform 1 0 1784 0 1 370
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1710841341
transform 1 0 1776 0 1 370
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1710841341
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1710841341
transform 1 0 1696 0 1 370
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1710841341
transform 1 0 1688 0 1 370
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1710841341
transform 1 0 1648 0 1 370
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1710841341
transform 1 0 1600 0 1 370
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1710841341
transform 1 0 1592 0 1 370
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1710841341
transform 1 0 1584 0 1 370
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1710841341
transform 1 0 1544 0 1 370
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1710841341
transform 1 0 1504 0 1 370
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1710841341
transform 1 0 1496 0 1 370
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1710841341
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1710841341
transform 1 0 1448 0 1 370
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1710841341
transform 1 0 1440 0 1 370
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1710841341
transform 1 0 1400 0 1 370
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1710841341
transform 1 0 1368 0 1 370
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1710841341
transform 1 0 1360 0 1 370
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1710841341
transform 1 0 1336 0 1 370
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1710841341
transform 1 0 1328 0 1 370
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1710841341
transform 1 0 1320 0 1 370
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1710841341
transform 1 0 1280 0 1 370
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1710841341
transform 1 0 1272 0 1 370
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1710841341
transform 1 0 1232 0 1 370
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1710841341
transform 1 0 1224 0 1 370
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1710841341
transform 1 0 1216 0 1 370
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1710841341
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1710841341
transform 1 0 1160 0 1 370
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1710841341
transform 1 0 1136 0 1 370
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1710841341
transform 1 0 1128 0 1 370
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1710841341
transform 1 0 1120 0 1 370
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1710841341
transform 1 0 1072 0 1 370
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1710841341
transform 1 0 1064 0 1 370
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1710841341
transform 1 0 1040 0 1 370
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1710841341
transform 1 0 1032 0 1 370
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1710841341
transform 1 0 1000 0 1 370
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1710841341
transform 1 0 992 0 1 370
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1710841341
transform 1 0 960 0 1 370
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1710841341
transform 1 0 952 0 1 370
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1710841341
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1710841341
transform 1 0 904 0 1 370
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1710841341
transform 1 0 896 0 1 370
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1710841341
transform 1 0 888 0 1 370
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1710841341
transform 1 0 848 0 1 370
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1710841341
transform 1 0 840 0 1 370
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1710841341
transform 1 0 832 0 1 370
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1710841341
transform 1 0 824 0 1 370
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1710841341
transform 1 0 784 0 1 370
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1710841341
transform 1 0 776 0 1 370
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1710841341
transform 1 0 768 0 1 370
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1710841341
transform 1 0 728 0 1 370
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1710841341
transform 1 0 720 0 1 370
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1710841341
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1710841341
transform 1 0 688 0 1 370
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1710841341
transform 1 0 680 0 1 370
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1710841341
transform 1 0 640 0 1 370
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1710841341
transform 1 0 632 0 1 370
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1710841341
transform 1 0 608 0 1 370
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1710841341
transform 1 0 600 0 1 370
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1710841341
transform 1 0 592 0 1 370
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1710841341
transform 1 0 552 0 1 370
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1710841341
transform 1 0 512 0 1 370
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1710841341
transform 1 0 504 0 1 370
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1710841341
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1710841341
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1710841341
transform 1 0 448 0 1 370
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1710841341
transform 1 0 440 0 1 370
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1710841341
transform 1 0 392 0 1 370
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1710841341
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1710841341
transform 1 0 376 0 1 370
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1710841341
transform 1 0 352 0 1 370
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1710841341
transform 1 0 344 0 1 370
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1710841341
transform 1 0 304 0 1 370
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1710841341
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1710841341
transform 1 0 288 0 1 370
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1710841341
transform 1 0 280 0 1 370
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1710841341
transform 1 0 232 0 1 370
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1710841341
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1710841341
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1710841341
transform 1 0 176 0 1 370
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1710841341
transform 1 0 168 0 1 370
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1710841341
transform 1 0 160 0 1 370
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1710841341
transform 1 0 152 0 1 370
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1710841341
transform 1 0 144 0 1 370
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1710841341
transform 1 0 120 0 1 370
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1710841341
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1710841341
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1710841341
transform 1 0 2664 0 -1 370
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1710841341
transform 1 0 2656 0 -1 370
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1710841341
transform 1 0 2648 0 -1 370
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1710841341
transform 1 0 2592 0 -1 370
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1710841341
transform 1 0 2584 0 -1 370
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1710841341
transform 1 0 2576 0 -1 370
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1710841341
transform 1 0 2568 0 -1 370
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1710841341
transform 1 0 2520 0 -1 370
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1710841341
transform 1 0 2512 0 -1 370
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1710841341
transform 1 0 2504 0 -1 370
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1710841341
transform 1 0 2480 0 -1 370
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1710841341
transform 1 0 2472 0 -1 370
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1710841341
transform 1 0 2440 0 -1 370
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1710841341
transform 1 0 2432 0 -1 370
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1710841341
transform 1 0 2424 0 -1 370
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1710841341
transform 1 0 2416 0 -1 370
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1710841341
transform 1 0 2384 0 -1 370
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1710841341
transform 1 0 2376 0 -1 370
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1710841341
transform 1 0 2336 0 -1 370
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1710841341
transform 1 0 2328 0 -1 370
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1710841341
transform 1 0 2320 0 -1 370
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1710841341
transform 1 0 2312 0 -1 370
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1710841341
transform 1 0 2280 0 -1 370
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1710841341
transform 1 0 2272 0 -1 370
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1710841341
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1710841341
transform 1 0 2224 0 -1 370
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1710841341
transform 1 0 2192 0 -1 370
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1710841341
transform 1 0 2184 0 -1 370
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1710841341
transform 1 0 2176 0 -1 370
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1710841341
transform 1 0 2128 0 -1 370
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1710841341
transform 1 0 2120 0 -1 370
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1710841341
transform 1 0 2096 0 -1 370
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1710841341
transform 1 0 2088 0 -1 370
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1710841341
transform 1 0 2080 0 -1 370
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1710841341
transform 1 0 2016 0 -1 370
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1710841341
transform 1 0 2008 0 -1 370
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1710841341
transform 1 0 2000 0 -1 370
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1710841341
transform 1 0 1976 0 -1 370
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1710841341
transform 1 0 1928 0 -1 370
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1710841341
transform 1 0 1920 0 -1 370
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1710841341
transform 1 0 1912 0 -1 370
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1710841341
transform 1 0 1872 0 -1 370
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1710841341
transform 1 0 1864 0 -1 370
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1710841341
transform 1 0 1824 0 -1 370
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1710841341
transform 1 0 1800 0 -1 370
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1710841341
transform 1 0 1792 0 -1 370
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1710841341
transform 1 0 1784 0 -1 370
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1710841341
transform 1 0 1736 0 -1 370
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1710841341
transform 1 0 1728 0 -1 370
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1710841341
transform 1 0 1696 0 -1 370
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1710841341
transform 1 0 1688 0 -1 370
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1710841341
transform 1 0 1664 0 -1 370
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1710841341
transform 1 0 1624 0 -1 370
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1710841341
transform 1 0 1616 0 -1 370
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1710841341
transform 1 0 1608 0 -1 370
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1710841341
transform 1 0 1568 0 -1 370
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1710841341
transform 1 0 1528 0 -1 370
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1710841341
transform 1 0 1520 0 -1 370
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1710841341
transform 1 0 1512 0 -1 370
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1710841341
transform 1 0 1504 0 -1 370
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1710841341
transform 1 0 1496 0 -1 370
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1710841341
transform 1 0 1440 0 -1 370
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1710841341
transform 1 0 1432 0 -1 370
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1710841341
transform 1 0 1376 0 -1 370
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1710841341
transform 1 0 1368 0 -1 370
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1710841341
transform 1 0 1360 0 -1 370
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1710841341
transform 1 0 1328 0 -1 370
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1710841341
transform 1 0 1320 0 -1 370
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1710841341
transform 1 0 1280 0 -1 370
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1710841341
transform 1 0 1272 0 -1 370
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1710841341
transform 1 0 1264 0 -1 370
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1710841341
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1710841341
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1710841341
transform 1 0 1184 0 -1 370
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1710841341
transform 1 0 1176 0 -1 370
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1710841341
transform 1 0 1168 0 -1 370
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1710841341
transform 1 0 1160 0 -1 370
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1710841341
transform 1 0 1112 0 -1 370
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1710841341
transform 1 0 1104 0 -1 370
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1710841341
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1710841341
transform 1 0 1064 0 -1 370
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1710841341
transform 1 0 1056 0 -1 370
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1710841341
transform 1 0 1048 0 -1 370
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1710841341
transform 1 0 992 0 -1 370
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1710841341
transform 1 0 984 0 -1 370
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1710841341
transform 1 0 976 0 -1 370
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1710841341
transform 1 0 968 0 -1 370
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1710841341
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1710841341
transform 1 0 896 0 -1 370
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1710841341
transform 1 0 888 0 -1 370
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1710841341
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1710841341
transform 1 0 840 0 -1 370
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1710841341
transform 1 0 832 0 -1 370
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1710841341
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1710841341
transform 1 0 776 0 -1 370
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1710841341
transform 1 0 768 0 -1 370
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1710841341
transform 1 0 760 0 -1 370
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1710841341
transform 1 0 704 0 -1 370
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1710841341
transform 1 0 696 0 -1 370
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1710841341
transform 1 0 688 0 -1 370
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1710841341
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1710841341
transform 1 0 648 0 -1 370
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1710841341
transform 1 0 640 0 -1 370
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1710841341
transform 1 0 592 0 -1 370
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1710841341
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1710841341
transform 1 0 576 0 -1 370
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1710841341
transform 1 0 568 0 -1 370
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1710841341
transform 1 0 536 0 -1 370
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1710841341
transform 1 0 528 0 -1 370
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1710841341
transform 1 0 504 0 -1 370
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1710841341
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1710841341
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1710841341
transform 1 0 456 0 -1 370
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1710841341
transform 1 0 448 0 -1 370
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1710841341
transform 1 0 400 0 -1 370
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1710841341
transform 1 0 392 0 -1 370
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1710841341
transform 1 0 384 0 -1 370
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1710841341
transform 1 0 376 0 -1 370
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1710841341
transform 1 0 328 0 -1 370
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1710841341
transform 1 0 320 0 -1 370
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1710841341
transform 1 0 312 0 -1 370
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1710841341
transform 1 0 304 0 -1 370
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1710841341
transform 1 0 256 0 -1 370
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1710841341
transform 1 0 248 0 -1 370
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1710841341
transform 1 0 240 0 -1 370
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1710841341
transform 1 0 232 0 -1 370
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1710841341
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1710841341
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1710841341
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1710841341
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1710841341
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1710841341
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1710841341
transform 1 0 2664 0 1 170
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1710841341
transform 1 0 2640 0 1 170
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1710841341
transform 1 0 2632 0 1 170
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1710841341
transform 1 0 2624 0 1 170
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1710841341
transform 1 0 2576 0 1 170
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1710841341
transform 1 0 2568 0 1 170
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1710841341
transform 1 0 2560 0 1 170
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1710841341
transform 1 0 2552 0 1 170
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1710841341
transform 1 0 2520 0 1 170
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1710841341
transform 1 0 2512 0 1 170
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1710841341
transform 1 0 2504 0 1 170
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1710841341
transform 1 0 2464 0 1 170
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1710841341
transform 1 0 2456 0 1 170
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1710841341
transform 1 0 2448 0 1 170
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1710841341
transform 1 0 2440 0 1 170
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1710841341
transform 1 0 2408 0 1 170
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1710841341
transform 1 0 2400 0 1 170
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1710841341
transform 1 0 2392 0 1 170
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1710841341
transform 1 0 2344 0 1 170
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1710841341
transform 1 0 2336 0 1 170
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1710841341
transform 1 0 2328 0 1 170
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1710841341
transform 1 0 2320 0 1 170
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1710841341
transform 1 0 2312 0 1 170
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1710841341
transform 1 0 2272 0 1 170
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1710841341
transform 1 0 2264 0 1 170
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1710841341
transform 1 0 2256 0 1 170
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1710841341
transform 1 0 2216 0 1 170
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1710841341
transform 1 0 2208 0 1 170
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1710841341
transform 1 0 2200 0 1 170
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1710841341
transform 1 0 2168 0 1 170
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1710841341
transform 1 0 2160 0 1 170
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1710841341
transform 1 0 2152 0 1 170
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1710841341
transform 1 0 2144 0 1 170
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1710841341
transform 1 0 2136 0 1 170
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1710841341
transform 1 0 2104 0 1 170
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1710841341
transform 1 0 2096 0 1 170
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1710841341
transform 1 0 2064 0 1 170
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1710841341
transform 1 0 2056 0 1 170
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1710841341
transform 1 0 2048 0 1 170
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1710841341
transform 1 0 2040 0 1 170
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1710841341
transform 1 0 2032 0 1 170
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1710841341
transform 1 0 2024 0 1 170
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1710841341
transform 1 0 2016 0 1 170
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1710841341
transform 1 0 2008 0 1 170
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1710841341
transform 1 0 1968 0 1 170
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1710841341
transform 1 0 1960 0 1 170
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1710841341
transform 1 0 1952 0 1 170
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1710841341
transform 1 0 1944 0 1 170
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1710841341
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1710841341
transform 1 0 1896 0 1 170
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1710841341
transform 1 0 1888 0 1 170
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1710841341
transform 1 0 1856 0 1 170
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1710841341
transform 1 0 1848 0 1 170
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1710841341
transform 1 0 1840 0 1 170
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1710841341
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1710841341
transform 1 0 1784 0 1 170
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1710841341
transform 1 0 1776 0 1 170
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1710841341
transform 1 0 1768 0 1 170
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1710841341
transform 1 0 1760 0 1 170
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1710841341
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1710841341
transform 1 0 1712 0 1 170
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1710841341
transform 1 0 1704 0 1 170
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1710841341
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1710841341
transform 1 0 1648 0 1 170
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1710841341
transform 1 0 1640 0 1 170
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1710841341
transform 1 0 1632 0 1 170
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1710841341
transform 1 0 1624 0 1 170
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1710841341
transform 1 0 1616 0 1 170
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1710841341
transform 1 0 1560 0 1 170
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1710841341
transform 1 0 1552 0 1 170
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1710841341
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1710841341
transform 1 0 1512 0 1 170
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1710841341
transform 1 0 1504 0 1 170
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1710841341
transform 1 0 1456 0 1 170
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1710841341
transform 1 0 1448 0 1 170
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1710841341
transform 1 0 1440 0 1 170
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1710841341
transform 1 0 1416 0 1 170
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1710841341
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1710841341
transform 1 0 1376 0 1 170
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1710841341
transform 1 0 1344 0 1 170
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1710841341
transform 1 0 1336 0 1 170
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1710841341
transform 1 0 1328 0 1 170
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1710841341
transform 1 0 1288 0 1 170
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1710841341
transform 1 0 1280 0 1 170
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1710841341
transform 1 0 1272 0 1 170
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1710841341
transform 1 0 1232 0 1 170
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1710841341
transform 1 0 1224 0 1 170
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1710841341
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1710841341
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1710841341
transform 1 0 1184 0 1 170
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1710841341
transform 1 0 1136 0 1 170
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1710841341
transform 1 0 1128 0 1 170
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1710841341
transform 1 0 1120 0 1 170
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1710841341
transform 1 0 1112 0 1 170
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1710841341
transform 1 0 1072 0 1 170
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1710841341
transform 1 0 1064 0 1 170
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1710841341
transform 1 0 1056 0 1 170
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1710841341
transform 1 0 1048 0 1 170
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1710841341
transform 1 0 1040 0 1 170
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1710841341
transform 1 0 1000 0 1 170
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1710841341
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1710841341
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1710841341
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1710841341
transform 1 0 912 0 1 170
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1710841341
transform 1 0 904 0 1 170
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1710841341
transform 1 0 896 0 1 170
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1710841341
transform 1 0 888 0 1 170
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1710841341
transform 1 0 880 0 1 170
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1710841341
transform 1 0 840 0 1 170
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1710841341
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1710841341
transform 1 0 792 0 1 170
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1710841341
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1710841341
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1710841341
transform 1 0 768 0 1 170
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1710841341
transform 1 0 760 0 1 170
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1710841341
transform 1 0 720 0 1 170
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1710841341
transform 1 0 712 0 1 170
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1710841341
transform 1 0 680 0 1 170
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1710841341
transform 1 0 672 0 1 170
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1710841341
transform 1 0 664 0 1 170
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1710841341
transform 1 0 632 0 1 170
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1710841341
transform 1 0 624 0 1 170
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1710841341
transform 1 0 616 0 1 170
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1710841341
transform 1 0 576 0 1 170
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1710841341
transform 1 0 568 0 1 170
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1710841341
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1710841341
transform 1 0 520 0 1 170
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1710841341
transform 1 0 512 0 1 170
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1710841341
transform 1 0 504 0 1 170
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1710841341
transform 1 0 480 0 1 170
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1710841341
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1710841341
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1710841341
transform 1 0 424 0 1 170
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1710841341
transform 1 0 416 0 1 170
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1710841341
transform 1 0 408 0 1 170
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1710841341
transform 1 0 360 0 1 170
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1710841341
transform 1 0 352 0 1 170
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1710841341
transform 1 0 344 0 1 170
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1710841341
transform 1 0 336 0 1 170
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1710841341
transform 1 0 328 0 1 170
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1710841341
transform 1 0 320 0 1 170
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1710841341
transform 1 0 280 0 1 170
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1710841341
transform 1 0 272 0 1 170
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1710841341
transform 1 0 264 0 1 170
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1710841341
transform 1 0 256 0 1 170
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1710841341
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1710841341
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1710841341
transform 1 0 136 0 1 170
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1710841341
transform 1 0 128 0 1 170
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1710841341
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1710841341
transform 1 0 112 0 1 170
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1710841341
transform 1 0 104 0 1 170
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1710841341
transform 1 0 96 0 1 170
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1710841341
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1710841341
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1710841341
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1710841341
transform 1 0 2664 0 -1 170
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1710841341
transform 1 0 2656 0 -1 170
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1710841341
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1710841341
transform 1 0 2584 0 -1 170
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1710841341
transform 1 0 2576 0 -1 170
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1710841341
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1710841341
transform 1 0 2464 0 -1 170
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1710841341
transform 1 0 2456 0 -1 170
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1710841341
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1710841341
transform 1 0 2440 0 -1 170
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1710841341
transform 1 0 2400 0 -1 170
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1710841341
transform 1 0 2392 0 -1 170
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1710841341
transform 1 0 2384 0 -1 170
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1710841341
transform 1 0 2376 0 -1 170
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1710841341
transform 1 0 2368 0 -1 170
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1710841341
transform 1 0 2320 0 -1 170
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1710841341
transform 1 0 2312 0 -1 170
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1710841341
transform 1 0 2304 0 -1 170
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1710841341
transform 1 0 2296 0 -1 170
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1710841341
transform 1 0 2288 0 -1 170
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1710841341
transform 1 0 2256 0 -1 170
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1710841341
transform 1 0 2224 0 -1 170
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1710841341
transform 1 0 2216 0 -1 170
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1710841341
transform 1 0 2208 0 -1 170
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1710841341
transform 1 0 2200 0 -1 170
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1710841341
transform 1 0 2192 0 -1 170
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1710841341
transform 1 0 2152 0 -1 170
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1710841341
transform 1 0 2144 0 -1 170
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1710841341
transform 1 0 2136 0 -1 170
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1710841341
transform 1 0 2096 0 -1 170
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1710841341
transform 1 0 2088 0 -1 170
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1710841341
transform 1 0 1984 0 -1 170
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1710841341
transform 1 0 1976 0 -1 170
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1710841341
transform 1 0 1968 0 -1 170
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1710841341
transform 1 0 1944 0 -1 170
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1710841341
transform 1 0 1936 0 -1 170
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1710841341
transform 1 0 1928 0 -1 170
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1710841341
transform 1 0 1824 0 -1 170
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1710841341
transform 1 0 1816 0 -1 170
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1710841341
transform 1 0 1784 0 -1 170
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1710841341
transform 1 0 1776 0 -1 170
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1710841341
transform 1 0 1736 0 -1 170
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1710841341
transform 1 0 1728 0 -1 170
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1710841341
transform 1 0 1720 0 -1 170
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1710841341
transform 1 0 1616 0 -1 170
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1710841341
transform 1 0 1608 0 -1 170
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1710841341
transform 1 0 1600 0 -1 170
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1710841341
transform 1 0 1560 0 -1 170
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1710841341
transform 1 0 1552 0 -1 170
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1710841341
transform 1 0 1544 0 -1 170
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1710841341
transform 1 0 1536 0 -1 170
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1710841341
transform 1 0 1528 0 -1 170
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1710841341
transform 1 0 1480 0 -1 170
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1710841341
transform 1 0 1472 0 -1 170
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1710841341
transform 1 0 1464 0 -1 170
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1710841341
transform 1 0 1456 0 -1 170
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1710841341
transform 1 0 1408 0 -1 170
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1710841341
transform 1 0 1400 0 -1 170
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1710841341
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1710841341
transform 1 0 1360 0 -1 170
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1710841341
transform 1 0 1352 0 -1 170
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1710841341
transform 1 0 1344 0 -1 170
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1710841341
transform 1 0 1296 0 -1 170
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1710841341
transform 1 0 1288 0 -1 170
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1710841341
transform 1 0 1280 0 -1 170
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1710841341
transform 1 0 1248 0 -1 170
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1710841341
transform 1 0 1240 0 -1 170
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1710841341
transform 1 0 1208 0 -1 170
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1710841341
transform 1 0 1200 0 -1 170
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1710841341
transform 1 0 1160 0 -1 170
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1710841341
transform 1 0 1152 0 -1 170
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1710841341
transform 1 0 1048 0 -1 170
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1710841341
transform 1 0 1008 0 -1 170
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1710841341
transform 1 0 1000 0 -1 170
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1710841341
transform 1 0 968 0 -1 170
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1710841341
transform 1 0 960 0 -1 170
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1710841341
transform 1 0 928 0 -1 170
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1710841341
transform 1 0 920 0 -1 170
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1710841341
transform 1 0 872 0 -1 170
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1710841341
transform 1 0 864 0 -1 170
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1710841341
transform 1 0 832 0 -1 170
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1710841341
transform 1 0 824 0 -1 170
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1710841341
transform 1 0 720 0 -1 170
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1710841341
transform 1 0 712 0 -1 170
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1710841341
transform 1 0 704 0 -1 170
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1710841341
transform 1 0 672 0 -1 170
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1710841341
transform 1 0 664 0 -1 170
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1710841341
transform 1 0 624 0 -1 170
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1710841341
transform 1 0 616 0 -1 170
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1710841341
transform 1 0 608 0 -1 170
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1710841341
transform 1 0 600 0 -1 170
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1710841341
transform 1 0 568 0 -1 170
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1710841341
transform 1 0 536 0 -1 170
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1710841341
transform 1 0 528 0 -1 170
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1710841341
transform 1 0 520 0 -1 170
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1710841341
transform 1 0 512 0 -1 170
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1710841341
transform 1 0 464 0 -1 170
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1710841341
transform 1 0 456 0 -1 170
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1710841341
transform 1 0 432 0 -1 170
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1710841341
transform 1 0 424 0 -1 170
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1710841341
transform 1 0 416 0 -1 170
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1710841341
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1710841341
transform 1 0 344 0 -1 170
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1710841341
transform 1 0 336 0 -1 170
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1710841341
transform 1 0 232 0 -1 170
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1710841341
transform 1 0 224 0 -1 170
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1710841341
transform 1 0 216 0 -1 170
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1710841341
transform 1 0 208 0 -1 170
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1710841341
transform 1 0 200 0 -1 170
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1710841341
transform 1 0 192 0 -1 170
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1710841341
transform 1 0 184 0 -1 170
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1710841341
transform 1 0 176 0 -1 170
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1710841341
transform 1 0 168 0 -1 170
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1710841341
transform 1 0 160 0 -1 170
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1710841341
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1710841341
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1710841341
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1710841341
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1710841341
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1710841341
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1710841341
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1710841341
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1710841341
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1710841341
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1710841341
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1710841341
transform 1 0 72 0 -1 1770
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1710841341
transform 1 0 72 0 -1 1970
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1710841341
transform 1 0 72 0 1 1970
box -5 -3 84 105
use INVX1  INVX1_0
timestamp 1710841341
transform 1 0 2632 0 -1 170
box -9 -3 26 105
use INVX1  INVX1_1
timestamp 1710841341
transform 1 0 80 0 -1 1370
box -9 -3 26 105
use INVX1  INVX1_2
timestamp 1710841341
transform 1 0 352 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_0
timestamp 1710841341
transform 1 0 504 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1710841341
transform 1 0 744 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1710841341
transform 1 0 1392 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1710841341
transform 1 0 1608 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1710841341
transform 1 0 1048 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1710841341
transform 1 0 1344 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1710841341
transform 1 0 1064 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1710841341
transform 1 0 1848 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1710841341
transform 1 0 1376 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1710841341
transform 1 0 1360 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1710841341
transform 1 0 1344 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1710841341
transform 1 0 1504 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1710841341
transform 1 0 616 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1710841341
transform 1 0 1984 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1710841341
transform 1 0 2296 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1710841341
transform 1 0 1504 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1710841341
transform 1 0 504 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1710841341
transform 1 0 744 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1710841341
transform 1 0 2192 0 1 570
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1710841341
transform 1 0 2384 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1710841341
transform 1 0 408 0 1 570
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1710841341
transform 1 0 1488 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1710841341
transform 1 0 2408 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1710841341
transform 1 0 1512 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1710841341
transform 1 0 2288 0 1 970
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1710841341
transform 1 0 1488 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1710841341
transform 1 0 1776 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1710841341
transform 1 0 2272 0 1 970
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1710841341
transform 1 0 1544 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1710841341
transform 1 0 1408 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1710841341
transform 1 0 440 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1710841341
transform 1 0 432 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1710841341
transform 1 0 2520 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1710841341
transform 1 0 1800 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1710841341
transform 1 0 1592 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1710841341
transform 1 0 1128 0 1 570
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1710841341
transform 1 0 2016 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1710841341
transform 1 0 2080 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1710841341
transform 1 0 1072 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1710841341
transform 1 0 952 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1710841341
transform 1 0 1512 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1710841341
transform 1 0 368 0 1 770
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1710841341
transform 1 0 1312 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1710841341
transform 1 0 2128 0 1 370
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1710841341
transform 1 0 2096 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1710841341
transform 1 0 1992 0 1 370
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1710841341
transform 1 0 1560 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1710841341
transform 1 0 504 0 1 570
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1710841341
transform 1 0 2360 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1710841341
transform 1 0 2496 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1710841341
transform 1 0 1480 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1710841341
transform 1 0 656 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1710841341
transform 1 0 584 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1710841341
transform 1 0 1160 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1710841341
transform 1 0 544 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1710841341
transform 1 0 520 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1710841341
transform 1 0 600 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1710841341
transform 1 0 2016 0 1 570
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1710841341
transform 1 0 2264 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1710841341
transform 1 0 896 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1710841341
transform 1 0 1056 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1710841341
transform 1 0 1136 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1710841341
transform 1 0 936 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1710841341
transform 1 0 2040 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1710841341
transform 1 0 2144 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1710841341
transform 1 0 312 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1710841341
transform 1 0 968 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1710841341
transform 1 0 792 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1710841341
transform 1 0 808 0 1 570
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1710841341
transform 1 0 1992 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1710841341
transform 1 0 1728 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1710841341
transform 1 0 560 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1710841341
transform 1 0 792 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1710841341
transform 1 0 984 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1710841341
transform 1 0 904 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1710841341
transform 1 0 2032 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1710841341
transform 1 0 2136 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1710841341
transform 1 0 784 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1710841341
transform 1 0 720 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1710841341
transform 1 0 736 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1710841341
transform 1 0 616 0 1 570
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1710841341
transform 1 0 1632 0 1 570
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1710841341
transform 1 0 2528 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1710841341
transform 1 0 928 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1710841341
transform 1 0 1168 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1710841341
transform 1 0 1344 0 1 370
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1710841341
transform 1 0 1944 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1710841341
transform 1 0 1704 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1710841341
transform 1 0 232 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1710841341
transform 1 0 376 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1710841341
transform 1 0 288 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1710841341
transform 1 0 352 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1710841341
transform 1 0 112 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1710841341
transform 1 0 200 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1710841341
transform 1 0 440 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1710841341
transform 1 0 520 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1710841341
transform 1 0 416 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1710841341
transform 1 0 232 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1710841341
transform 1 0 288 0 1 570
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1710841341
transform 1 0 184 0 1 570
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1710841341
transform 1 0 416 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1710841341
transform 1 0 544 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1710841341
transform 1 0 392 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1710841341
transform 1 0 504 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1710841341
transform 1 0 552 0 1 970
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1710841341
transform 1 0 664 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1710841341
transform 1 0 776 0 1 770
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1710841341
transform 1 0 776 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1710841341
transform 1 0 760 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1710841341
transform 1 0 1216 0 1 770
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1710841341
transform 1 0 1120 0 1 770
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1710841341
transform 1 0 864 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1710841341
transform 1 0 1224 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1710841341
transform 1 0 992 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1710841341
transform 1 0 368 0 1 570
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1710841341
transform 1 0 360 0 1 370
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1710841341
transform 1 0 488 0 1 170
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1710841341
transform 1 0 704 0 1 370
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1710841341
transform 1 0 616 0 1 370
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1710841341
transform 1 0 440 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1710841341
transform 1 0 792 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1710841341
transform 1 0 1048 0 1 370
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1710841341
transform 1 0 1144 0 1 370
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1710841341
transform 1 0 1032 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1710841341
transform 1 0 984 0 1 170
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1710841341
transform 1 0 1120 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1710841341
transform 1 0 1296 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1710841341
transform 1 0 1320 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1710841341
transform 1 0 1208 0 1 570
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1710841341
transform 1 0 1208 0 1 170
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1710841341
transform 1 0 1480 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1710841341
transform 1 0 1384 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1710841341
transform 1 0 1728 0 1 170
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1710841341
transform 1 0 1744 0 1 170
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1710841341
transform 1 0 1600 0 1 170
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1710841341
transform 1 0 1672 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1710841341
transform 1 0 1656 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1710841341
transform 1 0 1808 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1710841341
transform 1 0 1856 0 1 370
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1710841341
transform 1 0 1944 0 1 570
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1710841341
transform 1 0 1784 0 1 770
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1710841341
transform 1 0 1680 0 1 770
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1710841341
transform 1 0 1488 0 1 770
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1710841341
transform 1 0 1840 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1710841341
transform 1 0 1528 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1710841341
transform 1 0 2352 0 1 770
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1710841341
transform 1 0 2328 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1710841341
transform 1 0 2320 0 1 770
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1710841341
transform 1 0 2152 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1710841341
transform 1 0 2280 0 1 170
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1710841341
transform 1 0 2248 0 1 370
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1710841341
transform 1 0 2288 0 1 370
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1710841341
transform 1 0 2296 0 1 170
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1710841341
transform 1 0 2488 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1710841341
transform 1 0 2152 0 1 370
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1710841341
transform 1 0 2024 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1710841341
transform 1 0 2104 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1710841341
transform 1 0 2648 0 1 170
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1710841341
transform 1 0 2600 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1710841341
transform 1 0 2464 0 1 970
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1710841341
transform 1 0 2368 0 1 970
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1710841341
transform 1 0 2648 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1710841341
transform 1 0 2456 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1710841341
transform 1 0 2200 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1710841341
transform 1 0 2296 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1710841341
transform 1 0 1992 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1710841341
transform 1 0 2248 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1710841341
transform 1 0 2432 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1710841341
transform 1 0 2120 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1710841341
transform 1 0 1800 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1710841341
transform 1 0 1744 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1710841341
transform 1 0 2080 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1710841341
transform 1 0 1848 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1710841341
transform 1 0 1720 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1710841341
transform 1 0 2432 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1710841341
transform 1 0 2512 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1710841341
transform 1 0 2592 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1710841341
transform 1 0 2416 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1710841341
transform 1 0 2408 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1710841341
transform 1 0 2360 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1710841341
transform 1 0 2512 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1710841341
transform 1 0 2320 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1710841341
transform 1 0 2224 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1710841341
transform 1 0 2192 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1710841341
transform 1 0 2288 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1710841341
transform 1 0 2288 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1710841341
transform 1 0 2016 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1710841341
transform 1 0 1856 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1710841341
transform 1 0 2008 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1710841341
transform 1 0 1976 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1710841341
transform 1 0 1920 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1710841341
transform 1 0 1608 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1710841341
transform 1 0 1520 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1710841341
transform 1 0 1688 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1710841341
transform 1 0 1736 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1710841341
transform 1 0 1640 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1710841341
transform 1 0 1704 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1710841341
transform 1 0 832 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1710841341
transform 1 0 752 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1710841341
transform 1 0 264 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1710841341
transform 1 0 1488 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1710841341
transform 1 0 1936 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1710841341
transform 1 0 2464 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1710841341
transform 1 0 2560 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1710841341
transform 1 0 2560 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1710841341
transform 1 0 576 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1710841341
transform 1 0 96 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1710841341
transform 1 0 80 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1710841341
transform 1 0 128 0 1 370
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1710841341
transform 1 0 744 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1710841341
transform 1 0 920 0 1 770
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1710841341
transform 1 0 2272 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1710841341
transform 1 0 1472 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1710841341
transform 1 0 512 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1710841341
transform 1 0 2376 0 1 370
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1710841341
transform 1 0 2528 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1710841341
transform 1 0 1344 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1710841341
transform 1 0 1424 0 1 170
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1710841341
transform 1 0 2520 0 1 970
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1710841341
transform 1 0 1384 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1710841341
transform 1 0 1208 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1710841341
transform 1 0 944 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1710841341
transform 1 0 784 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_223
timestamp 1710841341
transform 1 0 72 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1710841341
transform 1 0 304 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_225
timestamp 1710841341
transform 1 0 208 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_226
timestamp 1710841341
transform 1 0 112 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_227
timestamp 1710841341
transform 1 0 112 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_228
timestamp 1710841341
transform 1 0 320 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_229
timestamp 1710841341
transform 1 0 280 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_230
timestamp 1710841341
transform 1 0 272 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1710841341
transform 1 0 1640 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_232
timestamp 1710841341
transform 1 0 648 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1710841341
transform 1 0 1800 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_234
timestamp 1710841341
transform 1 0 1568 0 1 770
box -9 -3 26 105
use INVX2  INVX2_235
timestamp 1710841341
transform 1 0 536 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_236
timestamp 1710841341
transform 1 0 512 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_237
timestamp 1710841341
transform 1 0 808 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1710841341
transform 1 0 1640 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_239
timestamp 1710841341
transform 1 0 664 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1710841341
transform 1 0 656 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_241
timestamp 1710841341
transform 1 0 1032 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_242
timestamp 1710841341
transform 1 0 1624 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_243
timestamp 1710841341
transform 1 0 1320 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_244
timestamp 1710841341
transform 1 0 424 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_245
timestamp 1710841341
transform 1 0 1472 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1710841341
transform 1 0 1224 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_247
timestamp 1710841341
transform 1 0 1856 0 1 970
box -9 -3 26 105
use INVX2  INVX2_248
timestamp 1710841341
transform 1 0 2320 0 1 570
box -9 -3 26 105
use INVX2  INVX2_249
timestamp 1710841341
transform 1 0 1904 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_250
timestamp 1710841341
transform 1 0 2000 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_251
timestamp 1710841341
transform 1 0 240 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_252
timestamp 1710841341
transform 1 0 368 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_253
timestamp 1710841341
transform 1 0 200 0 1 970
box -9 -3 26 105
use INVX2  INVX2_254
timestamp 1710841341
transform 1 0 216 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_255
timestamp 1710841341
transform 1 0 1656 0 1 170
box -9 -3 26 105
use INVX2  INVX2_256
timestamp 1710841341
transform 1 0 1952 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_257
timestamp 1710841341
transform 1 0 2608 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_258
timestamp 1710841341
transform 1 0 2552 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_259
timestamp 1710841341
transform 1 0 2536 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_260
timestamp 1710841341
transform 1 0 2552 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_261
timestamp 1710841341
transform 1 0 1400 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_262
timestamp 1710841341
transform 1 0 1224 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_263
timestamp 1710841341
transform 1 0 1080 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_264
timestamp 1710841341
transform 1 0 928 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_265
timestamp 1710841341
transform 1 0 472 0 -1 1570
box -9 -3 26 105
use INVX8  INVX8_0
timestamp 1710841341
transform 1 0 2592 0 -1 170
box -9 -3 45 105
use M2_M1  M2_M1_0
timestamp 1710841341
transform 1 0 532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1710841341
transform 1 0 532 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1710841341
transform 1 0 500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1710841341
transform 1 0 492 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1710841341
transform 1 0 508 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1710841341
transform 1 0 508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1710841341
transform 1 0 468 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1710841341
transform 1 0 468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1710841341
transform 1 0 108 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1710841341
transform 1 0 84 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1710841341
transform 1 0 100 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1710841341
transform 1 0 84 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1710841341
transform 1 0 100 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1710841341
transform 1 0 76 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1710841341
transform 1 0 692 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1710841341
transform 1 0 660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1710841341
transform 1 0 660 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1710841341
transform 1 0 564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1710841341
transform 1 0 564 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1710841341
transform 1 0 540 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1710841341
transform 1 0 652 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1710841341
transform 1 0 596 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1710841341
transform 1 0 580 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1710841341
transform 1 0 556 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1710841341
transform 1 0 548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1710841341
transform 1 0 524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1710841341
transform 1 0 652 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1710841341
transform 1 0 644 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1710841341
transform 1 0 612 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1710841341
transform 1 0 588 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1710841341
transform 1 0 588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1710841341
transform 1 0 540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1710841341
transform 1 0 676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1710841341
transform 1 0 580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1710841341
transform 1 0 556 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1710841341
transform 1 0 492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1710841341
transform 1 0 644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1710841341
transform 1 0 604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1710841341
transform 1 0 508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1710841341
transform 1 0 388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1710841341
transform 1 0 2596 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1710841341
transform 1 0 2564 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1710841341
transform 1 0 2196 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1710841341
transform 1 0 2148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1710841341
transform 1 0 2100 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1710841341
transform 1 0 1980 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1710841341
transform 1 0 1236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1710841341
transform 1 0 836 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1710841341
transform 1 0 836 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1710841341
transform 1 0 748 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1710841341
transform 1 0 676 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1710841341
transform 1 0 676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1710841341
transform 1 0 652 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1710841341
transform 1 0 604 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1710841341
transform 1 0 524 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1710841341
transform 1 0 292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1710841341
transform 1 0 244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1710841341
transform 1 0 244 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1710841341
transform 1 0 204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1710841341
transform 1 0 204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1710841341
transform 1 0 740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1710841341
transform 1 0 676 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1710841341
transform 1 0 676 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1710841341
transform 1 0 668 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1710841341
transform 1 0 1476 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1710841341
transform 1 0 1468 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1710841341
transform 1 0 1420 0 1 1655
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1710841341
transform 1 0 1404 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1710841341
transform 1 0 1396 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1710841341
transform 1 0 1364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1710841341
transform 1 0 1364 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1710841341
transform 1 0 1340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1710841341
transform 1 0 428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1710841341
transform 1 0 420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1710841341
transform 1 0 1452 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1710841341
transform 1 0 1388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1710841341
transform 1 0 1388 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1710841341
transform 1 0 1380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1710841341
transform 1 0 1348 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1710841341
transform 1 0 492 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1710841341
transform 1 0 348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1710841341
transform 1 0 340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1710841341
transform 1 0 308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1710841341
transform 1 0 1052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1710841341
transform 1 0 956 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1710841341
transform 1 0 956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1710841341
transform 1 0 452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1710841341
transform 1 0 388 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1710841341
transform 1 0 316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1710841341
transform 1 0 1140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1710841341
transform 1 0 1092 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1710841341
transform 1 0 1004 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1710841341
transform 1 0 996 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1710841341
transform 1 0 348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1710841341
transform 1 0 220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1710841341
transform 1 0 836 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1710841341
transform 1 0 796 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1710841341
transform 1 0 764 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1710841341
transform 1 0 748 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1710841341
transform 1 0 716 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1710841341
transform 1 0 684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1710841341
transform 1 0 652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1710841341
transform 1 0 652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1710841341
transform 1 0 748 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1710841341
transform 1 0 700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1710841341
transform 1 0 524 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1710841341
transform 1 0 636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1710841341
transform 1 0 572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1710841341
transform 1 0 500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1710841341
transform 1 0 444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1710841341
transform 1 0 588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1710841341
transform 1 0 572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1710841341
transform 1 0 292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1710841341
transform 1 0 228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1710841341
transform 1 0 108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1710841341
transform 1 0 84 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1710841341
transform 1 0 84 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1710841341
transform 1 0 492 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1710841341
transform 1 0 492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1710841341
transform 1 0 428 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1710841341
transform 1 0 356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1710841341
transform 1 0 276 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1710841341
transform 1 0 220 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1710841341
transform 1 0 76 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1710841341
transform 1 0 76 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1710841341
transform 1 0 484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1710841341
transform 1 0 452 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1710841341
transform 1 0 292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1710841341
transform 1 0 76 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1710841341
transform 1 0 428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1710841341
transform 1 0 380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1710841341
transform 1 0 228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1710841341
transform 1 0 228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1710841341
transform 1 0 164 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1710841341
transform 1 0 76 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1710841341
transform 1 0 332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1710841341
transform 1 0 236 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1710841341
transform 1 0 204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1710841341
transform 1 0 132 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1710841341
transform 1 0 180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1710841341
transform 1 0 172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1710841341
transform 1 0 292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1710841341
transform 1 0 220 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1710841341
transform 1 0 180 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1710841341
transform 1 0 268 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1710841341
transform 1 0 228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1710841341
transform 1 0 188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1710841341
transform 1 0 268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1710841341
transform 1 0 204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1710841341
transform 1 0 812 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1710841341
transform 1 0 788 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1710841341
transform 1 0 764 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1710841341
transform 1 0 652 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1710841341
transform 1 0 524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1710841341
transform 1 0 804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1710841341
transform 1 0 780 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1710841341
transform 1 0 780 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1710841341
transform 1 0 780 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1710841341
transform 1 0 724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1710841341
transform 1 0 708 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1710841341
transform 1 0 1444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1710841341
transform 1 0 1404 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1710841341
transform 1 0 1348 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1710841341
transform 1 0 1324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1710841341
transform 1 0 1260 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1710841341
transform 1 0 1252 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1710841341
transform 1 0 2084 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1710841341
transform 1 0 2068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1710841341
transform 1 0 2060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1710841341
transform 1 0 2044 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1710841341
transform 1 0 2028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1710841341
transform 1 0 2012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1710841341
transform 1 0 1636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1710841341
transform 1 0 1548 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1710841341
transform 1 0 1516 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1710841341
transform 1 0 1004 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1710841341
transform 1 0 972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1710841341
transform 1 0 932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1710841341
transform 1 0 892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1710841341
transform 1 0 844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1710841341
transform 1 0 812 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1710841341
transform 1 0 796 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1710841341
transform 1 0 708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1710841341
transform 1 0 1620 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1710841341
transform 1 0 1580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1710841341
transform 1 0 1340 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1710841341
transform 1 0 1340 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1710841341
transform 1 0 1316 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1710841341
transform 1 0 1284 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1710841341
transform 1 0 1276 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1710841341
transform 1 0 1164 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1710841341
transform 1 0 1124 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1710841341
transform 1 0 1124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1710841341
transform 1 0 1108 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1710841341
transform 1 0 1108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1710841341
transform 1 0 1108 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1710841341
transform 1 0 1068 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1710841341
transform 1 0 1028 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1710841341
transform 1 0 1028 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1710841341
transform 1 0 1532 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1710841341
transform 1 0 1444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1710841341
transform 1 0 1060 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1710841341
transform 1 0 2060 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1710841341
transform 1 0 2044 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1710841341
transform 1 0 1820 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1710841341
transform 1 0 1644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1710841341
transform 1 0 1588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1710841341
transform 1 0 1452 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1710841341
transform 1 0 1324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1710841341
transform 1 0 1148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1710841341
transform 1 0 1124 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1710841341
transform 1 0 1124 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1710841341
transform 1 0 1100 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1710841341
transform 1 0 1100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1710841341
transform 1 0 1740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1710841341
transform 1 0 1700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1710841341
transform 1 0 1620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1710841341
transform 1 0 1524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1710841341
transform 1 0 1524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1710841341
transform 1 0 1452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1710841341
transform 1 0 1332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1710841341
transform 1 0 1332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1710841341
transform 1 0 1284 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1710841341
transform 1 0 1212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1710841341
transform 1 0 1212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1710841341
transform 1 0 1964 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1710841341
transform 1 0 1916 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1710841341
transform 1 0 1900 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1710841341
transform 1 0 1900 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1710841341
transform 1 0 1892 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1710841341
transform 1 0 1876 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1710841341
transform 1 0 1468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1710841341
transform 1 0 1396 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1710841341
transform 1 0 1396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1710841341
transform 1 0 1340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1710841341
transform 1 0 1412 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1710841341
transform 1 0 1380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1710841341
transform 1 0 1356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1710841341
transform 1 0 1356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1710841341
transform 1 0 1332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1710841341
transform 1 0 1332 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1710841341
transform 1 0 1332 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1710841341
transform 1 0 1420 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1710841341
transform 1 0 1420 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1710841341
transform 1 0 1380 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1710841341
transform 1 0 1364 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1710841341
transform 1 0 1348 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1710841341
transform 1 0 1652 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1710841341
transform 1 0 1612 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1710841341
transform 1 0 1516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1710841341
transform 1 0 1284 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1710841341
transform 1 0 1268 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1710841341
transform 1 0 860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1710841341
transform 1 0 796 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1710841341
transform 1 0 708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1710841341
transform 1 0 668 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1710841341
transform 1 0 2644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1710841341
transform 1 0 1996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1710841341
transform 1 0 1740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1710841341
transform 1 0 2324 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1710841341
transform 1 0 2316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1710841341
transform 1 0 2284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1710841341
transform 1 0 2260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1710841341
transform 1 0 1748 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1710841341
transform 1 0 1564 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1710841341
transform 1 0 1516 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1710841341
transform 1 0 1468 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1710841341
transform 1 0 1092 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1710841341
transform 1 0 684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1710841341
transform 1 0 492 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1710841341
transform 1 0 220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1710841341
transform 1 0 180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1710841341
transform 1 0 1876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1710841341
transform 1 0 828 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1710841341
transform 1 0 772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1710841341
transform 1 0 668 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1710841341
transform 1 0 636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1710841341
transform 1 0 2436 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1710841341
transform 1 0 2292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1710841341
transform 1 0 2284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1710841341
transform 1 0 2228 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1710841341
transform 1 0 2204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1710841341
transform 1 0 2180 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1710841341
transform 1 0 2548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1710841341
transform 1 0 2436 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1710841341
transform 1 0 2396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1710841341
transform 1 0 1604 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1710841341
transform 1 0 812 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1710841341
transform 1 0 388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1710841341
transform 1 0 380 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1710841341
transform 1 0 236 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1710841341
transform 1 0 180 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1710841341
transform 1 0 2228 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1710841341
transform 1 0 2220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1710841341
transform 1 0 1644 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1710841341
transform 1 0 1628 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1710841341
transform 1 0 1476 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1710841341
transform 1 0 1308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1710841341
transform 1 0 1260 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1710841341
transform 1 0 2532 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1710841341
transform 1 0 2484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1710841341
transform 1 0 2468 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1710841341
transform 1 0 2420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1710841341
transform 1 0 2380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1710841341
transform 1 0 2340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1710841341
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1710841341
transform 1 0 2052 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1710841341
transform 1 0 1876 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1710841341
transform 1 0 1820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1710841341
transform 1 0 1492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1710841341
transform 1 0 948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1710841341
transform 1 0 900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1710841341
transform 1 0 2436 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1710841341
transform 1 0 2340 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1710841341
transform 1 0 2308 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1710841341
transform 1 0 2164 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1710841341
transform 1 0 1764 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1710841341
transform 1 0 1700 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1710841341
transform 1 0 1644 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1710841341
transform 1 0 1604 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1710841341
transform 1 0 1492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1710841341
transform 1 0 1404 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1710841341
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1710841341
transform 1 0 1756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1710841341
transform 1 0 1756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1710841341
transform 1 0 1716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1710841341
transform 1 0 2340 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1710841341
transform 1 0 2316 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1710841341
transform 1 0 2308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1710841341
transform 1 0 2284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1710841341
transform 1 0 2284 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1710841341
transform 1 0 2252 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1710841341
transform 1 0 1604 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1710841341
transform 1 0 1580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1710841341
transform 1 0 1436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1710841341
transform 1 0 1420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1710841341
transform 1 0 1412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1710841341
transform 1 0 1292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1710841341
transform 1 0 1092 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1710841341
transform 1 0 444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1710841341
transform 1 0 436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1710841341
transform 1 0 292 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1710841341
transform 1 0 1508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1710841341
transform 1 0 476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1710841341
transform 1 0 476 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1710841341
transform 1 0 2596 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1710841341
transform 1 0 2556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1710841341
transform 1 0 2556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1710841341
transform 1 0 1836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1710841341
transform 1 0 1828 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1710841341
transform 1 0 1796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1710841341
transform 1 0 1476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1710841341
transform 1 0 1692 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1710841341
transform 1 0 1692 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1710841341
transform 1 0 1668 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1710841341
transform 1 0 1668 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1710841341
transform 1 0 1620 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1710841341
transform 1 0 1252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1710841341
transform 1 0 1236 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1710841341
transform 1 0 1276 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1710841341
transform 1 0 1148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1710841341
transform 1 0 1124 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1710841341
transform 1 0 2492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1710841341
transform 1 0 1996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1710841341
transform 1 0 1972 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1710841341
transform 1 0 1972 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1710841341
transform 1 0 2308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1710841341
transform 1 0 2084 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1710841341
transform 1 0 1980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1710841341
transform 1 0 1964 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1710841341
transform 1 0 1068 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1710841341
transform 1 0 1044 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1710841341
transform 1 0 948 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1710841341
transform 1 0 884 0 1 2007
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1710841341
transform 1 0 1748 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1710841341
transform 1 0 1508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1710841341
transform 1 0 1484 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1710841341
transform 1 0 1412 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1710841341
transform 1 0 1148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1710841341
transform 1 0 996 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1710841341
transform 1 0 380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1710841341
transform 1 0 228 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1710841341
transform 1 0 188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1710841341
transform 1 0 172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1710841341
transform 1 0 1404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1710841341
transform 1 0 1300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1710841341
transform 1 0 1108 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1710841341
transform 1 0 1020 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1710841341
transform 1 0 956 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1710841341
transform 1 0 2628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1710841341
transform 1 0 2556 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1710841341
transform 1 0 2476 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1710841341
transform 1 0 2140 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1710841341
transform 1 0 2108 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1710841341
transform 1 0 2100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1710841341
transform 1 0 2092 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1710841341
transform 1 0 2196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1710841341
transform 1 0 2156 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1710841341
transform 1 0 2116 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1710841341
transform 1 0 2116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1710841341
transform 1 0 2060 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1710841341
transform 1 0 1516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1710841341
transform 1 0 1460 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1710841341
transform 1 0 2268 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1710841341
transform 1 0 2260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1710841341
transform 1 0 2236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1710841341
transform 1 0 2004 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1710841341
transform 1 0 1492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1710841341
transform 1 0 1468 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1710841341
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1710841341
transform 1 0 1388 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1710841341
transform 1 0 1572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1710841341
transform 1 0 1556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1710841341
transform 1 0 1284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1710841341
transform 1 0 1268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1710841341
transform 1 0 580 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1710841341
transform 1 0 484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1710841341
transform 1 0 468 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1710841341
transform 1 0 436 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1710841341
transform 1 0 412 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1710841341
transform 1 0 2356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1710841341
transform 1 0 2324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1710841341
transform 1 0 2308 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1710841341
transform 1 0 2564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1710841341
transform 1 0 2508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1710841341
transform 1 0 1612 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1710841341
transform 1 0 1492 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1710841341
transform 1 0 1412 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1710841341
transform 1 0 700 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1710841341
transform 1 0 684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1710841341
transform 1 0 668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1710841341
transform 1 0 676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1710841341
transform 1 0 612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1710841341
transform 1 0 596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1710841341
transform 1 0 1260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1710841341
transform 1 0 1236 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1710841341
transform 1 0 1228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1710841341
transform 1 0 1196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1710841341
transform 1 0 700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1710841341
transform 1 0 660 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1710841341
transform 1 0 604 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1710841341
transform 1 0 556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1710841341
transform 1 0 540 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1710841341
transform 1 0 684 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1710841341
transform 1 0 660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1710841341
transform 1 0 652 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1710841341
transform 1 0 628 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1710841341
transform 1 0 612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1710841341
transform 1 0 532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1710841341
transform 1 0 644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1710841341
transform 1 0 620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1710841341
transform 1 0 596 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1710841341
transform 1 0 588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1710841341
transform 1 0 444 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1710841341
transform 1 0 2092 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1710841341
transform 1 0 2044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1710841341
transform 1 0 1980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1710841341
transform 1 0 1556 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1710841341
transform 1 0 1540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1710841341
transform 1 0 1356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1710841341
transform 1 0 2572 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1710841341
transform 1 0 2276 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1710841341
transform 1 0 2260 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1710841341
transform 1 0 2244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1710841341
transform 1 0 2020 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1710841341
transform 1 0 1828 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1710841341
transform 1 0 1700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1710841341
transform 1 0 1972 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1710841341
transform 1 0 1236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1710841341
transform 1 0 1196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1710841341
transform 1 0 1196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1710841341
transform 1 0 1188 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1710841341
transform 1 0 1164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1710841341
transform 1 0 996 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1710841341
transform 1 0 916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1710841341
transform 1 0 916 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1710841341
transform 1 0 900 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1710841341
transform 1 0 1116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1710841341
transform 1 0 1100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1710841341
transform 1 0 1572 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1710841341
transform 1 0 1548 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1710841341
transform 1 0 1340 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1710841341
transform 1 0 1148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1710841341
transform 1 0 1148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1710841341
transform 1 0 1148 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1710841341
transform 1 0 956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1710841341
transform 1 0 956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1710841341
transform 1 0 924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1710841341
transform 1 0 852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1710841341
transform 1 0 2100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1710841341
transform 1 0 2068 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1710841341
transform 1 0 2068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1710841341
transform 1 0 300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1710841341
transform 1 0 268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1710841341
transform 1 0 1036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1710841341
transform 1 0 932 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1710841341
transform 1 0 844 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1710841341
transform 1 0 1604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1710841341
transform 1 0 1276 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1710841341
transform 1 0 1220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1710841341
transform 1 0 1068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1710841341
transform 1 0 1060 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1710841341
transform 1 0 1012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1710841341
transform 1 0 812 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1710841341
transform 1 0 804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1710841341
transform 1 0 764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1710841341
transform 1 0 884 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1710841341
transform 1 0 804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1710841341
transform 1 0 740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1710841341
transform 1 0 2076 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1710841341
transform 1 0 1996 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1710841341
transform 1 0 1980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1710841341
transform 1 0 2004 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1710841341
transform 1 0 1900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1710841341
transform 1 0 1708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1710841341
transform 1 0 1620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1710841341
transform 1 0 1308 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1710841341
transform 1 0 1252 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1710841341
transform 1 0 644 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1710841341
transform 1 0 620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1710841341
transform 1 0 612 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1710841341
transform 1 0 588 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1710841341
transform 1 0 588 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1710841341
transform 1 0 1820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1710841341
transform 1 0 1636 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1710841341
transform 1 0 828 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1710841341
transform 1 0 564 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1710841341
transform 1 0 2004 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1710841341
transform 1 0 1924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1710841341
transform 1 0 1084 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1710841341
transform 1 0 996 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1710841341
transform 1 0 948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1710841341
transform 1 0 996 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1710841341
transform 1 0 892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1710841341
transform 1 0 796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1710841341
transform 1 0 2076 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1710841341
transform 1 0 2036 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1710841341
transform 1 0 1964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1710841341
transform 1 0 2140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1710841341
transform 1 0 2140 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1710841341
transform 1 0 2068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1710841341
transform 1 0 1004 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1710841341
transform 1 0 836 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1710841341
transform 1 0 796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1710841341
transform 1 0 1812 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1710841341
transform 1 0 1364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1710841341
transform 1 0 1316 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1710841341
transform 1 0 1204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1710841341
transform 1 0 1116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1710841341
transform 1 0 1076 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1710841341
transform 1 0 1076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1710841341
transform 1 0 948 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1710841341
transform 1 0 836 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1710841341
transform 1 0 732 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1710841341
transform 1 0 1660 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1710841341
transform 1 0 1300 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1710841341
transform 1 0 1260 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1710841341
transform 1 0 916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1710841341
transform 1 0 892 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1710841341
transform 1 0 764 0 1 1695
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1710841341
transform 1 0 764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1710841341
transform 1 0 756 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1710841341
transform 1 0 1076 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1710841341
transform 1 0 828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1710841341
transform 1 0 828 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1710841341
transform 1 0 604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1710841341
transform 1 0 596 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1710841341
transform 1 0 2116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1710841341
transform 1 0 2052 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1710841341
transform 1 0 1996 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1710841341
transform 1 0 1732 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1710841341
transform 1 0 1620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1710841341
transform 1 0 1620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1710841341
transform 1 0 2516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1710841341
transform 1 0 2508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1710841341
transform 1 0 2204 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1710841341
transform 1 0 2108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1710841341
transform 1 0 1956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1710841341
transform 1 0 1876 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1710841341
transform 1 0 980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1710841341
transform 1 0 964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1710841341
transform 1 0 1532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1710841341
transform 1 0 1500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1710841341
transform 1 0 1220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1710841341
transform 1 0 1188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1710841341
transform 1 0 1180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1710841341
transform 1 0 1180 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1710841341
transform 1 0 1580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1710841341
transform 1 0 1420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1710841341
transform 1 0 1348 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1710841341
transform 1 0 964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1710841341
transform 1 0 740 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1710841341
transform 1 0 2028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1710841341
transform 1 0 2028 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1710841341
transform 1 0 2020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1710841341
transform 1 0 1964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1710841341
transform 1 0 2156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1710841341
transform 1 0 2020 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1710841341
transform 1 0 1676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1710841341
transform 1 0 1588 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1710841341
transform 1 0 1452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1710841341
transform 1 0 1452 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1710841341
transform 1 0 364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1710841341
transform 1 0 348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1710841341
transform 1 0 284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1710841341
transform 1 0 268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1710841341
transform 1 0 244 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1710841341
transform 1 0 204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1710841341
transform 1 0 364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1710841341
transform 1 0 364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1710841341
transform 1 0 340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1710841341
transform 1 0 316 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1710841341
transform 1 0 300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1710841341
transform 1 0 300 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1710841341
transform 1 0 276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1710841341
transform 1 0 308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1710841341
transform 1 0 236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1710841341
transform 1 0 196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1710841341
transform 1 0 164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1710841341
transform 1 0 204 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1710841341
transform 1 0 164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1710841341
transform 1 0 436 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1710841341
transform 1 0 428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1710841341
transform 1 0 412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1710841341
transform 1 0 524 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1710841341
transform 1 0 524 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1710841341
transform 1 0 484 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1710841341
transform 1 0 484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1710841341
transform 1 0 396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1710841341
transform 1 0 356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1710841341
transform 1 0 356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1710841341
transform 1 0 260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1710841341
transform 1 0 260 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1710841341
transform 1 0 252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1710841341
transform 1 0 188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1710841341
transform 1 0 188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1710841341
transform 1 0 164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1710841341
transform 1 0 668 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1710841341
transform 1 0 660 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1710841341
transform 1 0 452 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1710841341
transform 1 0 524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1710841341
transform 1 0 500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1710841341
transform 1 0 444 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1710841341
transform 1 0 412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1710841341
transform 1 0 740 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1710841341
transform 1 0 740 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1710841341
transform 1 0 708 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1710841341
transform 1 0 548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1710841341
transform 1 0 556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1710841341
transform 1 0 548 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1710841341
transform 1 0 684 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1710841341
transform 1 0 684 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1710841341
transform 1 0 636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1710841341
transform 1 0 484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1710841341
transform 1 0 1124 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1710841341
transform 1 0 1060 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1710841341
transform 1 0 900 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1710841341
transform 1 0 764 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1710841341
transform 1 0 764 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1710841341
transform 1 0 788 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1710841341
transform 1 0 700 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1710841341
transform 1 0 716 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1710841341
transform 1 0 700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1710841341
transform 1 0 1236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1710841341
transform 1 0 1236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1710841341
transform 1 0 1116 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1710841341
transform 1 0 1100 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1710841341
transform 1 0 1084 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1710841341
transform 1 0 940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1710841341
transform 1 0 892 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1710841341
transform 1 0 1340 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1710841341
transform 1 0 1268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1710841341
transform 1 0 996 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1710841341
transform 1 0 996 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1710841341
transform 1 0 348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1710841341
transform 1 0 340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1710841341
transform 1 0 380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1710841341
transform 1 0 372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1710841341
transform 1 0 588 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1710841341
transform 1 0 532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1710841341
transform 1 0 532 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1710841341
transform 1 0 684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1710841341
transform 1 0 668 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1710841341
transform 1 0 668 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1710841341
transform 1 0 612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1710841341
transform 1 0 604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1710841341
transform 1 0 436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1710841341
transform 1 0 436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1710841341
transform 1 0 836 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1710841341
transform 1 0 812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1710841341
transform 1 0 812 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1710841341
transform 1 0 1092 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1710841341
transform 1 0 1060 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1710841341
transform 1 0 1060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1710841341
transform 1 0 1116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1710841341
transform 1 0 1052 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1710841341
transform 1 0 1220 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1710841341
transform 1 0 1140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1710841341
transform 1 0 1284 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1710841341
transform 1 0 1284 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1710841341
transform 1 0 1268 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1710841341
transform 1 0 1244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1710841341
transform 1 0 1244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1710841341
transform 1 0 1500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1710841341
transform 1 0 1500 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1710841341
transform 1 0 1396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1710841341
transform 1 0 1396 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1710841341
transform 1 0 1708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1710841341
transform 1 0 1700 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1710841341
transform 1 0 1612 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1710841341
transform 1 0 1516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1710841341
transform 1 0 1828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1710841341
transform 1 0 1796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1710841341
transform 1 0 1596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1710841341
transform 1 0 1572 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1710841341
transform 1 0 1796 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1710841341
transform 1 0 1692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1710841341
transform 1 0 1692 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1710841341
transform 1 0 1676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1710841341
transform 1 0 1548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1710841341
transform 1 0 1932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1710841341
transform 1 0 1892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1710841341
transform 1 0 1956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1710841341
transform 1 0 1956 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1710841341
transform 1 0 1892 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1710841341
transform 1 0 1828 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1710841341
transform 1 0 1820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1710841341
transform 1 0 1660 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1710841341
transform 1 0 1660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1710841341
transform 1 0 1628 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1710841341
transform 1 0 1484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1710841341
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1710841341
transform 1 0 1924 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1710841341
transform 1 0 1876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1710841341
transform 1 0 1940 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1710841341
transform 1 0 1516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1710841341
transform 1 0 1428 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1710841341
transform 1 0 2348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1710841341
transform 1 0 2172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1710841341
transform 1 0 2172 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1710841341
transform 1 0 2164 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1710841341
transform 1 0 2404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1710841341
transform 1 0 2372 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1710841341
transform 1 0 2340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1710841341
transform 1 0 2300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1710841341
transform 1 0 2164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1710841341
transform 1 0 2124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1710841341
transform 1 0 2252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1710841341
transform 1 0 2092 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1710841341
transform 1 0 2076 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1710841341
transform 1 0 2292 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1710841341
transform 1 0 2268 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1710841341
transform 1 0 2268 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1710841341
transform 1 0 2228 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1710841341
transform 1 0 2212 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1710841341
transform 1 0 2388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1710841341
transform 1 0 2356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1710841341
transform 1 0 2540 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1710841341
transform 1 0 2508 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1710841341
transform 1 0 2508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1710841341
transform 1 0 2148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1710841341
transform 1 0 2060 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1710841341
transform 1 0 2044 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1710841341
transform 1 0 2172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1710841341
transform 1 0 2140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1710841341
transform 1 0 2596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1710841341
transform 1 0 2540 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1710841341
transform 1 0 2540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1710841341
transform 1 0 2444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1710841341
transform 1 0 2316 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1710841341
transform 1 0 2220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1710841341
transform 1 0 2156 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1710841341
transform 1 0 2436 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1710841341
transform 1 0 2396 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1710841341
transform 1 0 2668 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1710841341
transform 1 0 2668 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1710841341
transform 1 0 2452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1710841341
transform 1 0 2452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1710841341
transform 1 0 2164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1710841341
transform 1 0 2148 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1710841341
transform 1 0 2316 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1710841341
transform 1 0 2284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1710841341
transform 1 0 2228 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1710841341
transform 1 0 2172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1710841341
transform 1 0 2020 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1710841341
transform 1 0 2324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1710841341
transform 1 0 2284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1710841341
transform 1 0 2516 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1710841341
transform 1 0 2484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1710841341
transform 1 0 2300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1710841341
transform 1 0 2292 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1710841341
transform 1 0 2148 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1710841341
transform 1 0 1820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1710841341
transform 1 0 1820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1710841341
transform 1 0 1756 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1710841341
transform 1 0 1724 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1710841341
transform 1 0 1716 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1710841341
transform 1 0 1828 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1710841341
transform 1 0 1820 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1710841341
transform 1 0 2084 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1710841341
transform 1 0 1724 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1710841341
transform 1 0 1724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1710841341
transform 1 0 2452 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1710841341
transform 1 0 2388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1710841341
transform 1 0 2540 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1710841341
transform 1 0 2524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1710841341
transform 1 0 2588 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1710841341
transform 1 0 2572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1710841341
transform 1 0 2556 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1710841341
transform 1 0 2396 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1710841341
transform 1 0 2396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1710841341
transform 1 0 2356 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1710841341
transform 1 0 2348 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1710841341
transform 1 0 2380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1710841341
transform 1 0 2380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1710841341
transform 1 0 2596 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1710841341
transform 1 0 2564 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1710841341
transform 1 0 2284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1710841341
transform 1 0 2268 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1710841341
transform 1 0 2228 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1710841341
transform 1 0 2212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1710841341
transform 1 0 2196 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1710841341
transform 1 0 2156 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1710841341
transform 1 0 2140 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1710841341
transform 1 0 2308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1710841341
transform 1 0 2308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1710841341
transform 1 0 2372 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1710841341
transform 1 0 2340 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1710841341
transform 1 0 1996 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1710841341
transform 1 0 1972 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1710841341
transform 1 0 1948 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1710841341
transform 1 0 1924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1710841341
transform 1 0 1844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1710841341
transform 1 0 1844 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1710841341
transform 1 0 1828 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1710841341
transform 1 0 1988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1710841341
transform 1 0 1948 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1710841341
transform 1 0 2116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1710841341
transform 1 0 1988 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1710841341
transform 1 0 2044 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1710841341
transform 1 0 1940 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1710841341
transform 1 0 1684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1710841341
transform 1 0 1652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1710841341
transform 1 0 1548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1710841341
transform 1 0 1548 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1710841341
transform 1 0 1540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1710841341
transform 1 0 1724 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1710841341
transform 1 0 1708 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1710841341
transform 1 0 1748 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1710841341
transform 1 0 1660 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1710841341
transform 1 0 1796 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1710841341
transform 1 0 1756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1710841341
transform 1 0 844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1710841341
transform 1 0 844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1710841341
transform 1 0 788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1710841341
transform 1 0 772 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1710841341
transform 1 0 300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1710841341
transform 1 0 276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1710841341
transform 1 0 1524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1710841341
transform 1 0 1508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1710841341
transform 1 0 1972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1710841341
transform 1 0 1956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1710841341
transform 1 0 2500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1710841341
transform 1 0 2484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1710841341
transform 1 0 2596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1710841341
transform 1 0 2580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1710841341
transform 1 0 2604 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1710841341
transform 1 0 2588 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1710841341
transform 1 0 1172 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1710841341
transform 1 0 1124 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1710841341
transform 1 0 1084 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1710841341
transform 1 0 700 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1710841341
transform 1 0 692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1710841341
transform 1 0 564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1710841341
transform 1 0 476 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1710841341
transform 1 0 1468 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1710841341
transform 1 0 1340 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1710841341
transform 1 0 1340 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1710841341
transform 1 0 1292 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1710841341
transform 1 0 1284 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1710841341
transform 1 0 1268 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1710841341
transform 1 0 1212 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1710841341
transform 1 0 1108 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1710841341
transform 1 0 908 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1710841341
transform 1 0 892 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1710841341
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1710841341
transform 1 0 412 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1710841341
transform 1 0 396 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1710841341
transform 1 0 396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1710841341
transform 1 0 372 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1710841341
transform 1 0 332 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1710841341
transform 1 0 164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1710841341
transform 1 0 156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1710841341
transform 1 0 140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1710841341
transform 1 0 132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1710841341
transform 1 0 164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1710841341
transform 1 0 124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1710841341
transform 1 0 164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1710841341
transform 1 0 108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1710841341
transform 1 0 124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1710841341
transform 1 0 124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1710841341
transform 1 0 756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1710841341
transform 1 0 756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1710841341
transform 1 0 1004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1710841341
transform 1 0 956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1710841341
transform 1 0 2380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1710841341
transform 1 0 2300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1710841341
transform 1 0 2332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1710841341
transform 1 0 2284 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1710841341
transform 1 0 1484 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1710841341
transform 1 0 772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1710841341
transform 1 0 508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1710841341
transform 1 0 484 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1710841341
transform 1 0 2532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1710841341
transform 1 0 2516 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1710841341
transform 1 0 2172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1710841341
transform 1 0 1380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1710841341
transform 1 0 1356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1710841341
transform 1 0 1004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1710841341
transform 1 0 1540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1710841341
transform 1 0 1468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1710841341
transform 1 0 2556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1710841341
transform 1 0 2540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1710841341
transform 1 0 1468 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1710841341
transform 1 0 1396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1710841341
transform 1 0 1220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1710841341
transform 1 0 1156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1710841341
transform 1 0 1020 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1710841341
transform 1 0 980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1710841341
transform 1 0 852 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1710841341
transform 1 0 812 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1710841341
transform 1 0 164 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1710841341
transform 1 0 84 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1710841341
transform 1 0 308 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1710841341
transform 1 0 244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1710841341
transform 1 0 284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1710841341
transform 1 0 236 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1710841341
transform 1 0 268 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1710841341
transform 1 0 252 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1710841341
transform 1 0 244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1710841341
transform 1 0 188 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1710841341
transform 1 0 140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1710841341
transform 1 0 124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1710841341
transform 1 0 116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1710841341
transform 1 0 76 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1710841341
transform 1 0 460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1710841341
transform 1 0 372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1710841341
transform 1 0 348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1710841341
transform 1 0 372 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1710841341
transform 1 0 324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1710841341
transform 1 0 324 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1710841341
transform 1 0 292 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1710841341
transform 1 0 292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1710841341
transform 1 0 284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1710841341
transform 1 0 252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1710841341
transform 1 0 252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1710841341
transform 1 0 244 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1710841341
transform 1 0 2628 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1710841341
transform 1 0 2556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1710841341
transform 1 0 2540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1710841341
transform 1 0 2492 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1710841341
transform 1 0 2492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1710841341
transform 1 0 2356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1710841341
transform 1 0 2284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1710841341
transform 1 0 2244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1710841341
transform 1 0 2076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1710841341
transform 1 0 1908 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1710841341
transform 1 0 1900 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1710841341
transform 1 0 1884 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1710841341
transform 1 0 1788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1710841341
transform 1 0 1756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1710841341
transform 1 0 1444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1710841341
transform 1 0 1332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1710841341
transform 1 0 1284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1710841341
transform 1 0 908 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1710841341
transform 1 0 668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1710841341
transform 1 0 636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1710841341
transform 1 0 500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1710841341
transform 1 0 316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1710841341
transform 1 0 68 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1710841341
transform 1 0 68 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1710841341
transform 1 0 68 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1710841341
transform 1 0 2108 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1710841341
transform 1 0 2076 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1710841341
transform 1 0 2068 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1710841341
transform 1 0 2068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1710841341
transform 1 0 1996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1710841341
transform 1 0 1900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1710841341
transform 1 0 1596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1710841341
transform 1 0 1500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1710841341
transform 1 0 1212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1710841341
transform 1 0 1140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1710841341
transform 1 0 1076 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1710841341
transform 1 0 876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1710841341
transform 1 0 756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1710841341
transform 1 0 716 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1710841341
transform 1 0 676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1710841341
transform 1 0 628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1710841341
transform 1 0 628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1710841341
transform 1 0 2620 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1710841341
transform 1 0 2580 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1710841341
transform 1 0 2540 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1710841341
transform 1 0 2516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1710841341
transform 1 0 2252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1710841341
transform 1 0 2036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1710841341
transform 1 0 2036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1710841341
transform 1 0 1948 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1710841341
transform 1 0 1948 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1710841341
transform 1 0 1908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1710841341
transform 1 0 1572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1710841341
transform 1 0 1556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1710841341
transform 1 0 1476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1710841341
transform 1 0 1252 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1710841341
transform 1 0 1172 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1710841341
transform 1 0 1084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1710841341
transform 1 0 1052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1710841341
transform 1 0 852 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1710841341
transform 1 0 2252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1710841341
transform 1 0 2172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1710841341
transform 1 0 2092 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1710841341
transform 1 0 2076 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1710841341
transform 1 0 2060 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1710841341
transform 1 0 2052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1710841341
transform 1 0 1924 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1710841341
transform 1 0 1500 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1710841341
transform 1 0 996 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1710841341
transform 1 0 828 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1710841341
transform 1 0 692 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1710841341
transform 1 0 524 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1710841341
transform 1 0 476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1710841341
transform 1 0 428 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1710841341
transform 1 0 348 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1710841341
transform 1 0 324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1710841341
transform 1 0 316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1710841341
transform 1 0 308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1710841341
transform 1 0 2628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1710841341
transform 1 0 2596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1710841341
transform 1 0 2572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1710841341
transform 1 0 2380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1710841341
transform 1 0 2364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1710841341
transform 1 0 2348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1710841341
transform 1 0 2020 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1710841341
transform 1 0 1804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1710841341
transform 1 0 1796 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1710841341
transform 1 0 1796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1710841341
transform 1 0 1660 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1710841341
transform 1 0 1348 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1710841341
transform 1 0 1204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1710841341
transform 1 0 1164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1710841341
transform 1 0 1156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1710841341
transform 1 0 1116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1710841341
transform 1 0 1004 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1710841341
transform 1 0 932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1710841341
transform 1 0 644 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1710841341
transform 1 0 548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1710841341
transform 1 0 412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1710841341
transform 1 0 332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1710841341
transform 1 0 212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1710841341
transform 1 0 196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1710841341
transform 1 0 196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1710841341
transform 1 0 2572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1710841341
transform 1 0 2516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1710841341
transform 1 0 2508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1710841341
transform 1 0 2332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1710841341
transform 1 0 2300 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1710841341
transform 1 0 2204 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1710841341
transform 1 0 1852 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1710841341
transform 1 0 1724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1710841341
transform 1 0 1396 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1710841341
transform 1 0 1340 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1710841341
transform 1 0 1284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1710841341
transform 1 0 1204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1710841341
transform 1 0 1004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1710841341
transform 1 0 908 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1710841341
transform 1 0 868 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1710841341
transform 1 0 484 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1710841341
transform 1 0 2676 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1710841341
transform 1 0 2556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1710841341
transform 1 0 2468 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1710841341
transform 1 0 2428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1710841341
transform 1 0 2372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1710841341
transform 1 0 2052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1710841341
transform 1 0 1988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1710841341
transform 1 0 1652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1710841341
transform 1 0 1556 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1710841341
transform 1 0 1540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1710841341
transform 1 0 1212 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1710841341
transform 1 0 1140 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1710841341
transform 1 0 932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1710841341
transform 1 0 708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1710841341
transform 1 0 1668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1710841341
transform 1 0 1612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1710841341
transform 1 0 1612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1710841341
transform 1 0 1372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1710841341
transform 1 0 1156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1710841341
transform 1 0 932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1710841341
transform 1 0 836 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1710841341
transform 1 0 812 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1710841341
transform 1 0 764 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1710841341
transform 1 0 764 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1710841341
transform 1 0 2100 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1710841341
transform 1 0 2100 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1710841341
transform 1 0 2092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1710841341
transform 1 0 2060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1710841341
transform 1 0 2052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1710841341
transform 1 0 2052 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1710841341
transform 1 0 1636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1710841341
transform 1 0 1436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1710841341
transform 1 0 1244 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1710841341
transform 1 0 1060 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1710841341
transform 1 0 988 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1710841341
transform 1 0 948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1710841341
transform 1 0 940 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1710841341
transform 1 0 900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1710841341
transform 1 0 876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1710841341
transform 1 0 820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1710841341
transform 1 0 788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1710841341
transform 1 0 2236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1710841341
transform 1 0 2164 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1710841341
transform 1 0 2124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1710841341
transform 1 0 2084 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1710841341
transform 1 0 1492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1710841341
transform 1 0 1236 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1710841341
transform 1 0 1196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1710841341
transform 1 0 948 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1710841341
transform 1 0 860 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1710841341
transform 1 0 2148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1710841341
transform 1 0 2148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1710841341
transform 1 0 2132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1710841341
transform 1 0 2100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1710841341
transform 1 0 2084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1710841341
transform 1 0 2036 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1710841341
transform 1 0 2028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1710841341
transform 1 0 1916 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1710841341
transform 1 0 1604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1710841341
transform 1 0 1364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1710841341
transform 1 0 1220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1710841341
transform 1 0 972 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1710841341
transform 1 0 900 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1710841341
transform 1 0 868 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1710841341
transform 1 0 836 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1710841341
transform 1 0 836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1710841341
transform 1 0 764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1710841341
transform 1 0 708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1710841341
transform 1 0 2612 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1710841341
transform 1 0 2468 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1710841341
transform 1 0 2460 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1710841341
transform 1 0 2412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1710841341
transform 1 0 2100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1710841341
transform 1 0 1380 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1710841341
transform 1 0 1380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1710841341
transform 1 0 1236 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1710841341
transform 1 0 1236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1710841341
transform 1 0 1908 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1710841341
transform 1 0 1844 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1710841341
transform 1 0 1836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1710841341
transform 1 0 1820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1710841341
transform 1 0 1780 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1710841341
transform 1 0 1772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1710841341
transform 1 0 1772 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1710841341
transform 1 0 1756 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1710841341
transform 1 0 1692 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1710841341
transform 1 0 1692 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1710841341
transform 1 0 2092 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1710841341
transform 1 0 1948 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1710841341
transform 1 0 1364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1710841341
transform 1 0 1180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1710841341
transform 1 0 2308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1710841341
transform 1 0 1916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1710841341
transform 1 0 1380 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1710841341
transform 1 0 1372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1710841341
transform 1 0 2532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1710841341
transform 1 0 2508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1710841341
transform 1 0 2460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1710841341
transform 1 0 1236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1710841341
transform 1 0 652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1710841341
transform 1 0 2460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1710841341
transform 1 0 1804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1710841341
transform 1 0 1740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1710841341
transform 1 0 1316 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1710841341
transform 1 0 1308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1710841341
transform 1 0 2324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1710841341
transform 1 0 2252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1710841341
transform 1 0 1316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1710841341
transform 1 0 404 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1710841341
transform 1 0 364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1710841341
transform 1 0 2052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1710841341
transform 1 0 1924 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1710841341
transform 1 0 1772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1710841341
transform 1 0 1388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1710841341
transform 1 0 612 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1710841341
transform 1 0 1244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1710841341
transform 1 0 1220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1710841341
transform 1 0 1348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1710841341
transform 1 0 1292 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1710841341
transform 1 0 2396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1710841341
transform 1 0 2308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1710841341
transform 1 0 2300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1710841341
transform 1 0 2164 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1710841341
transform 1 0 2156 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1710841341
transform 1 0 2132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1710841341
transform 1 0 2108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1710841341
transform 1 0 2028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1710841341
transform 1 0 1772 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1710841341
transform 1 0 1548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1710841341
transform 1 0 1492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1710841341
transform 1 0 1476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1710841341
transform 1 0 540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1710841341
transform 1 0 420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1710841341
transform 1 0 2428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1710841341
transform 1 0 2164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1710841341
transform 1 0 1844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1710841341
transform 1 0 1180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1710841341
transform 1 0 1108 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1710841341
transform 1 0 1484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1710841341
transform 1 0 1228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1710841341
transform 1 0 1204 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1710841341
transform 1 0 708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1710841341
transform 1 0 348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1710841341
transform 1 0 2372 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1710841341
transform 1 0 2356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1710841341
transform 1 0 2132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1710841341
transform 1 0 1172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1710841341
transform 1 0 964 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1710841341
transform 1 0 1188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1710841341
transform 1 0 1180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1710841341
transform 1 0 1164 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1710841341
transform 1 0 1156 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1710841341
transform 1 0 2452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1710841341
transform 1 0 2404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1710841341
transform 1 0 2404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1710841341
transform 1 0 2348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1710841341
transform 1 0 2332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1710841341
transform 1 0 2260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1710841341
transform 1 0 2148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1710841341
transform 1 0 2068 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1710841341
transform 1 0 2012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1710841341
transform 1 0 1828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1710841341
transform 1 0 1828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1710841341
transform 1 0 1812 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1710841341
transform 1 0 1780 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1710841341
transform 1 0 1636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1710841341
transform 1 0 1476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1710841341
transform 1 0 1196 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1710841341
transform 1 0 1076 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1710841341
transform 1 0 548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1710841341
transform 1 0 548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1710841341
transform 1 0 1884 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1710841341
transform 1 0 1804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1710841341
transform 1 0 1788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1710841341
transform 1 0 1708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1710841341
transform 1 0 1668 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1710841341
transform 1 0 1668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1710841341
transform 1 0 1620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1710841341
transform 1 0 1620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1710841341
transform 1 0 1620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1710841341
transform 1 0 1572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1710841341
transform 1 0 1572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1710841341
transform 1 0 1164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1710841341
transform 1 0 1068 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1710841341
transform 1 0 1068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1710841341
transform 1 0 1012 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1710841341
transform 1 0 1012 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1710841341
transform 1 0 940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1710841341
transform 1 0 684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1710841341
transform 1 0 684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1710841341
transform 1 0 636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1710841341
transform 1 0 620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1710841341
transform 1 0 612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1710841341
transform 1 0 612 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1710841341
transform 1 0 572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1710841341
transform 1 0 2476 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1710841341
transform 1 0 2476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1710841341
transform 1 0 2436 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1710841341
transform 1 0 2388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1710841341
transform 1 0 2340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1710841341
transform 1 0 2332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1710841341
transform 1 0 2268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1710841341
transform 1 0 2068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1710841341
transform 1 0 2012 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1710841341
transform 1 0 1980 0 1 1085
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1710841341
transform 1 0 1972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1710841341
transform 1 0 1972 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1710841341
transform 1 0 1796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1710841341
transform 1 0 1780 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1710841341
transform 1 0 1764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1710841341
transform 1 0 1620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1710841341
transform 1 0 1388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1710841341
transform 1 0 1196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1710841341
transform 1 0 628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1710841341
transform 1 0 532 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1710841341
transform 1 0 524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1710841341
transform 1 0 508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1710841341
transform 1 0 1692 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1710841341
transform 1 0 1684 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1710841341
transform 1 0 1620 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1710841341
transform 1 0 1580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1710841341
transform 1 0 1356 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1710841341
transform 1 0 876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1710841341
transform 1 0 876 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1710841341
transform 1 0 836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1710841341
transform 1 0 812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1710841341
transform 1 0 804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1710841341
transform 1 0 2644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1710841341
transform 1 0 2612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1710841341
transform 1 0 2588 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1710841341
transform 1 0 2396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1710841341
transform 1 0 2380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1710841341
transform 1 0 2364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1710841341
transform 1 0 2036 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1710841341
transform 1 0 1820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1710841341
transform 1 0 1812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1710841341
transform 1 0 1812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1710841341
transform 1 0 1676 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1710841341
transform 1 0 1468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1710841341
transform 1 0 1308 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1710841341
transform 1 0 1308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1710841341
transform 1 0 1284 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1710841341
transform 1 0 1228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1710841341
transform 1 0 1172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1710841341
transform 1 0 948 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1710841341
transform 1 0 924 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1710841341
transform 1 0 524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1710841341
transform 1 0 516 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1710841341
transform 1 0 436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1710841341
transform 1 0 396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1710841341
transform 1 0 364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1710841341
transform 1 0 1636 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1710841341
transform 1 0 1540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1710841341
transform 1 0 1540 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1710841341
transform 1 0 1484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1710841341
transform 1 0 1284 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1710841341
transform 1 0 916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1710841341
transform 1 0 796 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1710841341
transform 1 0 748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1710841341
transform 1 0 716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1710841341
transform 1 0 716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1710841341
transform 1 0 700 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1710841341
transform 1 0 2204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1710841341
transform 1 0 1668 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1710841341
transform 1 0 1012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1710841341
transform 1 0 964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1710841341
transform 1 0 740 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1710841341
transform 1 0 660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1710841341
transform 1 0 548 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1710841341
transform 1 0 2308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1710841341
transform 1 0 2244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1710841341
transform 1 0 2236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1710841341
transform 1 0 1828 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1710841341
transform 1 0 908 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1710841341
transform 1 0 908 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1710841341
transform 1 0 892 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1710841341
transform 1 0 892 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1710841341
transform 1 0 876 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1710841341
transform 1 0 740 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1710841341
transform 1 0 2372 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1710841341
transform 1 0 2332 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1710841341
transform 1 0 2324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1710841341
transform 1 0 2300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1710841341
transform 1 0 2220 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1710841341
transform 1 0 2188 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1710841341
transform 1 0 2172 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1710841341
transform 1 0 2148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1710841341
transform 1 0 2124 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1710841341
transform 1 0 1916 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1710841341
transform 1 0 1564 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1710841341
transform 1 0 1444 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1710841341
transform 1 0 1052 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1710841341
transform 1 0 732 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1710841341
transform 1 0 716 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1710841341
transform 1 0 500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1710841341
transform 1 0 460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1710841341
transform 1 0 340 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1710841341
transform 1 0 292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1710841341
transform 1 0 276 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1710841341
transform 1 0 244 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1710841341
transform 1 0 2620 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1710841341
transform 1 0 2588 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1710841341
transform 1 0 2588 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1710841341
transform 1 0 2588 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1710841341
transform 1 0 2588 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1710841341
transform 1 0 2588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1710841341
transform 1 0 2588 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1710841341
transform 1 0 2484 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1710841341
transform 1 0 2460 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1710841341
transform 1 0 2452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1710841341
transform 1 0 2444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1710841341
transform 1 0 2420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1710841341
transform 1 0 2420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1710841341
transform 1 0 2068 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1710841341
transform 1 0 2004 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1710841341
transform 1 0 1932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1710841341
transform 1 0 1852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1710841341
transform 1 0 1844 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1710841341
transform 1 0 1636 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1710841341
transform 1 0 1628 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1710841341
transform 1 0 1444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1710841341
transform 1 0 1108 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1710841341
transform 1 0 1068 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1710841341
transform 1 0 996 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1710841341
transform 1 0 988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1710841341
transform 1 0 828 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1710841341
transform 1 0 740 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1710841341
transform 1 0 668 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1710841341
transform 1 0 660 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1710841341
transform 1 0 540 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1710841341
transform 1 0 492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1710841341
transform 1 0 412 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1710841341
transform 1 0 372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1710841341
transform 1 0 340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1710841341
transform 1 0 292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1710841341
transform 1 0 252 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1710841341
transform 1 0 172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1710841341
transform 1 0 140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1710841341
transform 1 0 132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1710841341
transform 1 0 124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1710841341
transform 1 0 100 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1710841341
transform 1 0 84 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1710841341
transform 1 0 2628 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1710841341
transform 1 0 2596 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1710841341
transform 1 0 2660 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1710841341
transform 1 0 2660 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1710841341
transform 1 0 2660 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1710841341
transform 1 0 2612 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1710841341
transform 1 0 2564 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1710841341
transform 1 0 2548 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1710841341
transform 1 0 2500 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1710841341
transform 1 0 2500 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1710841341
transform 1 0 2484 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1710841341
transform 1 0 2428 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1710841341
transform 1 0 2388 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1710841341
transform 1 0 2036 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1710841341
transform 1 0 1940 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1710841341
transform 1 0 1916 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1710841341
transform 1 0 1900 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1710841341
transform 1 0 1788 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1710841341
transform 1 0 1772 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1710841341
transform 1 0 1596 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1710841341
transform 1 0 1196 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1710841341
transform 1 0 1068 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1710841341
transform 1 0 1044 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1710841341
transform 1 0 780 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1710841341
transform 1 0 764 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1710841341
transform 1 0 636 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1710841341
transform 1 0 540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1710841341
transform 1 0 524 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1710841341
transform 1 0 404 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1710841341
transform 1 0 380 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1710841341
transform 1 0 380 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1710841341
transform 1 0 364 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1710841341
transform 1 0 252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1710841341
transform 1 0 220 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1710841341
transform 1 0 204 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1710841341
transform 1 0 1300 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1710841341
transform 1 0 1172 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1710841341
transform 1 0 988 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1710841341
transform 1 0 892 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1710841341
transform 1 0 476 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1710841341
transform 1 0 436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1710841341
transform 1 0 228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1710841341
transform 1 0 148 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1710841341
transform 1 0 132 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1710841341
transform 1 0 116 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1710841341
transform 1 0 92 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1710841341
transform 1 0 668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1710841341
transform 1 0 588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1710841341
transform 1 0 572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1710841341
transform 1 0 564 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1710841341
transform 1 0 548 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1710841341
transform 1 0 468 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1710841341
transform 1 0 452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1710841341
transform 1 0 420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1710841341
transform 1 0 404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1710841341
transform 1 0 396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1710841341
transform 1 0 372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1710841341
transform 1 0 340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1710841341
transform 1 0 308 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1710841341
transform 1 0 268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1710841341
transform 1 0 268 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1710841341
transform 1 0 260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1710841341
transform 1 0 228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1710841341
transform 1 0 372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1710841341
transform 1 0 252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1710841341
transform 1 0 556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1710841341
transform 1 0 556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1710841341
transform 1 0 2420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1710841341
transform 1 0 2420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1710841341
transform 1 0 2348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1710841341
transform 1 0 2324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1710841341
transform 1 0 1764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1710841341
transform 1 0 1724 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1710841341
transform 1 0 1828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1710841341
transform 1 0 1788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1710841341
transform 1 0 2468 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1710841341
transform 1 0 2420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1710841341
transform 1 0 996 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1710841341
transform 1 0 932 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1710841341
transform 1 0 828 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1710841341
transform 1 0 2188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1710841341
transform 1 0 2156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1710841341
transform 1 0 2124 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1710841341
transform 1 0 1668 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1710841341
transform 1 0 1636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1710841341
transform 1 0 1572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1710841341
transform 1 0 332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1710841341
transform 1 0 300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1710841341
transform 1 0 2284 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1710841341
transform 1 0 2276 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1710841341
transform 1 0 2220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1710841341
transform 1 0 2076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1710841341
transform 1 0 1964 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1710841341
transform 1 0 1516 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1710841341
transform 1 0 1428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1710841341
transform 1 0 2092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1710841341
transform 1 0 1988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1710841341
transform 1 0 1892 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1710841341
transform 1 0 1876 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1710841341
transform 1 0 1548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1710841341
transform 1 0 1316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1710841341
transform 1 0 1220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1710841341
transform 1 0 1212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1710841341
transform 1 0 1132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1710841341
transform 1 0 868 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1710841341
transform 1 0 1660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1710841341
transform 1 0 1476 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1710841341
transform 1 0 1252 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1710841341
transform 1 0 996 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1710841341
transform 1 0 1220 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1710841341
transform 1 0 1164 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1710841341
transform 1 0 964 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1710841341
transform 1 0 948 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1710841341
transform 1 0 916 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1710841341
transform 1 0 804 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1710841341
transform 1 0 724 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1710841341
transform 1 0 716 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1710841341
transform 1 0 652 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1710841341
transform 1 0 588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1710841341
transform 1 0 564 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1710841341
transform 1 0 1972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1710841341
transform 1 0 1924 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1710841341
transform 1 0 1572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1710841341
transform 1 0 1524 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1710841341
transform 1 0 1524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1710841341
transform 1 0 1524 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1710841341
transform 1 0 1300 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1710841341
transform 1 0 1260 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1710841341
transform 1 0 1244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1710841341
transform 1 0 1228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1710841341
transform 1 0 1172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1710841341
transform 1 0 660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1710841341
transform 1 0 1972 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1710841341
transform 1 0 1964 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1710841341
transform 1 0 1956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1710841341
transform 1 0 1876 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1710841341
transform 1 0 1796 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1710841341
transform 1 0 1788 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1710841341
transform 1 0 1764 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1710841341
transform 1 0 1660 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1710841341
transform 1 0 1660 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1710841341
transform 1 0 1612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1710841341
transform 1 0 1556 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1710841341
transform 1 0 724 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1710841341
transform 1 0 1836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1710841341
transform 1 0 1644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1710841341
transform 1 0 1548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1710841341
transform 1 0 908 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1710841341
transform 1 0 852 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1710841341
transform 1 0 820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1710841341
transform 1 0 748 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1710841341
transform 1 0 724 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1710841341
transform 1 0 692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1710841341
transform 1 0 676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1710841341
transform 1 0 116 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1710841341
transform 1 0 116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1710841341
transform 1 0 108 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1710841341
transform 1 0 196 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1710841341
transform 1 0 172 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1710841341
transform 1 0 148 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1710841341
transform 1 0 148 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1710841341
transform 1 0 308 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1710841341
transform 1 0 292 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1710841341
transform 1 0 212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1710841341
transform 1 0 220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1710841341
transform 1 0 148 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1710841341
transform 1 0 276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1710841341
transform 1 0 188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1710841341
transform 1 0 196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1710841341
transform 1 0 156 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1710841341
transform 1 0 188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1710841341
transform 1 0 148 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1710841341
transform 1 0 220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1710841341
transform 1 0 140 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1710841341
transform 1 0 220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1710841341
transform 1 0 132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1710841341
transform 1 0 612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1710841341
transform 1 0 268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1710841341
transform 1 0 364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1710841341
transform 1 0 348 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1710841341
transform 1 0 300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1710841341
transform 1 0 284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1710841341
transform 1 0 396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1710841341
transform 1 0 372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1710841341
transform 1 0 292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1710841341
transform 1 0 292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1710841341
transform 1 0 596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1710841341
transform 1 0 500 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1710841341
transform 1 0 444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1710841341
transform 1 0 436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1710841341
transform 1 0 1436 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1710841341
transform 1 0 1364 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1710841341
transform 1 0 1364 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1710841341
transform 1 0 1364 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1710841341
transform 1 0 1364 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1710841341
transform 1 0 1348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1710841341
transform 1 0 668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1710841341
transform 1 0 532 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1710841341
transform 1 0 556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1710841341
transform 1 0 540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1710841341
transform 1 0 452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1710841341
transform 1 0 452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1710841341
transform 1 0 460 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1710841341
transform 1 0 420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1710841341
transform 1 0 220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1710841341
transform 1 0 180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1710841341
transform 1 0 172 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1710841341
transform 1 0 132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1710841341
transform 1 0 756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1710841341
transform 1 0 716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1710841341
transform 1 0 628 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1710841341
transform 1 0 588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1710841341
transform 1 0 1756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1710841341
transform 1 0 1676 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1710841341
transform 1 0 2092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1710841341
transform 1 0 2052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1710841341
transform 1 0 2444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1710841341
transform 1 0 2404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1710841341
transform 1 0 2660 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1710841341
transform 1 0 2636 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1710841341
transform 1 0 2676 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1710841341
transform 1 0 2636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1710841341
transform 1 0 1956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1710841341
transform 1 0 1916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1710841341
transform 1 0 2668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1710841341
transform 1 0 2636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1710841341
transform 1 0 2612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1710841341
transform 1 0 2556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1710841341
transform 1 0 2612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1710841341
transform 1 0 2564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1710841341
transform 1 0 2620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1710841341
transform 1 0 2620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1710841341
transform 1 0 2508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1710841341
transform 1 0 2508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1710841341
transform 1 0 2476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1710841341
transform 1 0 2468 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1710841341
transform 1 0 2484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1710841341
transform 1 0 2444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1710841341
transform 1 0 1908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1710841341
transform 1 0 1900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1710841341
transform 1 0 2028 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1710841341
transform 1 0 1972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1710841341
transform 1 0 1868 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1710841341
transform 1 0 1796 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1710841341
transform 1 0 1660 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1710841341
transform 1 0 1620 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1710841341
transform 1 0 1196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1710841341
transform 1 0 1116 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1710841341
transform 1 0 1044 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1710841341
transform 1 0 788 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1710841341
transform 1 0 380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1710841341
transform 1 0 300 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1710841341
transform 1 0 316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1710841341
transform 1 0 220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1710841341
transform 1 0 1068 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1710841341
transform 1 0 1036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1710841341
transform 1 0 772 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1710841341
transform 1 0 708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1710841341
transform 1 0 524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1710841341
transform 1 0 388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1710841341
transform 1 0 388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1710841341
transform 1 0 340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1710841341
transform 1 0 732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1710841341
transform 1 0 260 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1710841341
transform 1 0 1660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1710841341
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1710841341
transform 1 0 1972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1710841341
transform 1 0 1964 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1710841341
transform 1 0 2532 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1710841341
transform 1 0 2516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1710841341
transform 1 0 2564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1710841341
transform 1 0 2092 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1710841341
transform 1 0 2524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1710841341
transform 1 0 2164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1710841341
transform 1 0 2572 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1710841341
transform 1 0 2164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1710841341
transform 1 0 1412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1710841341
transform 1 0 1364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1710841341
transform 1 0 1244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1710841341
transform 1 0 1244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1710841341
transform 1 0 1140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1710841341
transform 1 0 1092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1710841341
transform 1 0 940 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1710841341
transform 1 0 924 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1710841341
transform 1 0 556 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1710841341
transform 1 0 492 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1710841341
transform 1 0 484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1710841341
transform 1 0 380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1710841341
transform 1 0 340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1710841341
transform 1 0 2116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1710841341
transform 1 0 2068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1710841341
transform 1 0 2532 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1710841341
transform 1 0 2508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1710841341
transform 1 0 668 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1710841341
transform 1 0 628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1710841341
transform 1 0 212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1710841341
transform 1 0 84 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1710841341
transform 1 0 1244 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1710841341
transform 1 0 1228 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1710841341
transform 1 0 1876 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1710841341
transform 1 0 1780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1710841341
transform 1 0 1580 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1710841341
transform 1 0 1548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1710841341
transform 1 0 1548 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1710841341
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1710841341
transform 1 0 572 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1710841341
transform 1 0 1788 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1710841341
transform 1 0 1780 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1710841341
transform 1 0 1548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1710841341
transform 1 0 1244 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1710841341
transform 1 0 1204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1710841341
transform 1 0 1196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1710841341
transform 1 0 1092 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1710841341
transform 1 0 1076 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1710841341
transform 1 0 964 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1710841341
transform 1 0 956 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1710841341
transform 1 0 156 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1710841341
transform 1 0 92 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1710841341
transform 1 0 164 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1710841341
transform 1 0 84 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1710841341
transform 1 0 1300 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1710841341
transform 1 0 1076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1710841341
transform 1 0 964 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1710841341
transform 1 0 956 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1710841341
transform 1 0 2636 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1710841341
transform 1 0 2540 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1710841341
transform 1 0 1908 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1710841341
transform 1 0 1860 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1710841341
transform 1 0 2252 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1710841341
transform 1 0 2212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1710841341
transform 1 0 1652 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1710841341
transform 1 0 1636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1710841341
transform 1 0 1604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1710841341
transform 1 0 1588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1710841341
transform 1 0 1572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1710841341
transform 1 0 1444 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1710841341
transform 1 0 1396 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1710841341
transform 1 0 1380 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1710841341
transform 1 0 1340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1710841341
transform 1 0 1020 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1710841341
transform 1 0 948 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1710841341
transform 1 0 2364 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1710841341
transform 1 0 2284 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1710841341
transform 1 0 2452 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1710841341
transform 1 0 2340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1710841341
transform 1 0 2212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1710841341
transform 1 0 2116 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1710841341
transform 1 0 2556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1710841341
transform 1 0 2508 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1710841341
transform 1 0 1852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1710841341
transform 1 0 1828 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1710841341
transform 1 0 1828 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1710841341
transform 1 0 1780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1710841341
transform 1 0 1748 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1710841341
transform 1 0 1740 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1710841341
transform 1 0 1724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1710841341
transform 1 0 1708 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1710841341
transform 1 0 1708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1710841341
transform 1 0 1644 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1710841341
transform 1 0 1644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1710841341
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1710841341
transform 1 0 1596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1710841341
transform 1 0 1172 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1710841341
transform 1 0 564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1710841341
transform 1 0 508 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1710841341
transform 1 0 1932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1710841341
transform 1 0 1892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1710841341
transform 1 0 1452 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1710841341
transform 1 0 1444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1710841341
transform 1 0 1940 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1710841341
transform 1 0 1900 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1710841341
transform 1 0 676 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1710841341
transform 1 0 620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1710841341
transform 1 0 1844 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1710841341
transform 1 0 1748 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1710841341
transform 1 0 1780 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1710841341
transform 1 0 1732 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1710841341
transform 1 0 1500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1710841341
transform 1 0 1092 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1710841341
transform 1 0 1060 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1710841341
transform 1 0 1028 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1710841341
transform 1 0 956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1710841341
transform 1 0 1412 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1710841341
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1710841341
transform 1 0 1844 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1710841341
transform 1 0 1796 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1710841341
transform 1 0 1324 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1710841341
transform 1 0 1316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1710841341
transform 1 0 1844 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1710841341
transform 1 0 1804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1710841341
transform 1 0 1660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1710841341
transform 1 0 1140 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1710841341
transform 1 0 1140 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1710841341
transform 1 0 2284 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1710841341
transform 1 0 2284 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1710841341
transform 1 0 1892 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1710841341
transform 1 0 1852 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1710841341
transform 1 0 2460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1710841341
transform 1 0 2452 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1710841341
transform 1 0 2436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1710841341
transform 1 0 2244 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1710841341
transform 1 0 2052 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1710841341
transform 1 0 2028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1710841341
transform 1 0 1996 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1710841341
transform 1 0 1900 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1710841341
transform 1 0 2204 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1710841341
transform 1 0 2196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1710841341
transform 1 0 660 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1710841341
transform 1 0 628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1710841341
transform 1 0 508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1710841341
transform 1 0 444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1710841341
transform 1 0 396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1710841341
transform 1 0 996 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1710841341
transform 1 0 980 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1710841341
transform 1 0 2268 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1710841341
transform 1 0 2148 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1710841341
transform 1 0 2396 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1710841341
transform 1 0 2388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1710841341
transform 1 0 2364 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1710841341
transform 1 0 420 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1710841341
transform 1 0 356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1710841341
transform 1 0 1620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1710841341
transform 1 0 1612 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1710841341
transform 1 0 2316 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1710841341
transform 1 0 2268 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1710841341
transform 1 0 2332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1710841341
transform 1 0 2324 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1710841341
transform 1 0 500 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1710841341
transform 1 0 468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1710841341
transform 1 0 964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1710841341
transform 1 0 940 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1710841341
transform 1 0 2524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1710841341
transform 1 0 2516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1710841341
transform 1 0 2060 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1710841341
transform 1 0 1988 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1710841341
transform 1 0 1700 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1710841341
transform 1 0 1684 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1710841341
transform 1 0 1556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1710841341
transform 1 0 1500 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1710841341
transform 1 0 1324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1710841341
transform 1 0 1260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1710841341
transform 1 0 1196 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1710841341
transform 1 0 2332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1710841341
transform 1 0 2188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1710841341
transform 1 0 2068 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1710841341
transform 1 0 2004 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1710841341
transform 1 0 2636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1710841341
transform 1 0 2612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1710841341
transform 1 0 2652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1710841341
transform 1 0 2652 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1710841341
transform 1 0 660 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1710841341
transform 1 0 444 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1710841341
transform 1 0 1788 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1710841341
transform 1 0 1788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1710841341
transform 1 0 1500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1710841341
transform 1 0 1500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1710841341
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1710841341
transform 1 0 1892 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1710841341
transform 1 0 1324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1710841341
transform 1 0 1212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1710841341
transform 1 0 1044 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1710841341
transform 1 0 988 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1710841341
transform 1 0 388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1710841341
transform 1 0 356 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1710841341
transform 1 0 1204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1710841341
transform 1 0 1116 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1710841341
transform 1 0 484 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1710841341
transform 1 0 484 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1710841341
transform 1 0 908 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1710841341
transform 1 0 892 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1710841341
transform 1 0 268 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1710841341
transform 1 0 260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1710841341
transform 1 0 2236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1710841341
transform 1 0 2156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1710841341
transform 1 0 2036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1710841341
transform 1 0 2036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1710841341
transform 1 0 1908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1710841341
transform 1 0 1884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1710841341
transform 1 0 1476 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1710841341
transform 1 0 780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1710841341
transform 1 0 540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1710841341
transform 1 0 500 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1710841341
transform 1 0 460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1710841341
transform 1 0 412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1710841341
transform 1 0 2396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1710841341
transform 1 0 2396 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1710841341
transform 1 0 2316 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1710841341
transform 1 0 2284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1710841341
transform 1 0 2476 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1710841341
transform 1 0 2420 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1710841341
transform 1 0 2404 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1710841341
transform 1 0 2396 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1710841341
transform 1 0 2388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1710841341
transform 1 0 2364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1710841341
transform 1 0 2316 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1710841341
transform 1 0 2132 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1710841341
transform 1 0 2116 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1710841341
transform 1 0 1596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1710841341
transform 1 0 2116 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1710841341
transform 1 0 2028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1710841341
transform 1 0 1908 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1710841341
transform 1 0 1828 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1710841341
transform 1 0 1780 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1710841341
transform 1 0 2380 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1710841341
transform 1 0 2268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1710841341
transform 1 0 2196 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1710841341
transform 1 0 2148 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1710841341
transform 1 0 1940 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1710841341
transform 1 0 788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1710841341
transform 1 0 780 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1710841341
transform 1 0 1740 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1710841341
transform 1 0 1580 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1710841341
transform 1 0 1564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1710841341
transform 1 0 748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1710841341
transform 1 0 684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1710841341
transform 1 0 660 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1710841341
transform 1 0 2180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1710841341
transform 1 0 2012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1710841341
transform 1 0 1964 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1710841341
transform 1 0 1908 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1710841341
transform 1 0 1892 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1710841341
transform 1 0 2012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1710841341
transform 1 0 1924 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1710841341
transform 1 0 1876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1710841341
transform 1 0 1860 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1710841341
transform 1 0 1740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1710841341
transform 1 0 1628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1710841341
transform 1 0 1612 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1710841341
transform 1 0 1588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1710841341
transform 1 0 1556 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1710841341
transform 1 0 1516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1710841341
transform 1 0 2148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1710841341
transform 1 0 1476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1710841341
transform 1 0 1404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1710841341
transform 1 0 1388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1710841341
transform 1 0 1356 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1710841341
transform 1 0 772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1710841341
transform 1 0 612 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1710841341
transform 1 0 564 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1710841341
transform 1 0 532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1710841341
transform 1 0 404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1710841341
transform 1 0 2428 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1710841341
transform 1 0 2348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1710841341
transform 1 0 2340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1710841341
transform 1 0 2252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1710841341
transform 1 0 2036 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1710841341
transform 1 0 2020 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1710841341
transform 1 0 1980 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1710841341
transform 1 0 1908 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1710841341
transform 1 0 1844 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1710841341
transform 1 0 1764 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1710841341
transform 1 0 1588 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1710841341
transform 1 0 1476 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1710841341
transform 1 0 1476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1710841341
transform 1 0 2236 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1710841341
transform 1 0 2220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1710841341
transform 1 0 2212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1710841341
transform 1 0 2204 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1710841341
transform 1 0 1164 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1710841341
transform 1 0 1108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1710841341
transform 1 0 1108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1710841341
transform 1 0 2124 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1710841341
transform 1 0 2068 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1710841341
transform 1 0 2020 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1710841341
transform 1 0 1852 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1710841341
transform 1 0 1764 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1710841341
transform 1 0 1764 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1710841341
transform 1 0 1684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1710841341
transform 1 0 2436 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1710841341
transform 1 0 2292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1710841341
transform 1 0 1980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1710841341
transform 1 0 1972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1710841341
transform 1 0 1652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1710841341
transform 1 0 1580 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1710841341
transform 1 0 1508 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1710841341
transform 1 0 1508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1710841341
transform 1 0 1468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1710841341
transform 1 0 1524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1710841341
transform 1 0 1476 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1710841341
transform 1 0 1468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1710841341
transform 1 0 2540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1710841341
transform 1 0 2228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1710841341
transform 1 0 2140 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1710841341
transform 1 0 2132 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1710841341
transform 1 0 2604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1710841341
transform 1 0 2596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1710841341
transform 1 0 2540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1710841341
transform 1 0 2540 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1710841341
transform 1 0 1932 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1710841341
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1710841341
transform 1 0 1500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1710841341
transform 1 0 1428 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1710841341
transform 1 0 1164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1710841341
transform 1 0 1124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1710841341
transform 1 0 1124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1710841341
transform 1 0 1124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1710841341
transform 1 0 1740 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1710841341
transform 1 0 1684 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1710841341
transform 1 0 1468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1710841341
transform 1 0 1308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1710841341
transform 1 0 1124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1710841341
transform 1 0 1068 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1710841341
transform 1 0 332 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1710841341
transform 1 0 308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1710841341
transform 1 0 300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1710841341
transform 1 0 220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1710841341
transform 1 0 204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1710841341
transform 1 0 1228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1710841341
transform 1 0 644 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1710841341
transform 1 0 580 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1710841341
transform 1 0 492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1710841341
transform 1 0 492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1710841341
transform 1 0 460 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1710841341
transform 1 0 772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1710841341
transform 1 0 700 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1710841341
transform 1 0 1652 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1710841341
transform 1 0 1492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1710841341
transform 1 0 1484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1710841341
transform 1 0 1476 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1710841341
transform 1 0 1812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1710841341
transform 1 0 1772 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1710841341
transform 1 0 1276 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1710841341
transform 1 0 1212 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1710841341
transform 1 0 1084 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1710841341
transform 1 0 1036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1710841341
transform 1 0 2340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1710841341
transform 1 0 2244 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1710841341
transform 1 0 2084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1710841341
transform 1 0 2076 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1710841341
transform 1 0 2348 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1710841341
transform 1 0 2316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1710841341
transform 1 0 2252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1710841341
transform 1 0 2212 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1710841341
transform 1 0 2116 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1710841341
transform 1 0 2108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1710841341
transform 1 0 1980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1710841341
transform 1 0 1860 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1710841341
transform 1 0 2284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1710841341
transform 1 0 2172 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1710841341
transform 1 0 468 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1710841341
transform 1 0 436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1710841341
transform 1 0 2452 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1710841341
transform 1 0 2436 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1710841341
transform 1 0 468 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1710841341
transform 1 0 364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1710841341
transform 1 0 1412 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1710841341
transform 1 0 1412 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1710841341
transform 1 0 1372 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1710841341
transform 1 0 1340 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1710841341
transform 1 0 1292 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1710841341
transform 1 0 1284 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1710841341
transform 1 0 1132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1710841341
transform 1 0 196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1710841341
transform 1 0 132 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1710841341
transform 1 0 188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1710841341
transform 1 0 100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1710841341
transform 1 0 148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1710841341
transform 1 0 100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1710841341
transform 1 0 1172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1710841341
transform 1 0 1116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1710841341
transform 1 0 996 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1710841341
transform 1 0 324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1710841341
transform 1 0 252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1710841341
transform 1 0 204 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1710841341
transform 1 0 2332 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1710841341
transform 1 0 2316 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1710841341
transform 1 0 2292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1710841341
transform 1 0 2220 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1710841341
transform 1 0 2196 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1710841341
transform 1 0 2180 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1710841341
transform 1 0 1956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1710841341
transform 1 0 1676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1710841341
transform 1 0 2620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1710841341
transform 1 0 2532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1710841341
transform 1 0 2196 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1710841341
transform 1 0 2012 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1710841341
transform 1 0 1988 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1710841341
transform 1 0 1988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1710841341
transform 1 0 1708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1710841341
transform 1 0 1620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1710841341
transform 1 0 1612 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1710841341
transform 1 0 1596 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1710841341
transform 1 0 2236 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1710841341
transform 1 0 2140 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1710841341
transform 1 0 2108 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1710841341
transform 1 0 2084 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1710841341
transform 1 0 1988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1710841341
transform 1 0 1868 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1710841341
transform 1 0 1716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1710841341
transform 1 0 1436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1710841341
transform 1 0 1412 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1710841341
transform 1 0 228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1710841341
transform 1 0 228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1710841341
transform 1 0 148 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1710841341
transform 1 0 284 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1710841341
transform 1 0 172 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1710841341
transform 1 0 1612 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1710841341
transform 1 0 1596 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1710841341
transform 1 0 1476 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1710841341
transform 1 0 1372 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1710841341
transform 1 0 1916 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1710841341
transform 1 0 1876 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1710841341
transform 1 0 2268 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1710841341
transform 1 0 2220 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1710841341
transform 1 0 2292 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1710841341
transform 1 0 2260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1710841341
transform 1 0 1132 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1710841341
transform 1 0 940 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1710841341
transform 1 0 764 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1710841341
transform 1 0 556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1710841341
transform 1 0 396 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1710841341
transform 1 0 324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1710841341
transform 1 0 2532 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1710841341
transform 1 0 2316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1710841341
transform 1 0 2228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1710841341
transform 1 0 516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1710841341
transform 1 0 476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1710841341
transform 1 0 2356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1710841341
transform 1 0 2324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1710841341
transform 1 0 2284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1710841341
transform 1 0 2284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1710841341
transform 1 0 708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1710841341
transform 1 0 668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1710841341
transform 1 0 1644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1710841341
transform 1 0 1588 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1710841341
transform 1 0 1620 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1710841341
transform 1 0 1452 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1710841341
transform 1 0 1324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1710841341
transform 1 0 484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1710841341
transform 1 0 428 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1710841341
transform 1 0 428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1710841341
transform 1 0 396 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1710841341
transform 1 0 716 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1710841341
transform 1 0 644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1710841341
transform 1 0 596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1710841341
transform 1 0 556 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1710841341
transform 1 0 2516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1710841341
transform 1 0 2412 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1710841341
transform 1 0 2380 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1710841341
transform 1 0 2348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1710841341
transform 1 0 1940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1710841341
transform 1 0 2244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1710841341
transform 1 0 2148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1710841341
transform 1 0 2180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1710841341
transform 1 0 2132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1710841341
transform 1 0 2492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1710841341
transform 1 0 2404 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1710841341
transform 1 0 1244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1710841341
transform 1 0 1196 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1710841341
transform 1 0 1444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1710841341
transform 1 0 1420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1710841341
transform 1 0 2356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1710841341
transform 1 0 2260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1710841341
transform 1 0 2388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1710841341
transform 1 0 2348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1710841341
transform 1 0 1836 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1710841341
transform 1 0 1740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1710841341
transform 1 0 2252 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1710841341
transform 1 0 2228 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1710841341
transform 1 0 2220 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1710841341
transform 1 0 2220 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1710841341
transform 1 0 2204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1710841341
transform 1 0 2196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1710841341
transform 1 0 1756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1710841341
transform 1 0 884 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1710841341
transform 1 0 876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1710841341
transform 1 0 1820 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1710841341
transform 1 0 1788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1710841341
transform 1 0 2148 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1710841341
transform 1 0 2124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1710841341
transform 1 0 2092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1710841341
transform 1 0 2036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1710841341
transform 1 0 1820 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1710841341
transform 1 0 1772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1710841341
transform 1 0 1068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1710841341
transform 1 0 1012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1710841341
transform 1 0 2156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1710841341
transform 1 0 2132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1710841341
transform 1 0 2076 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1710841341
transform 1 0 1404 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1710841341
transform 1 0 1020 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1710841341
transform 1 0 2068 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1710841341
transform 1 0 2036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1710841341
transform 1 0 2220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1710841341
transform 1 0 2212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1710841341
transform 1 0 1988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1710841341
transform 1 0 1444 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1710841341
transform 1 0 860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1710841341
transform 1 0 860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1710841341
transform 1 0 844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1710841341
transform 1 0 844 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1710841341
transform 1 0 1684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1710841341
transform 1 0 1604 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1710841341
transform 1 0 2348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1710841341
transform 1 0 2236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1710841341
transform 1 0 2508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1710841341
transform 1 0 2460 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1710841341
transform 1 0 2444 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1710841341
transform 1 0 2404 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1710841341
transform 1 0 2268 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1710841341
transform 1 0 1692 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1710841341
transform 1 0 1420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1710841341
transform 1 0 1420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1710841341
transform 1 0 1332 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1710841341
transform 1 0 956 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1710841341
transform 1 0 852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1710841341
transform 1 0 628 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1710841341
transform 1 0 516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1710841341
transform 1 0 284 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1710841341
transform 1 0 172 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1710841341
transform 1 0 292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1710841341
transform 1 0 164 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1710841341
transform 1 0 1964 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1710841341
transform 1 0 1796 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1710841341
transform 1 0 1636 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1710841341
transform 1 0 1468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1710841341
transform 1 0 1460 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1710841341
transform 1 0 668 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1710841341
transform 1 0 548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1710841341
transform 1 0 484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1710841341
transform 1 0 2220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1710841341
transform 1 0 2212 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1710841341
transform 1 0 1452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1710841341
transform 1 0 1452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1710841341
transform 1 0 2484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1710841341
transform 1 0 2452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1710841341
transform 1 0 2180 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1710841341
transform 1 0 2020 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1710841341
transform 1 0 1828 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1710841341
transform 1 0 1796 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1710841341
transform 1 0 1780 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1710841341
transform 1 0 1780 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1710841341
transform 1 0 1620 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1710841341
transform 1 0 1580 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1710841341
transform 1 0 2484 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1710841341
transform 1 0 2476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1710841341
transform 1 0 1980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1710841341
transform 1 0 1908 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1710841341
transform 1 0 2276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1710841341
transform 1 0 2276 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1710841341
transform 1 0 2420 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1710841341
transform 1 0 2116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1710841341
transform 1 0 2388 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1710841341
transform 1 0 2364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1710841341
transform 1 0 2356 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1710841341
transform 1 0 2340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1710841341
transform 1 0 1436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1710841341
transform 1 0 1380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1710841341
transform 1 0 1212 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1710841341
transform 1 0 2028 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1710841341
transform 1 0 1988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1710841341
transform 1 0 2180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1710841341
transform 1 0 2100 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1710841341
transform 1 0 1212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1710841341
transform 1 0 1020 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1710841341
transform 1 0 132 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1710841341
transform 1 0 100 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1710841341
transform 1 0 116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1710841341
transform 1 0 108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1710841341
transform 1 0 228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1710841341
transform 1 0 116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1710841341
transform 1 0 292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1710841341
transform 1 0 268 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1710841341
transform 1 0 1052 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1710841341
transform 1 0 876 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1710841341
transform 1 0 628 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1710841341
transform 1 0 500 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1710841341
transform 1 0 484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1710841341
transform 1 0 380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1710841341
transform 1 0 268 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1710841341
transform 1 0 396 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1710841341
transform 1 0 380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1710841341
transform 1 0 324 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1710841341
transform 1 0 284 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1710841341
transform 1 0 140 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1710841341
transform 1 0 116 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1710841341
transform 1 0 452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1710841341
transform 1 0 116 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1710841341
transform 1 0 92 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1710841341
transform 1 0 92 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1710841341
transform 1 0 1956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1710841341
transform 1 0 1916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1710841341
transform 1 0 860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1710841341
transform 1 0 580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1710841341
transform 1 0 276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1710841341
transform 1 0 260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1710841341
transform 1 0 252 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1710841341
transform 1 0 252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1710841341
transform 1 0 564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1710841341
transform 1 0 348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1710841341
transform 1 0 332 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1710841341
transform 1 0 332 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1710841341
transform 1 0 284 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1710841341
transform 1 0 236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1710841341
transform 1 0 684 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1710841341
transform 1 0 604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1710841341
transform 1 0 316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1710841341
transform 1 0 140 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1710841341
transform 1 0 84 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1710841341
transform 1 0 228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1710841341
transform 1 0 116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1710841341
transform 1 0 308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1710841341
transform 1 0 244 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1710841341
transform 1 0 1156 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1710841341
transform 1 0 1156 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1710841341
transform 1 0 836 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1710841341
transform 1 0 364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1710841341
transform 1 0 348 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1710841341
transform 1 0 364 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1710841341
transform 1 0 300 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1710841341
transform 1 0 284 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1710841341
transform 1 0 284 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1710841341
transform 1 0 108 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1710841341
transform 1 0 108 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1710841341
transform 1 0 260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1710841341
transform 1 0 252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1710841341
transform 1 0 236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1710841341
transform 1 0 908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1710841341
transform 1 0 892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1710841341
transform 1 0 268 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1710841341
transform 1 0 204 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1710841341
transform 1 0 116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1710841341
transform 1 0 92 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1710841341
transform 1 0 212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1710841341
transform 1 0 100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1710841341
transform 1 0 276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1710841341
transform 1 0 228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1710841341
transform 1 0 212 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1710841341
transform 1 0 212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1710841341
transform 1 0 188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1710841341
transform 1 0 188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1710841341
transform 1 0 260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1710841341
transform 1 0 236 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1710841341
transform 1 0 340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1710841341
transform 1 0 268 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1710841341
transform 1 0 268 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1710841341
transform 1 0 244 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1710841341
transform 1 0 124 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1710841341
transform 1 0 108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1710841341
transform 1 0 268 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1710841341
transform 1 0 188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1710841341
transform 1 0 156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1710841341
transform 1 0 860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1710841341
transform 1 0 556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1710841341
transform 1 0 532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1710841341
transform 1 0 444 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1710841341
transform 1 0 428 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1710841341
transform 1 0 1356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1710841341
transform 1 0 1308 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1710841341
transform 1 0 1196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1710841341
transform 1 0 1092 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1710841341
transform 1 0 460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1710841341
transform 1 0 932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1710841341
transform 1 0 460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1710841341
transform 1 0 428 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1710841341
transform 1 0 388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1710841341
transform 1 0 276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1710841341
transform 1 0 180 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1710841341
transform 1 0 724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1710841341
transform 1 0 724 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1710841341
transform 1 0 620 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1710841341
transform 1 0 404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1710841341
transform 1 0 364 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1710841341
transform 1 0 436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1710841341
transform 1 0 356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1710841341
transform 1 0 364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1710841341
transform 1 0 364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1710841341
transform 1 0 540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1710841341
transform 1 0 348 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1710841341
transform 1 0 412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1710841341
transform 1 0 396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1710841341
transform 1 0 1364 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1710841341
transform 1 0 1332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1710841341
transform 1 0 1332 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1710841341
transform 1 0 1332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1710841341
transform 1 0 2140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1710841341
transform 1 0 1988 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1710841341
transform 1 0 1460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1710841341
transform 1 0 1460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1710841341
transform 1 0 1460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1710841341
transform 1 0 1060 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1710841341
transform 1 0 580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1710841341
transform 1 0 524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1710841341
transform 1 0 452 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1710841341
transform 1 0 444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1710841341
transform 1 0 724 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1710841341
transform 1 0 644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1710841341
transform 1 0 716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1710841341
transform 1 0 652 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1710841341
transform 1 0 884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1710841341
transform 1 0 692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1710841341
transform 1 0 644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1710841341
transform 1 0 612 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1710841341
transform 1 0 612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1710841341
transform 1 0 604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1710841341
transform 1 0 812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1710841341
transform 1 0 764 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1710841341
transform 1 0 868 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1710841341
transform 1 0 788 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1710841341
transform 1 0 620 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1710841341
transform 1 0 604 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1710841341
transform 1 0 596 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1710841341
transform 1 0 596 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1710841341
transform 1 0 516 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1710841341
transform 1 0 412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1710841341
transform 1 0 468 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1710841341
transform 1 0 420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1710841341
transform 1 0 428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1710841341
transform 1 0 420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1710841341
transform 1 0 628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1710841341
transform 1 0 452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1710841341
transform 1 0 468 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1710841341
transform 1 0 468 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1710841341
transform 1 0 1772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1710841341
transform 1 0 1724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1710841341
transform 1 0 892 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1710841341
transform 1 0 788 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1710841341
transform 1 0 788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1710841341
transform 1 0 604 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1710841341
transform 1 0 588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1710841341
transform 1 0 564 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1710841341
transform 1 0 660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1710841341
transform 1 0 564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1710841341
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1710841341
transform 1 0 492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1710841341
transform 1 0 492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1710841341
transform 1 0 500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1710841341
transform 1 0 500 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1710841341
transform 1 0 564 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1710841341
transform 1 0 516 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1710841341
transform 1 0 540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1710841341
transform 1 0 532 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1710841341
transform 1 0 660 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1710841341
transform 1 0 556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1710841341
transform 1 0 1220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1710841341
transform 1 0 1092 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1710841341
transform 1 0 668 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1710841341
transform 1 0 636 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1710841341
transform 1 0 620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1710841341
transform 1 0 612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1710841341
transform 1 0 596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1710841341
transform 1 0 1108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1710841341
transform 1 0 964 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1710841341
transform 1 0 604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1710841341
transform 1 0 604 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1710841341
transform 1 0 596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1710841341
transform 1 0 588 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1710841341
transform 1 0 540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1710841341
transform 1 0 564 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1710841341
transform 1 0 500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1710841341
transform 1 0 644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1710841341
transform 1 0 460 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1710841341
transform 1 0 484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1710841341
transform 1 0 428 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1710841341
transform 1 0 508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1710841341
transform 1 0 484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1710841341
transform 1 0 388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1710841341
transform 1 0 380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1710841341
transform 1 0 628 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1710841341
transform 1 0 396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1710841341
transform 1 0 588 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1710841341
transform 1 0 388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1710841341
transform 1 0 716 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1710841341
transform 1 0 716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1710841341
transform 1 0 660 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1710841341
transform 1 0 580 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1710841341
transform 1 0 1700 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1710841341
transform 1 0 1564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1710841341
transform 1 0 788 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1710841341
transform 1 0 692 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1710841341
transform 1 0 812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1710841341
transform 1 0 700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1710841341
transform 1 0 708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1710841341
transform 1 0 668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1710841341
transform 1 0 1804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1710841341
transform 1 0 1652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1710841341
transform 1 0 1108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1710841341
transform 1 0 1068 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1710841341
transform 1 0 692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1710841341
transform 1 0 820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1710841341
transform 1 0 748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1710841341
transform 1 0 756 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1710841341
transform 1 0 756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1710841341
transform 1 0 868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1710841341
transform 1 0 748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1710841341
transform 1 0 1068 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1710841341
transform 1 0 956 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1710841341
transform 1 0 916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1710841341
transform 1 0 916 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1710841341
transform 1 0 852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1710841341
transform 1 0 1004 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1710841341
transform 1 0 884 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1710841341
transform 1 0 884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1710841341
transform 1 0 724 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1710841341
transform 1 0 724 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1710841341
transform 1 0 868 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1710841341
transform 1 0 780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1710841341
transform 1 0 1284 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1710841341
transform 1 0 1172 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1710841341
transform 1 0 1124 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1710841341
transform 1 0 1068 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1710841341
transform 1 0 1012 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1710841341
transform 1 0 892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1710841341
transform 1 0 884 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1710841341
transform 1 0 844 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1710841341
transform 1 0 972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1710841341
transform 1 0 788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1710841341
transform 1 0 820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1710841341
transform 1 0 804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1710841341
transform 1 0 956 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1710841341
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1710841341
transform 1 0 916 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1710841341
transform 1 0 900 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1710841341
transform 1 0 1852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1710841341
transform 1 0 1780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1710841341
transform 1 0 1364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1710841341
transform 1 0 1316 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1710841341
transform 1 0 932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1710841341
transform 1 0 956 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1710841341
transform 1 0 932 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1710841341
transform 1 0 1852 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1710841341
transform 1 0 1844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1710841341
transform 1 0 1100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1710841341
transform 1 0 1044 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1710841341
transform 1 0 1908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1710841341
transform 1 0 1876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1710841341
transform 1 0 1156 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1710841341
transform 1 0 1132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1710841341
transform 1 0 1084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1710841341
transform 1 0 1084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1710841341
transform 1 0 1068 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1710841341
transform 1 0 924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1710841341
transform 1 0 908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1710841341
transform 1 0 828 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1710841341
transform 1 0 764 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1710841341
transform 1 0 740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1710841341
transform 1 0 684 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1710841341
transform 1 0 1244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1710841341
transform 1 0 1044 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1710841341
transform 1 0 980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1710841341
transform 1 0 980 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1710841341
transform 1 0 884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1710841341
transform 1 0 868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1710841341
transform 1 0 1148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1710841341
transform 1 0 1060 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1710841341
transform 1 0 828 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1710841341
transform 1 0 820 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1710841341
transform 1 0 804 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1710841341
transform 1 0 1044 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1710841341
transform 1 0 1028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1710841341
transform 1 0 844 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1710841341
transform 1 0 532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1710841341
transform 1 0 1036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1710841341
transform 1 0 1004 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1710841341
transform 1 0 1420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1710841341
transform 1 0 1404 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1710841341
transform 1 0 1380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1710841341
transform 1 0 1236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1710841341
transform 1 0 1204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1710841341
transform 1 0 1132 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1710841341
transform 1 0 1076 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1710841341
transform 1 0 820 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1710841341
transform 1 0 780 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1710841341
transform 1 0 1300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1710841341
transform 1 0 1276 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1710841341
transform 1 0 1292 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1710841341
transform 1 0 1220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1710841341
transform 1 0 1188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1710841341
transform 1 0 1084 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1710841341
transform 1 0 1764 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1710841341
transform 1 0 1732 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1710841341
transform 1 0 1204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1710841341
transform 1 0 1156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1710841341
transform 1 0 1196 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1710841341
transform 1 0 1140 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1710841341
transform 1 0 1228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1710841341
transform 1 0 1196 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1710841341
transform 1 0 1660 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1710841341
transform 1 0 1644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1710841341
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1710841341
transform 1 0 956 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1710841341
transform 1 0 1668 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1710841341
transform 1 0 1580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1710841341
transform 1 0 1204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1710841341
transform 1 0 1100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1710841341
transform 1 0 1052 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1710841341
transform 1 0 1164 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1710841341
transform 1 0 1132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1710841341
transform 1 0 1100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1710841341
transform 1 0 1020 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1710841341
transform 1 0 948 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1710841341
transform 1 0 940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1710841341
transform 1 0 292 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1710841341
transform 1 0 292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1710841341
transform 1 0 308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1710841341
transform 1 0 300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1710841341
transform 1 0 364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1710841341
transform 1 0 300 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1710841341
transform 1 0 540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1710841341
transform 1 0 324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1710841341
transform 1 0 604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1710841341
transform 1 0 524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1710841341
transform 1 0 492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1710841341
transform 1 0 452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1710841341
transform 1 0 404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1710841341
transform 1 0 620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1710841341
transform 1 0 452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1710841341
transform 1 0 452 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1710841341
transform 1 0 364 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1710841341
transform 1 0 364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1710841341
transform 1 0 356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1710841341
transform 1 0 284 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1710841341
transform 1 0 420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1710841341
transform 1 0 268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1710841341
transform 1 0 588 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1710841341
transform 1 0 484 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1710841341
transform 1 0 1364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1710841341
transform 1 0 1340 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1710841341
transform 1 0 1292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1710841341
transform 1 0 804 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1710841341
transform 1 0 572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1710841341
transform 1 0 444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1710841341
transform 1 0 580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1710841341
transform 1 0 580 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1710841341
transform 1 0 572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1710841341
transform 1 0 572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1710841341
transform 1 0 780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1710841341
transform 1 0 588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1710841341
transform 1 0 716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1710841341
transform 1 0 692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1710841341
transform 1 0 2004 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1710841341
transform 1 0 1948 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1710841341
transform 1 0 788 0 1 755
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1710841341
transform 1 0 780 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1710841341
transform 1 0 868 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1710841341
transform 1 0 524 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1710841341
transform 1 0 380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1710841341
transform 1 0 356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1710841341
transform 1 0 452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1710841341
transform 1 0 356 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1710841341
transform 1 0 620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1710841341
transform 1 0 500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1710841341
transform 1 0 740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1710841341
transform 1 0 684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1710841341
transform 1 0 668 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1710841341
transform 1 0 1260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1710841341
transform 1 0 996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1710841341
transform 1 0 700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1710841341
transform 1 0 700 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1710841341
transform 1 0 748 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1710841341
transform 1 0 516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1710841341
transform 1 0 828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1710841341
transform 1 0 716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1710841341
transform 1 0 692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1710841341
transform 1 0 596 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1710841341
transform 1 0 540 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1710841341
transform 1 0 540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1710841341
transform 1 0 756 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1710841341
transform 1 0 740 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1710841341
transform 1 0 1508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1710841341
transform 1 0 1348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1710841341
transform 1 0 796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1710841341
transform 1 0 780 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1710841341
transform 1 0 732 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1710841341
transform 1 0 620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1710841341
transform 1 0 596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1710841341
transform 1 0 668 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1710841341
transform 1 0 468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1710841341
transform 1 0 372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1710841341
transform 1 0 820 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1710841341
transform 1 0 812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1710841341
transform 1 0 1892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1710841341
transform 1 0 1492 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1710841341
transform 1 0 1484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1710841341
transform 1 0 1364 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1710841341
transform 1 0 1356 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1710841341
transform 1 0 956 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1710841341
transform 1 0 492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1710841341
transform 1 0 396 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1710841341
transform 1 0 412 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1710841341
transform 1 0 388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1710841341
transform 1 0 652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1710841341
transform 1 0 644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1710841341
transform 1 0 572 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1710841341
transform 1 0 556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1710841341
transform 1 0 540 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1710841341
transform 1 0 612 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1710841341
transform 1 0 596 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1710841341
transform 1 0 1044 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1710841341
transform 1 0 1028 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1710841341
transform 1 0 1100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1710841341
transform 1 0 1084 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1710841341
transform 1 0 1188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1710841341
transform 1 0 1124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1710841341
transform 1 0 1028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1710841341
transform 1 0 1012 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1710841341
transform 1 0 988 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1710841341
transform 1 0 972 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1710841341
transform 1 0 1388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1710841341
transform 1 0 1284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1710841341
transform 1 0 1060 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1710841341
transform 1 0 1052 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1710841341
transform 1 0 1004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1710841341
transform 1 0 924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1710841341
transform 1 0 852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1710841341
transform 1 0 852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1710841341
transform 1 0 964 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1710841341
transform 1 0 964 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1710841341
transform 1 0 1724 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1710841341
transform 1 0 1204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1710841341
transform 1 0 1084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1710841341
transform 1 0 1004 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1710841341
transform 1 0 940 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1710841341
transform 1 0 868 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1710841341
transform 1 0 868 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1710841341
transform 1 0 940 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1710841341
transform 1 0 924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1710841341
transform 1 0 892 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1710841341
transform 1 0 892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1710841341
transform 1 0 828 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1710841341
transform 1 0 796 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1710841341
transform 1 0 884 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1710841341
transform 1 0 868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1710841341
transform 1 0 972 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1710841341
transform 1 0 900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1710841341
transform 1 0 996 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1710841341
transform 1 0 940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1710841341
transform 1 0 1012 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1710841341
transform 1 0 1012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1710841341
transform 1 0 1052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1710841341
transform 1 0 1052 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1710841341
transform 1 0 924 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1710841341
transform 1 0 876 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1710841341
transform 1 0 836 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1710841341
transform 1 0 884 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1710841341
transform 1 0 884 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1710841341
transform 1 0 1196 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1710841341
transform 1 0 1164 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1710841341
transform 1 0 1180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1710841341
transform 1 0 1164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1710841341
transform 1 0 1220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1710841341
transform 1 0 1172 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1710841341
transform 1 0 1380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1710841341
transform 1 0 1188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1710841341
transform 1 0 1412 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1710841341
transform 1 0 1316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1710841341
transform 1 0 1300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1710841341
transform 1 0 1268 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1710841341
transform 1 0 1436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1710841341
transform 1 0 1436 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1710841341
transform 1 0 1412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1710841341
transform 1 0 1388 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1710841341
transform 1 0 1300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1710841341
transform 1 0 1276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1710841341
transform 1 0 1228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1710841341
transform 1 0 1196 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1710841341
transform 1 0 1332 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1710841341
transform 1 0 1332 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1710841341
transform 1 0 1596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1710841341
transform 1 0 1340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1710841341
transform 1 0 1268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1710841341
transform 1 0 1252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1710841341
transform 1 0 1244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1710841341
transform 1 0 1244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1710841341
transform 1 0 1396 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1710841341
transform 1 0 1396 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1710841341
transform 1 0 1356 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1710841341
transform 1 0 1348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1710841341
transform 1 0 1300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1710841341
transform 1 0 1260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1710841341
transform 1 0 1276 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1710841341
transform 1 0 1228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1710841341
transform 1 0 1268 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1710841341
transform 1 0 980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1710841341
transform 1 0 1324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1710841341
transform 1 0 1220 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1710841341
transform 1 0 1244 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1710841341
transform 1 0 1164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1710841341
transform 1 0 1340 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1710841341
transform 1 0 1308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1710841341
transform 1 0 1348 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1710841341
transform 1 0 1268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1710841341
transform 1 0 1260 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1710841341
transform 1 0 1268 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1710841341
transform 1 0 1268 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1710841341
transform 1 0 1564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1710841341
transform 1 0 1564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1710841341
transform 1 0 1508 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1710841341
transform 1 0 1484 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1710841341
transform 1 0 1436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1710841341
transform 1 0 1428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1710841341
transform 1 0 1492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1710841341
transform 1 0 1460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1710841341
transform 1 0 1420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1710841341
transform 1 0 1396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1710841341
transform 1 0 1388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1710841341
transform 1 0 1564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1710841341
transform 1 0 1524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1710841341
transform 1 0 1492 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1710841341
transform 1 0 1460 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1710841341
transform 1 0 1500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1710841341
transform 1 0 1468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1710841341
transform 1 0 2052 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1710841341
transform 1 0 1444 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1710841341
transform 1 0 972 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1710841341
transform 1 0 1388 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1710841341
transform 1 0 940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1710841341
transform 1 0 1508 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1710841341
transform 1 0 1436 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1710841341
transform 1 0 1484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1710841341
transform 1 0 1460 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1710841341
transform 1 0 1444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1710841341
transform 1 0 1404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1710841341
transform 1 0 1524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1710841341
transform 1 0 1476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1710841341
transform 1 0 1540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1710841341
transform 1 0 1508 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1710841341
transform 1 0 1556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1710841341
transform 1 0 1404 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1710841341
transform 1 0 1404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1710841341
transform 1 0 1588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1710841341
transform 1 0 1556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1710841341
transform 1 0 2100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1710841341
transform 1 0 2020 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1710841341
transform 1 0 2012 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1710841341
transform 1 0 1660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1710841341
transform 1 0 1628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1710841341
transform 1 0 1772 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1710841341
transform 1 0 1748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1710841341
transform 1 0 1724 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1710841341
transform 1 0 1724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1710841341
transform 1 0 1676 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1710841341
transform 1 0 1596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1710841341
transform 1 0 1692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1710841341
transform 1 0 1628 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1710841341
transform 1 0 1652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1710841341
transform 1 0 1644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1710841341
transform 1 0 1628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1710841341
transform 1 0 1628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1710841341
transform 1 0 1612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1710841341
transform 1 0 1588 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1710841341
transform 1 0 1556 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1710841341
transform 1 0 1716 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1710841341
transform 1 0 1692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1710841341
transform 1 0 1684 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1710841341
transform 1 0 1668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1710841341
transform 1 0 1596 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1710841341
transform 1 0 1572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1710841341
transform 1 0 1604 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1710841341
transform 1 0 1604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1710841341
transform 1 0 1780 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1710841341
transform 1 0 1764 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1710841341
transform 1 0 1812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1710841341
transform 1 0 1812 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1710841341
transform 1 0 2012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1710841341
transform 1 0 1764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1710841341
transform 1 0 1732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1710841341
transform 1 0 1748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1710841341
transform 1 0 1732 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1710841341
transform 1 0 1692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1710841341
transform 1 0 1692 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1710841341
transform 1 0 1660 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1710841341
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1710841341
transform 1 0 1596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1710841341
transform 1 0 1596 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1710841341
transform 1 0 1596 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1710841341
transform 1 0 1452 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1710841341
transform 1 0 1716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1710841341
transform 1 0 1660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1710841341
transform 1 0 1956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1710841341
transform 1 0 1908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1710841341
transform 1 0 1868 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1710841341
transform 1 0 1868 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1710841341
transform 1 0 1900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1710841341
transform 1 0 1820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1710841341
transform 1 0 1860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1710841341
transform 1 0 1780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1710841341
transform 1 0 1756 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1710841341
transform 1 0 1756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1710841341
transform 1 0 1700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1710841341
transform 1 0 1844 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1710841341
transform 1 0 1812 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1710841341
transform 1 0 1748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1710841341
transform 1 0 1740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1710841341
transform 1 0 1908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1710841341
transform 1 0 1876 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1710841341
transform 1 0 1956 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1710841341
transform 1 0 1916 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1710841341
transform 1 0 1940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1710841341
transform 1 0 1916 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1710841341
transform 1 0 1836 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1710841341
transform 1 0 1820 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1710841341
transform 1 0 1804 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1710841341
transform 1 0 1772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1710841341
transform 1 0 1884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1710841341
transform 1 0 1828 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1710841341
transform 1 0 1788 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1710841341
transform 1 0 1516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1710841341
transform 1 0 1844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1710841341
transform 1 0 1804 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1710841341
transform 1 0 1732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1710841341
transform 1 0 1668 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1710841341
transform 1 0 1668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1710841341
transform 1 0 1636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1710841341
transform 1 0 2140 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1710841341
transform 1 0 1756 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1710841341
transform 1 0 1708 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1710841341
transform 1 0 1708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1710841341
transform 1 0 1500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1710841341
transform 1 0 1476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1710841341
transform 1 0 1908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1710841341
transform 1 0 1820 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1710841341
transform 1 0 1844 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1710841341
transform 1 0 1804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1710841341
transform 1 0 1980 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1710841341
transform 1 0 1756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1710841341
transform 1 0 1684 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1710841341
transform 1 0 1756 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1710841341
transform 1 0 1756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1710841341
transform 1 0 1764 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1710841341
transform 1 0 1764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1710841341
transform 1 0 1596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1710841341
transform 1 0 1524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1710841341
transform 1 0 2596 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1710841341
transform 1 0 2580 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1710841341
transform 1 0 2412 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1710841341
transform 1 0 2020 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1710841341
transform 1 0 1948 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1710841341
transform 1 0 1540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1710841341
transform 1 0 2412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1710841341
transform 1 0 2404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1710841341
transform 1 0 2372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1710841341
transform 1 0 2372 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1710841341
transform 1 0 2260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1710841341
transform 1 0 2228 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1710841341
transform 1 0 2252 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1710841341
transform 1 0 2236 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1710841341
transform 1 0 2140 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1710841341
transform 1 0 2116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1710841341
transform 1 0 2348 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1710841341
transform 1 0 2212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1710841341
transform 1 0 2428 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1710841341
transform 1 0 2084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1710841341
transform 1 0 2444 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1710841341
transform 1 0 2388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1710841341
transform 1 0 2276 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1710841341
transform 1 0 2236 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1710841341
transform 1 0 2340 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1710841341
transform 1 0 2340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1710841341
transform 1 0 2204 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1710841341
transform 1 0 1996 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1710841341
transform 1 0 1708 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1710841341
transform 1 0 2172 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1710841341
transform 1 0 2036 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1710841341
transform 1 0 2092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1710841341
transform 1 0 1972 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1710841341
transform 1 0 2084 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1710841341
transform 1 0 2044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1710841341
transform 1 0 1980 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1710841341
transform 1 0 1588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1710841341
transform 1 0 2148 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1710841341
transform 1 0 2060 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1710841341
transform 1 0 2644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1710841341
transform 1 0 2636 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1710841341
transform 1 0 2380 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1710841341
transform 1 0 2356 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1710841341
transform 1 0 1948 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1710841341
transform 1 0 1716 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1710841341
transform 1 0 1556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1710841341
transform 1 0 2444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1710841341
transform 1 0 2444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1710841341
transform 1 0 2412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1710841341
transform 1 0 2332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1710841341
transform 1 0 2276 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1710841341
transform 1 0 2244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1710841341
transform 1 0 2228 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1710841341
transform 1 0 2244 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1710841341
transform 1 0 2220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1710841341
transform 1 0 2212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1710841341
transform 1 0 2012 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1710841341
transform 1 0 2372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1710841341
transform 1 0 2324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1710841341
transform 1 0 2220 0 1 385
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1710841341
transform 1 0 2220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1710841341
transform 1 0 2196 0 1 385
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1710841341
transform 1 0 2188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1710841341
transform 1 0 2236 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1710841341
transform 1 0 2228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1710841341
transform 1 0 2140 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1710841341
transform 1 0 2108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1710841341
transform 1 0 2372 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1710841341
transform 1 0 2284 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1710841341
transform 1 0 2372 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1710841341
transform 1 0 2348 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1710841341
transform 1 0 2284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1710841341
transform 1 0 2124 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1710841341
transform 1 0 2116 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1710841341
transform 1 0 1900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1710841341
transform 1 0 1836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1710841341
transform 1 0 2532 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1710841341
transform 1 0 2316 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1710841341
transform 1 0 2036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1710841341
transform 1 0 2004 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1710841341
transform 1 0 2380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1710841341
transform 1 0 2364 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1710841341
transform 1 0 2172 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1710841341
transform 1 0 2092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1710841341
transform 1 0 2396 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1710841341
transform 1 0 2348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1710841341
transform 1 0 2436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1710841341
transform 1 0 2372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1710841341
transform 1 0 2300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1710841341
transform 1 0 2276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1710841341
transform 1 0 2268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1710841341
transform 1 0 2236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1710841341
transform 1 0 2252 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1710841341
transform 1 0 2220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1710841341
transform 1 0 2252 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1710841341
transform 1 0 2236 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1710841341
transform 1 0 2188 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1710841341
transform 1 0 2156 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1710841341
transform 1 0 2500 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1710841341
transform 1 0 2476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1710841341
transform 1 0 2452 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1710841341
transform 1 0 2180 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1710841341
transform 1 0 2156 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1710841341
transform 1 0 2116 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1710841341
transform 1 0 2132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1710841341
transform 1 0 2060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1710841341
transform 1 0 2404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1710841341
transform 1 0 2180 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1710841341
transform 1 0 2172 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1710841341
transform 1 0 2156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1710841341
transform 1 0 2540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1710841341
transform 1 0 2500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1710841341
transform 1 0 2188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1710841341
transform 1 0 1956 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1710841341
transform 1 0 2340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1710841341
transform 1 0 2188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1710841341
transform 1 0 2628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1710841341
transform 1 0 2628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1710841341
transform 1 0 2580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1710841341
transform 1 0 2484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1710841341
transform 1 0 2380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1710841341
transform 1 0 2468 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1710841341
transform 1 0 2436 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1710841341
transform 1 0 2556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1710841341
transform 1 0 2556 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1710841341
transform 1 0 2516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1710841341
transform 1 0 2444 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1710841341
transform 1 0 2156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1710841341
transform 1 0 1964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1710841341
transform 1 0 1900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1710841341
transform 1 0 2460 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1710841341
transform 1 0 2460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1710841341
transform 1 0 2556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1710841341
transform 1 0 2476 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1710841341
transform 1 0 2460 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1710841341
transform 1 0 2452 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1710841341
transform 1 0 2172 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1710841341
transform 1 0 2084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1710841341
transform 1 0 2548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1710841341
transform 1 0 2532 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1710841341
transform 1 0 2604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1710841341
transform 1 0 2588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1710841341
transform 1 0 2660 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1710841341
transform 1 0 2548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1710841341
transform 1 0 2660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1710841341
transform 1 0 2628 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1710841341
transform 1 0 2604 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1710841341
transform 1 0 2660 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1710841341
transform 1 0 2620 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1710841341
transform 1 0 2636 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1710841341
transform 1 0 2580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1710841341
transform 1 0 2596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1710841341
transform 1 0 2556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1710841341
transform 1 0 2540 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1710841341
transform 1 0 2420 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1710841341
transform 1 0 2508 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1710841341
transform 1 0 2204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1710841341
transform 1 0 2508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1710841341
transform 1 0 2388 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1710841341
transform 1 0 2260 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1710841341
transform 1 0 1828 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1710841341
transform 1 0 2612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1710841341
transform 1 0 2484 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1710841341
transform 1 0 2468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1710841341
transform 1 0 2564 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1710841341
transform 1 0 2124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1710841341
transform 1 0 2612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1710841341
transform 1 0 2596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1710841341
transform 1 0 2580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1710841341
transform 1 0 2564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1710841341
transform 1 0 2564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1710841341
transform 1 0 2524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1710841341
transform 1 0 2660 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1710841341
transform 1 0 2628 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1710841341
transform 1 0 2636 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1710841341
transform 1 0 2620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1710841341
transform 1 0 2564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1710841341
transform 1 0 2532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1710841341
transform 1 0 2092 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1710841341
transform 1 0 1892 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1710841341
transform 1 0 1652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1710841341
transform 1 0 2620 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1710841341
transform 1 0 2620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1710841341
transform 1 0 2628 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1710841341
transform 1 0 2604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1710841341
transform 1 0 2604 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1710841341
transform 1 0 2556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1710841341
transform 1 0 2116 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1710841341
transform 1 0 2044 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1710841341
transform 1 0 2644 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1710841341
transform 1 0 2532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1710841341
transform 1 0 2660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1710841341
transform 1 0 2636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1710841341
transform 1 0 2604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1710841341
transform 1 0 2580 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1710841341
transform 1 0 2596 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1710841341
transform 1 0 2524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1710841341
transform 1 0 2540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1710841341
transform 1 0 2460 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1710841341
transform 1 0 2460 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1710841341
transform 1 0 2580 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1710841341
transform 1 0 2556 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1710841341
transform 1 0 2540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1710841341
transform 1 0 2244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1710841341
transform 1 0 2532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1710841341
transform 1 0 2468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1710841341
transform 1 0 2396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1710841341
transform 1 0 2396 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1710841341
transform 1 0 2372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1710841341
transform 1 0 2300 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1710841341
transform 1 0 2148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1710841341
transform 1 0 2428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1710841341
transform 1 0 2404 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1710841341
transform 1 0 2372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1710841341
transform 1 0 1900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1710841341
transform 1 0 2532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1710841341
transform 1 0 2276 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1710841341
transform 1 0 2068 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1710841341
transform 1 0 2020 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1710841341
transform 1 0 2052 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1710841341
transform 1 0 2036 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1710841341
transform 1 0 2068 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1710841341
transform 1 0 2052 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1710841341
transform 1 0 2196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1710841341
transform 1 0 2180 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1710841341
transform 1 0 2204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1710841341
transform 1 0 2164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1710841341
transform 1 0 2316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1710841341
transform 1 0 2284 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1710841341
transform 1 0 2388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1710841341
transform 1 0 2340 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1710841341
transform 1 0 2124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1710841341
transform 1 0 2124 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1710841341
transform 1 0 2108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1710841341
transform 1 0 2092 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1710841341
transform 1 0 2060 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1710841341
transform 1 0 2236 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1710841341
transform 1 0 2076 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1710841341
transform 1 0 2076 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1710841341
transform 1 0 2060 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1710841341
transform 1 0 1748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1710841341
transform 1 0 2532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1710841341
transform 1 0 2452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1710841341
transform 1 0 2436 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1710841341
transform 1 0 2188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1710841341
transform 1 0 2468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1710841341
transform 1 0 2396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1710841341
transform 1 0 2348 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1710841341
transform 1 0 2348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1710841341
transform 1 0 2324 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1710841341
transform 1 0 2236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1710841341
transform 1 0 1772 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1710841341
transform 1 0 2388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1710841341
transform 1 0 2356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1710841341
transform 1 0 1956 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1710841341
transform 1 0 1716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1710841341
transform 1 0 2220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1710841341
transform 1 0 2188 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1710841341
transform 1 0 2260 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1710841341
transform 1 0 2204 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1710841341
transform 1 0 2484 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1710841341
transform 1 0 2300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1710841341
transform 1 0 2468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1710841341
transform 1 0 2044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1710841341
transform 1 0 1940 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1710841341
transform 1 0 1892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1710841341
transform 1 0 1924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1710841341
transform 1 0 1900 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1710841341
transform 1 0 796 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1710841341
transform 1 0 772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1710841341
transform 1 0 772 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1710841341
transform 1 0 2340 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1710841341
transform 1 0 2300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1710841341
transform 1 0 1732 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1710841341
transform 1 0 1732 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1710841341
transform 1 0 844 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1710841341
transform 1 0 788 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1710841341
transform 1 0 804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1710841341
transform 1 0 804 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1710841341
transform 1 0 724 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1710841341
transform 1 0 724 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1710841341
transform 1 0 1036 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1710841341
transform 1 0 988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1710841341
transform 1 0 740 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1710841341
transform 1 0 708 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1710841341
transform 1 0 620 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1710841341
transform 1 0 1916 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1710841341
transform 1 0 1748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1710841341
transform 1 0 1540 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1710841341
transform 1 0 1412 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1710841341
transform 1 0 1412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1710841341
transform 1 0 1988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1710841341
transform 1 0 1844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1710841341
transform 1 0 2644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1710841341
transform 1 0 2524 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1710841341
transform 1 0 2484 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1710841341
transform 1 0 2372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1710841341
transform 1 0 2508 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1710841341
transform 1 0 2444 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1710841341
transform 1 0 2380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1710841341
transform 1 0 2228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1710841341
transform 1 0 2164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1710841341
transform 1 0 2068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1710841341
transform 1 0 1900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1710841341
transform 1 0 2100 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1710841341
transform 1 0 2052 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1710841341
transform 1 0 1972 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1710841341
transform 1 0 1804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1710841341
transform 1 0 2372 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1710841341
transform 1 0 2348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1710841341
transform 1 0 2580 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1710841341
transform 1 0 2500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1710841341
transform 1 0 2548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1710841341
transform 1 0 2052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1710841341
transform 1 0 1964 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1710841341
transform 1 0 1892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1710841341
transform 1 0 1932 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1710841341
transform 1 0 1900 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1710841341
transform 1 0 1100 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1710841341
transform 1 0 1060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1710841341
transform 1 0 884 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1710841341
transform 1 0 1116 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1710841341
transform 1 0 1068 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1710841341
transform 1 0 964 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1710841341
transform 1 0 844 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1710841341
transform 1 0 740 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1710841341
transform 1 0 1052 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1710841341
transform 1 0 1052 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1710841341
transform 1 0 2124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1710841341
transform 1 0 1972 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1710841341
transform 1 0 1940 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1710841341
transform 1 0 1892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1710841341
transform 1 0 2148 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1710841341
transform 1 0 1964 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1710841341
transform 1 0 2004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1710841341
transform 1 0 1980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1710841341
transform 1 0 2060 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1710841341
transform 1 0 2044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1710841341
transform 1 0 1988 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1710841341
transform 1 0 1868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1710841341
transform 1 0 1740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1710841341
transform 1 0 2284 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1710841341
transform 1 0 1996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1710841341
transform 1 0 1748 0 1 1695
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1710841341
transform 1 0 1748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1710841341
transform 1 0 2148 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1710841341
transform 1 0 2148 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1710841341
transform 1 0 1820 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1710841341
transform 1 0 1796 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1710841341
transform 1 0 1852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1710841341
transform 1 0 1804 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1710841341
transform 1 0 1932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1710841341
transform 1 0 1892 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1710841341
transform 1 0 1764 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1710841341
transform 1 0 1748 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1710841341
transform 1 0 1804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1710841341
transform 1 0 1796 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1710841341
transform 1 0 1820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1710841341
transform 1 0 1788 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1710841341
transform 1 0 1868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1710841341
transform 1 0 1852 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1710841341
transform 1 0 956 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1710841341
transform 1 0 916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1710841341
transform 1 0 732 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1710841341
transform 1 0 1164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1710841341
transform 1 0 852 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1710841341
transform 1 0 836 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1710841341
transform 1 0 684 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1710841341
transform 1 0 676 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1710841341
transform 1 0 932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1710841341
transform 1 0 924 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1710841341
transform 1 0 2140 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1710841341
transform 1 0 1940 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1710841341
transform 1 0 1908 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1710841341
transform 1 0 1668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1710841341
transform 1 0 1580 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1710841341
transform 1 0 1580 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1710841341
transform 1 0 2644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1710841341
transform 1 0 2492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1710841341
transform 1 0 2460 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1710841341
transform 1 0 2436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1710841341
transform 1 0 2476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1710841341
transform 1 0 2340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1710841341
transform 1 0 2476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1710841341
transform 1 0 2436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1710841341
transform 1 0 2332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1710841341
transform 1 0 2276 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1710841341
transform 1 0 2212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1710841341
transform 1 0 2412 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1710841341
transform 1 0 2404 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1710841341
transform 1 0 2580 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1710841341
transform 1 0 2524 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1710841341
transform 1 0 2556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1710841341
transform 1 0 2244 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1710841341
transform 1 0 2540 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1710841341
transform 1 0 2244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1710841341
transform 1 0 1716 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1710841341
transform 1 0 1604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1710841341
transform 1 0 1396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1710841341
transform 1 0 1268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1710841341
transform 1 0 2252 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1710841341
transform 1 0 2228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1710841341
transform 1 0 2172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1710841341
transform 1 0 1916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1710841341
transform 1 0 2156 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1710841341
transform 1 0 1932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1710841341
transform 1 0 1900 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1710841341
transform 1 0 1876 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1710841341
transform 1 0 804 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1710841341
transform 1 0 756 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1710841341
transform 1 0 884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1710841341
transform 1 0 820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1710841341
transform 1 0 700 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1710841341
transform 1 0 2188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1710841341
transform 1 0 1988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1710841341
transform 1 0 2636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1710841341
transform 1 0 2636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1710841341
transform 1 0 2612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1710841341
transform 1 0 2540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1710841341
transform 1 0 2508 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1710841341
transform 1 0 2364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1710841341
transform 1 0 2540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1710841341
transform 1 0 2468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1710841341
transform 1 0 2508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1710841341
transform 1 0 2436 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1710841341
transform 1 0 2436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1710841341
transform 1 0 2420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1710841341
transform 1 0 2452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1710841341
transform 1 0 2444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1710841341
transform 1 0 2244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1710841341
transform 1 0 2116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1710841341
transform 1 0 2412 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1710841341
transform 1 0 2404 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1710841341
transform 1 0 2364 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1710841341
transform 1 0 2356 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1710841341
transform 1 0 2444 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1710841341
transform 1 0 2188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1710841341
transform 1 0 2548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1710841341
transform 1 0 2532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1710841341
transform 1 0 2492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1710841341
transform 1 0 2484 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1710841341
transform 1 0 2532 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1710841341
transform 1 0 2516 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1710841341
transform 1 0 2508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1710841341
transform 1 0 2484 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1710841341
transform 1 0 2308 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1710841341
transform 1 0 2132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1710841341
transform 1 0 1956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1710841341
transform 1 0 2532 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1710841341
transform 1 0 2516 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1710841341
transform 1 0 2172 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1710841341
transform 1 0 2092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1710841341
transform 1 0 2620 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1710841341
transform 1 0 2620 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1710841341
transform 1 0 2652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1710841341
transform 1 0 2580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1710841341
transform 1 0 2532 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1710841341
transform 1 0 2460 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1710841341
transform 1 0 2580 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1710841341
transform 1 0 2548 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1710841341
transform 1 0 2524 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1710841341
transform 1 0 2628 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1710841341
transform 1 0 2596 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1710841341
transform 1 0 2348 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1710841341
transform 1 0 2332 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1710841341
transform 1 0 2372 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1710841341
transform 1 0 2372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1710841341
transform 1 0 2316 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1710841341
transform 1 0 2292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1710841341
transform 1 0 2348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1710841341
transform 1 0 2260 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1710841341
transform 1 0 2244 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1710841341
transform 1 0 2228 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1710841341
transform 1 0 2228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1710841341
transform 1 0 2268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1710841341
transform 1 0 2172 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1710841341
transform 1 0 2060 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1710841341
transform 1 0 2060 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1710841341
transform 1 0 2260 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1710841341
transform 1 0 2260 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1710841341
transform 1 0 2204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1710841341
transform 1 0 2180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1710841341
transform 1 0 2180 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1710841341
transform 1 0 2196 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1710841341
transform 1 0 2188 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1710841341
transform 1 0 2340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1710841341
transform 1 0 2180 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1710841341
transform 1 0 2436 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1710841341
transform 1 0 2340 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1710841341
transform 1 0 2324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1710841341
transform 1 0 2324 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1710841341
transform 1 0 2124 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1710841341
transform 1 0 1692 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1710841341
transform 1 0 1684 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1710841341
transform 1 0 1684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1710841341
transform 1 0 2308 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1710841341
transform 1 0 2236 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1710841341
transform 1 0 2356 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1710841341
transform 1 0 2356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1710841341
transform 1 0 2284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1710841341
transform 1 0 2244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1710841341
transform 1 0 2180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1710841341
transform 1 0 2156 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1710841341
transform 1 0 2204 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1710841341
transform 1 0 2164 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1710841341
transform 1 0 2276 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1710841341
transform 1 0 2268 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1710841341
transform 1 0 2180 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1710841341
transform 1 0 2276 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1710841341
transform 1 0 2268 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1710841341
transform 1 0 2028 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1710841341
transform 1 0 2020 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1710841341
transform 1 0 2100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1710841341
transform 1 0 2004 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1710841341
transform 1 0 2020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1710841341
transform 1 0 1964 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1710841341
transform 1 0 2020 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1710841341
transform 1 0 1972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1710841341
transform 1 0 1876 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1710841341
transform 1 0 1860 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1710841341
transform 1 0 1892 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1710841341
transform 1 0 1836 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1710841341
transform 1 0 1836 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1710841341
transform 1 0 1820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1710841341
transform 1 0 2076 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1710841341
transform 1 0 1932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1710841341
transform 1 0 1956 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1710841341
transform 1 0 1956 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1710841341
transform 1 0 1900 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1710841341
transform 1 0 1900 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1710841341
transform 1 0 1860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1710841341
transform 1 0 1956 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1710841341
transform 1 0 1916 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1710841341
transform 1 0 2036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1710841341
transform 1 0 1972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1710841341
transform 1 0 1844 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1710841341
transform 1 0 1820 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1710841341
transform 1 0 1780 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1710841341
transform 1 0 1564 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1710841341
transform 1 0 1260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1710841341
transform 1 0 940 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1710841341
transform 1 0 940 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1710841341
transform 1 0 908 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1710841341
transform 1 0 1876 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1710841341
transform 1 0 1852 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1710841341
transform 1 0 1700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1710841341
transform 1 0 1564 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1710841341
transform 1 0 1564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1710841341
transform 1 0 2036 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1710841341
transform 1 0 1884 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1710841341
transform 1 0 2108 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1710841341
transform 1 0 2036 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1710841341
transform 1 0 2012 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1710841341
transform 1 0 2012 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1710841341
transform 1 0 2068 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1710841341
transform 1 0 2044 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1710841341
transform 1 0 1948 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1710841341
transform 1 0 1892 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1710841341
transform 1 0 2028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1710841341
transform 1 0 2004 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1710841341
transform 1 0 1884 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1710841341
transform 1 0 1828 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1710841341
transform 1 0 1972 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1710841341
transform 1 0 1932 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1710841341
transform 1 0 1828 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1710841341
transform 1 0 1988 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1710841341
transform 1 0 1988 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1710841341
transform 1 0 1724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1710841341
transform 1 0 1724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1710841341
transform 1 0 1756 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1710841341
transform 1 0 1740 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1710841341
transform 1 0 1804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1710841341
transform 1 0 1764 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1710841341
transform 1 0 1780 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1710841341
transform 1 0 1772 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1710841341
transform 1 0 932 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1710841341
transform 1 0 868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1710841341
transform 1 0 868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1710841341
transform 1 0 1708 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1710841341
transform 1 0 1700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1710841341
transform 1 0 1684 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1710841341
transform 1 0 1588 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1710841341
transform 1 0 1540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1710841341
transform 1 0 1116 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1710841341
transform 1 0 932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1710841341
transform 1 0 844 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1710841341
transform 1 0 804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1710841341
transform 1 0 1788 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1710841341
transform 1 0 1684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1710841341
transform 1 0 1596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1710841341
transform 1 0 1524 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1710841341
transform 1 0 1484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1710841341
transform 1 0 1428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1710841341
transform 1 0 1396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1710841341
transform 1 0 1388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1710841341
transform 1 0 1196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1710841341
transform 1 0 836 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1710841341
transform 1 0 1668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1710841341
transform 1 0 1596 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1710841341
transform 1 0 1484 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1710841341
transform 1 0 1380 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1710841341
transform 1 0 1348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1710841341
transform 1 0 972 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1710841341
transform 1 0 1732 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1710841341
transform 1 0 1732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1710841341
transform 1 0 1748 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1710841341
transform 1 0 1668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1710841341
transform 1 0 1620 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1710841341
transform 1 0 1612 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1710841341
transform 1 0 1612 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1710841341
transform 1 0 1596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1710841341
transform 1 0 1540 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1710841341
transform 1 0 1532 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1710841341
transform 1 0 1508 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1710841341
transform 1 0 1356 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1710841341
transform 1 0 796 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1710841341
transform 1 0 780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1710841341
transform 1 0 780 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1710841341
transform 1 0 772 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1710841341
transform 1 0 1580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1710841341
transform 1 0 1516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1710841341
transform 1 0 1500 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1710841341
transform 1 0 1052 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1710841341
transform 1 0 1124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1710841341
transform 1 0 1084 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1710841341
transform 1 0 1004 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1710841341
transform 1 0 980 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1710841341
transform 1 0 964 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1710841341
transform 1 0 1556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1710841341
transform 1 0 1556 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1710841341
transform 1 0 1596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1710841341
transform 1 0 1572 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1710841341
transform 1 0 1516 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1710841341
transform 1 0 1492 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1710841341
transform 1 0 1356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1710841341
transform 1 0 1332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1710841341
transform 1 0 1292 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1710841341
transform 1 0 1268 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1710841341
transform 1 0 1356 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1710841341
transform 1 0 1276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1710841341
transform 1 0 1364 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1710841341
transform 1 0 1364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1710841341
transform 1 0 1332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1710841341
transform 1 0 1316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1710841341
transform 1 0 1444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1710841341
transform 1 0 1324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1710841341
transform 1 0 1404 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1710841341
transform 1 0 1396 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1710841341
transform 1 0 1388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1710841341
transform 1 0 772 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1710841341
transform 1 0 1572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1710841341
transform 1 0 1484 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1710841341
transform 1 0 1284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1710841341
transform 1 0 1276 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1710841341
transform 1 0 1276 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1710841341
transform 1 0 1268 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1710841341
transform 1 0 1340 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1710841341
transform 1 0 1252 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1710841341
transform 1 0 1356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1710841341
transform 1 0 1236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1710841341
transform 1 0 1388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1710841341
transform 1 0 1268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1710841341
transform 1 0 1236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1710841341
transform 1 0 1268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1710841341
transform 1 0 1204 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1710841341
transform 1 0 1132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1710841341
transform 1 0 1132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1710841341
transform 1 0 1396 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1710841341
transform 1 0 1332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1710841341
transform 1 0 1348 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1710841341
transform 1 0 1028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1710841341
transform 1 0 1476 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1710841341
transform 1 0 1412 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1710841341
transform 1 0 1492 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1710841341
transform 1 0 1436 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1710841341
transform 1 0 1228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1710841341
transform 1 0 1092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1710841341
transform 1 0 1236 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1710841341
transform 1 0 1132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1710841341
transform 1 0 1004 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1710841341
transform 1 0 1004 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1710841341
transform 1 0 1316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1710841341
transform 1 0 1300 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1710841341
transform 1 0 1372 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1710841341
transform 1 0 1300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1710841341
transform 1 0 1332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1710841341
transform 1 0 1284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1710841341
transform 1 0 1212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1710841341
transform 1 0 1052 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1710841341
transform 1 0 1412 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1710841341
transform 1 0 1340 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1710841341
transform 1 0 1316 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1710841341
transform 1 0 1140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1710841341
transform 1 0 1164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1710841341
transform 1 0 1132 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1710841341
transform 1 0 1124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1710841341
transform 1 0 1100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1710841341
transform 1 0 1068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1710841341
transform 1 0 1044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1710841341
transform 1 0 852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1710841341
transform 1 0 772 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1710841341
transform 1 0 724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1710841341
transform 1 0 1428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1710841341
transform 1 0 1404 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1710841341
transform 1 0 1196 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1710841341
transform 1 0 1188 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1710841341
transform 1 0 1164 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1710841341
transform 1 0 1148 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1710841341
transform 1 0 1236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1710841341
transform 1 0 1156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1710841341
transform 1 0 1284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1710841341
transform 1 0 1252 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1710841341
transform 1 0 1236 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1710841341
transform 1 0 1228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1710841341
transform 1 0 1404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1710841341
transform 1 0 1268 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1710841341
transform 1 0 1508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1710841341
transform 1 0 1404 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1710841341
transform 1 0 1572 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1710841341
transform 1 0 1540 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1710841341
transform 1 0 1508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1710841341
transform 1 0 1044 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1710841341
transform 1 0 1028 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1710841341
transform 1 0 916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1710841341
transform 1 0 892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1710841341
transform 1 0 1244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1710841341
transform 1 0 1180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1710841341
transform 1 0 1156 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1710841341
transform 1 0 1148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1710841341
transform 1 0 1220 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1710841341
transform 1 0 1188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1710841341
transform 1 0 1180 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1710841341
transform 1 0 1172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1710841341
transform 1 0 1276 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1710841341
transform 1 0 1188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1710841341
transform 1 0 1180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1710841341
transform 1 0 1212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1710841341
transform 1 0 1140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1710841341
transform 1 0 1164 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1710841341
transform 1 0 1132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1710841341
transform 1 0 1276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1710841341
transform 1 0 1220 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1710841341
transform 1 0 1300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1710841341
transform 1 0 1292 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1710841341
transform 1 0 1116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1710841341
transform 1 0 1116 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1710841341
transform 1 0 1196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1710841341
transform 1 0 1172 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1710841341
transform 1 0 1220 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1710841341
transform 1 0 1180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1710841341
transform 1 0 1292 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1710841341
transform 1 0 1204 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1710841341
transform 1 0 1284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1710841341
transform 1 0 1268 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1710841341
transform 1 0 988 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1710841341
transform 1 0 948 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1710841341
transform 1 0 1036 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1710841341
transform 1 0 964 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3699
timestamp 1710841341
transform 1 0 1044 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1710841341
transform 1 0 972 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1710841341
transform 1 0 1108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3702
timestamp 1710841341
transform 1 0 1076 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1710841341
transform 1 0 1068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1710841341
transform 1 0 1068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1710841341
transform 1 0 1124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1710841341
transform 1 0 1092 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3707
timestamp 1710841341
transform 1 0 1468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3708
timestamp 1710841341
transform 1 0 1132 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1710841341
transform 1 0 1084 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1710841341
transform 1 0 1068 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1710841341
transform 1 0 1060 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1710841341
transform 1 0 1052 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1710841341
transform 1 0 1164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1710841341
transform 1 0 1036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1710841341
transform 1 0 1012 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1710841341
transform 1 0 1028 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1710841341
transform 1 0 988 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1710841341
transform 1 0 740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1710841341
transform 1 0 716 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1710841341
transform 1 0 644 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1710841341
transform 1 0 972 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1710841341
transform 1 0 908 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1710841341
transform 1 0 924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1710841341
transform 1 0 916 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1710841341
transform 1 0 908 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1710841341
transform 1 0 884 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1710841341
transform 1 0 1556 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1710841341
transform 1 0 1492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1710841341
transform 1 0 1476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1710841341
transform 1 0 1028 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1710841341
transform 1 0 1020 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1710841341
transform 1 0 1020 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1710841341
transform 1 0 1004 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1710841341
transform 1 0 1068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1710841341
transform 1 0 1012 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1710841341
transform 1 0 868 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1710841341
transform 1 0 788 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1710841341
transform 1 0 812 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1710841341
transform 1 0 788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1710841341
transform 1 0 924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1710841341
transform 1 0 852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1710841341
transform 1 0 924 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1710841341
transform 1 0 924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1710841341
transform 1 0 908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1710841341
transform 1 0 884 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1710841341
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1710841341
transform 1 0 892 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1710841341
transform 1 0 1428 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1710841341
transform 1 0 996 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1710841341
transform 1 0 908 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1710841341
transform 1 0 828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1710841341
transform 1 0 836 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3753
timestamp 1710841341
transform 1 0 836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1710841341
transform 1 0 884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1710841341
transform 1 0 844 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1710841341
transform 1 0 852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1710841341
transform 1 0 828 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1710841341
transform 1 0 812 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1710841341
transform 1 0 780 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1710841341
transform 1 0 764 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1710841341
transform 1 0 940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1710841341
transform 1 0 860 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1710841341
transform 1 0 748 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1710841341
transform 1 0 748 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1710841341
transform 1 0 756 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3766
timestamp 1710841341
transform 1 0 612 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1710841341
transform 1 0 580 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1710841341
transform 1 0 532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1710841341
transform 1 0 780 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1710841341
transform 1 0 716 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1710841341
transform 1 0 828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1710841341
transform 1 0 708 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1710841341
transform 1 0 732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1710841341
transform 1 0 660 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1710841341
transform 1 0 428 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1710841341
transform 1 0 396 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1710841341
transform 1 0 492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1710841341
transform 1 0 444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1710841341
transform 1 0 372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1710841341
transform 1 0 340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1710841341
transform 1 0 508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1710841341
transform 1 0 300 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1710841341
transform 1 0 268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1710841341
transform 1 0 228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3785
timestamp 1710841341
transform 1 0 188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1710841341
transform 1 0 300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1710841341
transform 1 0 276 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1710841341
transform 1 0 196 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1710841341
transform 1 0 196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1710841341
transform 1 0 132 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1710841341
transform 1 0 116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1710841341
transform 1 0 260 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1710841341
transform 1 0 252 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1710841341
transform 1 0 252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1710841341
transform 1 0 276 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1710841341
transform 1 0 204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1710841341
transform 1 0 196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1710841341
transform 1 0 188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1710841341
transform 1 0 172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1710841341
transform 1 0 172 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1710841341
transform 1 0 164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1710841341
transform 1 0 164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1710841341
transform 1 0 148 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1710841341
transform 1 0 140 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1710841341
transform 1 0 212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1710841341
transform 1 0 212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1710841341
transform 1 0 212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3808
timestamp 1710841341
transform 1 0 204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1710841341
transform 1 0 196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1710841341
transform 1 0 188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1710841341
transform 1 0 180 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1710841341
transform 1 0 364 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1710841341
transform 1 0 204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1710841341
transform 1 0 284 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1710841341
transform 1 0 172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1710841341
transform 1 0 348 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1710841341
transform 1 0 180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1710841341
transform 1 0 268 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1710841341
transform 1 0 180 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1710841341
transform 1 0 228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1710841341
transform 1 0 204 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1710841341
transform 1 0 84 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1710841341
transform 1 0 380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1710841341
transform 1 0 292 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1710841341
transform 1 0 220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3826
timestamp 1710841341
transform 1 0 132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1710841341
transform 1 0 108 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1710841341
transform 1 0 108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1710841341
transform 1 0 340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1710841341
transform 1 0 316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1710841341
transform 1 0 180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1710841341
transform 1 0 276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1710841341
transform 1 0 268 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1710841341
transform 1 0 332 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1710841341
transform 1 0 244 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1710841341
transform 1 0 236 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1710841341
transform 1 0 92 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1710841341
transform 1 0 356 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1710841341
transform 1 0 108 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1710841341
transform 1 0 452 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1710841341
transform 1 0 444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1710841341
transform 1 0 348 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1710841341
transform 1 0 292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1710841341
transform 1 0 204 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1710841341
transform 1 0 388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1710841341
transform 1 0 212 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1710841341
transform 1 0 436 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1710841341
transform 1 0 420 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1710841341
transform 1 0 516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1710841341
transform 1 0 420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1710841341
transform 1 0 420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1710841341
transform 1 0 468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1710841341
transform 1 0 284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1710841341
transform 1 0 1228 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1710841341
transform 1 0 1212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1710841341
transform 1 0 1524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1710841341
transform 1 0 1404 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1710841341
transform 1 0 1708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1710841341
transform 1 0 1572 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1710841341
transform 1 0 2148 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1710841341
transform 1 0 2092 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1710841341
transform 1 0 2516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1710841341
transform 1 0 2420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1710841341
transform 1 0 2676 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1710841341
transform 1 0 2580 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1710841341
transform 1 0 2676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1710841341
transform 1 0 2556 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1710841341
transform 1 0 2012 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1710841341
transform 1 0 1916 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1710841341
transform 1 0 2668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1710841341
transform 1 0 2540 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1710841341
transform 1 0 2668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1710841341
transform 1 0 2556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1710841341
transform 1 0 2668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1710841341
transform 1 0 2612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1710841341
transform 1 0 2668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1710841341
transform 1 0 2540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1710841341
transform 1 0 2564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1710841341
transform 1 0 2412 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1710841341
transform 1 0 2508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1710841341
transform 1 0 2364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1710841341
transform 1 0 2532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1710841341
transform 1 0 2404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1710841341
transform 1 0 2084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1710841341
transform 1 0 1956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1710841341
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1710841341
transform 1 0 1948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1710841341
transform 1 0 1716 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1710841341
transform 1 0 1660 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1710841341
transform 1 0 1148 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1710841341
transform 1 0 1092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1710841341
transform 1 0 820 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1710841341
transform 1 0 812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1710841341
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1710841341
transform 1 0 348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1710841341
transform 1 0 252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1710841341
transform 1 0 220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1710841341
transform 1 0 212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1710841341
transform 1 0 204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1710841341
transform 1 0 204 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1710841341
transform 1 0 204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1710841341
transform 1 0 260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1710841341
transform 1 0 244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3904
timestamp 1710841341
transform 1 0 108 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1710841341
transform 1 0 76 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1710841341
transform 1 0 172 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1710841341
transform 1 0 108 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1710841341
transform 1 0 92 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1710841341
transform 1 0 532 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1710841341
transform 1 0 500 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1710841341
transform 1 0 692 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1710841341
transform 1 0 684 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1710841341
transform 1 0 660 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1710841341
transform 1 0 660 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1710841341
transform 1 0 564 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1710841341
transform 1 0 564 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1710841341
transform 1 0 540 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1710841341
transform 1 0 652 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1710841341
transform 1 0 596 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1710841341
transform 1 0 580 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1710841341
transform 1 0 556 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1710841341
transform 1 0 524 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1710841341
transform 1 0 572 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1710841341
transform 1 0 540 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1710841341
transform 1 0 684 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1710841341
transform 1 0 580 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1710841341
transform 1 0 500 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1710841341
transform 1 0 644 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1710841341
transform 1 0 604 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1710841341
transform 1 0 508 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1710841341
transform 1 0 388 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1710841341
transform 1 0 2596 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1710841341
transform 1 0 2596 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1710841341
transform 1 0 2564 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1710841341
transform 1 0 2196 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1710841341
transform 1 0 2148 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1710841341
transform 1 0 2148 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1710841341
transform 1 0 2100 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1710841341
transform 1 0 1980 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1710841341
transform 1 0 1236 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1710841341
transform 1 0 844 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1710841341
transform 1 0 836 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1710841341
transform 1 0 748 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1710841341
transform 1 0 732 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1710841341
transform 1 0 676 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1710841341
transform 1 0 676 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1710841341
transform 1 0 668 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1710841341
transform 1 0 652 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1710841341
transform 1 0 636 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1710841341
transform 1 0 636 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1710841341
transform 1 0 604 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1710841341
transform 1 0 524 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1710841341
transform 1 0 524 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1710841341
transform 1 0 340 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1710841341
transform 1 0 340 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1710841341
transform 1 0 292 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1710841341
transform 1 0 292 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1710841341
transform 1 0 292 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1710841341
transform 1 0 292 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1710841341
transform 1 0 228 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1710841341
transform 1 0 204 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1710841341
transform 1 0 740 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1710841341
transform 1 0 676 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1710841341
transform 1 0 1340 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1710841341
transform 1 0 420 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1710841341
transform 1 0 1452 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1710841341
transform 1 0 1396 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1710841341
transform 1 0 1388 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1710841341
transform 1 0 1388 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1710841341
transform 1 0 1380 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1710841341
transform 1 0 1348 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1710841341
transform 1 0 1348 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1710841341
transform 1 0 492 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1710841341
transform 1 0 348 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1710841341
transform 1 0 340 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1710841341
transform 1 0 1052 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1710841341
transform 1 0 956 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1710841341
transform 1 0 956 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1710841341
transform 1 0 452 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1710841341
transform 1 0 452 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1710841341
transform 1 0 388 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1710841341
transform 1 0 324 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1710841341
transform 1 0 1140 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1710841341
transform 1 0 1092 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1710841341
transform 1 0 1004 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1710841341
transform 1 0 996 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1710841341
transform 1 0 348 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1710841341
transform 1 0 220 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1710841341
transform 1 0 748 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1710841341
transform 1 0 700 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1710841341
transform 1 0 524 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1710841341
transform 1 0 644 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1710841341
transform 1 0 572 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1710841341
transform 1 0 492 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1710841341
transform 1 0 444 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1710841341
transform 1 0 572 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1710841341
transform 1 0 292 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1710841341
transform 1 0 228 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1710841341
transform 1 0 84 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1710841341
transform 1 0 492 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1710841341
transform 1 0 436 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1710841341
transform 1 0 356 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1710841341
transform 1 0 276 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1710841341
transform 1 0 220 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1710841341
transform 1 0 76 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1710841341
transform 1 0 484 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1710841341
transform 1 0 452 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1710841341
transform 1 0 292 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1710841341
transform 1 0 292 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1710841341
transform 1 0 76 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1710841341
transform 1 0 428 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1710841341
transform 1 0 380 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1710841341
transform 1 0 228 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1710841341
transform 1 0 164 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1710841341
transform 1 0 76 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1710841341
transform 1 0 332 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1710841341
transform 1 0 236 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1710841341
transform 1 0 132 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1710841341
transform 1 0 292 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1710841341
transform 1 0 220 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1710841341
transform 1 0 180 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1710841341
transform 1 0 268 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1710841341
transform 1 0 228 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1710841341
transform 1 0 188 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1710841341
transform 1 0 260 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1710841341
transform 1 0 204 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1710841341
transform 1 0 796 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1710841341
transform 1 0 764 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1710841341
transform 1 0 652 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1710841341
transform 1 0 652 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1710841341
transform 1 0 524 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1710841341
transform 1 0 1444 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1710841341
transform 1 0 1404 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1710841341
transform 1 0 1348 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1710841341
transform 1 0 1324 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1710841341
transform 1 0 1260 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1710841341
transform 1 0 2084 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1710841341
transform 1 0 2068 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1710841341
transform 1 0 2060 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1710841341
transform 1 0 2060 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1710841341
transform 1 0 2044 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1710841341
transform 1 0 2028 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1710841341
transform 1 0 2020 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1710841341
transform 1 0 2012 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1710841341
transform 1 0 2012 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1710841341
transform 1 0 1644 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1710841341
transform 1 0 1636 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1710841341
transform 1 0 1636 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1710841341
transform 1 0 1636 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1710841341
transform 1 0 1580 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1710841341
transform 1 0 1580 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1710841341
transform 1 0 1548 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1710841341
transform 1 0 1516 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1710841341
transform 1 0 1452 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1710841341
transform 1 0 1452 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1710841341
transform 1 0 1004 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1710841341
transform 1 0 1004 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1710841341
transform 1 0 972 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1710841341
transform 1 0 972 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1710841341
transform 1 0 932 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1710841341
transform 1 0 892 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1710841341
transform 1 0 844 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1710841341
transform 1 0 828 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1710841341
transform 1 0 796 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1710841341
transform 1 0 708 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1710841341
transform 1 0 1620 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1710841341
transform 1 0 1580 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1710841341
transform 1 0 1316 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1710841341
transform 1 0 1276 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1710841341
transform 1 0 1276 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1710841341
transform 1 0 1164 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1710841341
transform 1 0 1108 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1710841341
transform 1 0 1108 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1710841341
transform 1 0 1108 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1710841341
transform 1 0 1068 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1710841341
transform 1 0 1028 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1710841341
transform 1 0 1532 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1710841341
transform 1 0 1444 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1710841341
transform 1 0 1060 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1710841341
transform 1 0 2044 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1710841341
transform 1 0 1820 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1710841341
transform 1 0 1644 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1710841341
transform 1 0 1588 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1710841341
transform 1 0 1452 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1710841341
transform 1 0 1452 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1710841341
transform 1 0 1324 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1710841341
transform 1 0 1148 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1710841341
transform 1 0 1740 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1710841341
transform 1 0 1700 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1710841341
transform 1 0 1620 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1710841341
transform 1 0 1524 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1710841341
transform 1 0 1452 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1710841341
transform 1 0 1284 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1710841341
transform 1 0 1212 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1710841341
transform 1 0 1964 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1710841341
transform 1 0 1900 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1710841341
transform 1 0 1468 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1710841341
transform 1 0 1396 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1710841341
transform 1 0 1340 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1710841341
transform 1 0 1404 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1710841341
transform 1 0 1356 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1710841341
transform 1 0 1420 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1710841341
transform 1 0 1380 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1710841341
transform 1 0 1348 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1710841341
transform 1 0 1652 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1710841341
transform 1 0 1612 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1710841341
transform 1 0 1516 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1710841341
transform 1 0 1508 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1710841341
transform 1 0 1508 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1710841341
transform 1 0 1436 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1710841341
transform 1 0 1436 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1710841341
transform 1 0 1420 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1710841341
transform 1 0 1420 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1710841341
transform 1 0 1284 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1710841341
transform 1 0 1268 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1710841341
transform 1 0 860 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1710841341
transform 1 0 796 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1710841341
transform 1 0 788 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1710841341
transform 1 0 708 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1710841341
transform 1 0 668 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1710841341
transform 1 0 668 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1710841341
transform 1 0 2644 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1710841341
transform 1 0 1996 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1710841341
transform 1 0 1740 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1710841341
transform 1 0 1756 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1710841341
transform 1 0 1628 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1710841341
transform 1 0 1604 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1710841341
transform 1 0 1572 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1710841341
transform 1 0 1572 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1710841341
transform 1 0 1564 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1710841341
transform 1 0 1524 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1710841341
transform 1 0 1516 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1710841341
transform 1 0 1468 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1710841341
transform 1 0 1092 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1710841341
transform 1 0 684 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1710841341
transform 1 0 492 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1710841341
transform 1 0 220 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1710841341
transform 1 0 1876 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1710841341
transform 1 0 828 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1710841341
transform 1 0 772 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1710841341
transform 1 0 772 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1710841341
transform 1 0 668 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1710841341
transform 1 0 2436 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1710841341
transform 1 0 2276 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1710841341
transform 1 0 2276 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1710841341
transform 1 0 2244 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1710841341
transform 1 0 2204 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1710841341
transform 1 0 2180 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1710841341
transform 1 0 2556 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1710841341
transform 1 0 2436 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1710841341
transform 1 0 2396 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1710841341
transform 1 0 1604 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1710841341
transform 1 0 812 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1710841341
transform 1 0 388 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1710841341
transform 1 0 380 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1710841341
transform 1 0 236 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1710841341
transform 1 0 180 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1710841341
transform 1 0 2220 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1710841341
transform 1 0 1644 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1710841341
transform 1 0 1644 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1710841341
transform 1 0 1644 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1710841341
transform 1 0 1628 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1710841341
transform 1 0 1476 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1710841341
transform 1 0 1316 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1710841341
transform 1 0 1260 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1710841341
transform 1 0 2492 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1710841341
transform 1 0 2484 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1710841341
transform 1 0 2468 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1710841341
transform 1 0 2420 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1710841341
transform 1 0 2380 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1710841341
transform 1 0 2380 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1710841341
transform 1 0 2356 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1710841341
transform 1 0 2340 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1710841341
transform 1 0 2148 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1710841341
transform 1 0 2052 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1710841341
transform 1 0 1876 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1710841341
transform 1 0 1828 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1710841341
transform 1 0 1820 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1710841341
transform 1 0 1492 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1710841341
transform 1 0 948 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1710841341
transform 1 0 948 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1710841341
transform 1 0 900 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1710841341
transform 1 0 2436 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1710841341
transform 1 0 2348 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1710841341
transform 1 0 2308 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1710841341
transform 1 0 2164 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1710841341
transform 1 0 1764 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1710841341
transform 1 0 1764 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1710841341
transform 1 0 1700 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1710841341
transform 1 0 1644 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1710841341
transform 1 0 1604 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1710841341
transform 1 0 1492 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1710841341
transform 1 0 1492 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1710841341
transform 1 0 1404 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1710841341
transform 1 0 1316 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1710841341
transform 1 0 1756 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1710841341
transform 1 0 1716 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1710841341
transform 1 0 2340 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1710841341
transform 1 0 2308 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1710841341
transform 1 0 2308 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1710841341
transform 1 0 2284 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1710841341
transform 1 0 2252 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1710841341
transform 1 0 1412 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1710841341
transform 1 0 1292 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1710841341
transform 1 0 1092 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1710841341
transform 1 0 444 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1710841341
transform 1 0 292 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1710841341
transform 1 0 1508 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1710841341
transform 1 0 476 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1710841341
transform 1 0 2588 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1710841341
transform 1 0 2556 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1710841341
transform 1 0 1796 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1710841341
transform 1 0 1476 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1710841341
transform 1 0 1692 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1710841341
transform 1 0 1620 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1710841341
transform 1 0 1620 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1710841341
transform 1 0 1252 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1710841341
transform 1 0 1276 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1710841341
transform 1 0 1148 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1710841341
transform 1 0 2492 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1710841341
transform 1 0 1996 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1710841341
transform 1 0 1988 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1710841341
transform 1 0 1972 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1710841341
transform 1 0 1964 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1710841341
transform 1 0 2292 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1710841341
transform 1 0 2084 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1710841341
transform 1 0 2084 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1710841341
transform 1 0 1980 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1710841341
transform 1 0 1964 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1710841341
transform 1 0 948 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1710841341
transform 1 0 892 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1710841341
transform 1 0 1748 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1710841341
transform 1 0 1620 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1710841341
transform 1 0 1620 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1710841341
transform 1 0 1508 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1710841341
transform 1 0 1508 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1710841341
transform 1 0 1484 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1710841341
transform 1 0 1444 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1710841341
transform 1 0 1444 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1710841341
transform 1 0 1412 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1710841341
transform 1 0 1148 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1710841341
transform 1 0 996 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1710841341
transform 1 0 380 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1710841341
transform 1 0 228 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1710841341
transform 1 0 180 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1710841341
transform 1 0 1404 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1710841341
transform 1 0 1300 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1710841341
transform 1 0 1292 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1710841341
transform 1 0 1108 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1710841341
transform 1 0 1028 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1710841341
transform 1 0 1020 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1710841341
transform 1 0 956 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1710841341
transform 1 0 956 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1710841341
transform 1 0 2644 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1710841341
transform 1 0 2548 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1710841341
transform 1 0 2476 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1710841341
transform 1 0 2140 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1710841341
transform 1 0 2132 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1710841341
transform 1 0 2108 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1710841341
transform 1 0 2060 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1710841341
transform 1 0 1516 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1710841341
transform 1 0 1460 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1710841341
transform 1 0 2260 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1710841341
transform 1 0 2004 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1710841341
transform 1 0 1492 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1710841341
transform 1 0 1492 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1710841341
transform 1 0 1468 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1710841341
transform 1 0 1412 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1710841341
transform 1 0 1388 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1710841341
transform 1 0 1356 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1710841341
transform 1 0 1348 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1710841341
transform 1 0 1556 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1710841341
transform 1 0 1284 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1710841341
transform 1 0 564 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1710841341
transform 1 0 484 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1710841341
transform 1 0 436 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1710841341
transform 1 0 2356 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1710841341
transform 1 0 2324 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1710841341
transform 1 0 2564 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1710841341
transform 1 0 2508 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1710841341
transform 1 0 1612 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1710841341
transform 1 0 1492 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1710841341
transform 1 0 1412 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1710841341
transform 1 0 772 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1710841341
transform 1 0 772 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1710841341
transform 1 0 700 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1710841341
transform 1 0 692 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1710841341
transform 1 0 676 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1710841341
transform 1 0 612 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1710841341
transform 1 0 700 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1710841341
transform 1 0 660 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1710841341
transform 1 0 596 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1710841341
transform 1 0 572 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1710841341
transform 1 0 540 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1710841341
transform 1 0 684 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1710841341
transform 1 0 628 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1710841341
transform 1 0 532 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1710841341
transform 1 0 644 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1710841341
transform 1 0 588 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1710841341
transform 1 0 444 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1710841341
transform 1 0 2092 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1710841341
transform 1 0 2068 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1710841341
transform 1 0 2044 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1710841341
transform 1 0 1980 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1710841341
transform 1 0 1540 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1710841341
transform 1 0 1356 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1710841341
transform 1 0 2564 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1710841341
transform 1 0 2276 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1710841341
transform 1 0 2260 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1710841341
transform 1 0 2244 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1710841341
transform 1 0 2012 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1710841341
transform 1 0 1828 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1710841341
transform 1 0 1708 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1710841341
transform 1 0 1972 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1710841341
transform 1 0 1236 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1710841341
transform 1 0 1204 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1710841341
transform 1 0 1188 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1710841341
transform 1 0 1180 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1710841341
transform 1 0 1164 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1710841341
transform 1 0 996 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1710841341
transform 1 0 980 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1710841341
transform 1 0 972 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1710841341
transform 1 0 916 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1710841341
transform 1 0 900 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1710841341
transform 1 0 900 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1710841341
transform 1 0 1572 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1710841341
transform 1 0 1548 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1710841341
transform 1 0 1340 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1710841341
transform 1 0 1340 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1710841341
transform 1 0 1148 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1710841341
transform 1 0 1148 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1710841341
transform 1 0 924 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1710841341
transform 1 0 852 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1710841341
transform 1 0 2100 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1710841341
transform 1 0 2068 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1710841341
transform 1 0 1028 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1710841341
transform 1 0 932 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1710841341
transform 1 0 844 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1710841341
transform 1 0 1604 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1710841341
transform 1 0 1276 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1710841341
transform 1 0 1276 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1710841341
transform 1 0 1228 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1710841341
transform 1 0 1212 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1710841341
transform 1 0 1068 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1710841341
transform 1 0 1012 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1710841341
transform 1 0 812 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1710841341
transform 1 0 804 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1710841341
transform 1 0 756 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1710841341
transform 1 0 884 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1710841341
transform 1 0 804 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1710841341
transform 1 0 804 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1710841341
transform 1 0 740 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1710841341
transform 1 0 2068 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1710841341
transform 1 0 2004 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1710841341
transform 1 0 2004 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1710841341
transform 1 0 1900 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1710841341
transform 1 0 1900 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1710841341
transform 1 0 1708 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1710841341
transform 1 0 1620 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1710841341
transform 1 0 1308 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1710841341
transform 1 0 1308 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1710841341
transform 1 0 1252 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1710841341
transform 1 0 644 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1710841341
transform 1 0 588 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1710841341
transform 1 0 1820 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1710841341
transform 1 0 1676 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1710841341
transform 1 0 836 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1710841341
transform 1 0 828 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1710841341
transform 1 0 564 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1710841341
transform 1 0 1996 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1710841341
transform 1 0 1924 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1710841341
transform 1 0 1500 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1710841341
transform 1 0 1500 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1710841341
transform 1 0 1092 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1710841341
transform 1 0 1084 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1710841341
transform 1 0 996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1710841341
transform 1 0 996 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1710841341
transform 1 0 948 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1710841341
transform 1 0 940 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1710841341
transform 1 0 996 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1710841341
transform 1 0 892 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1710841341
transform 1 0 796 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1710841341
transform 1 0 2076 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1710841341
transform 1 0 2036 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1710841341
transform 1 0 1964 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1710841341
transform 1 0 1964 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1710841341
transform 1 0 2140 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1710841341
transform 1 0 2140 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1710841341
transform 1 0 2100 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1710841341
transform 1 0 2100 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1710841341
transform 1 0 2068 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1710841341
transform 1 0 996 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1710841341
transform 1 0 836 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1710841341
transform 1 0 796 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1710841341
transform 1 0 1804 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1710841341
transform 1 0 1364 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1710841341
transform 1 0 1316 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1710841341
transform 1 0 1308 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1710841341
transform 1 0 1204 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1710841341
transform 1 0 1116 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1710841341
transform 1 0 1076 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1710841341
transform 1 0 1076 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1710841341
transform 1 0 948 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1710841341
transform 1 0 836 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1710841341
transform 1 0 732 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1710841341
transform 1 0 1652 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1710841341
transform 1 0 1404 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1710841341
transform 1 0 1404 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1710841341
transform 1 0 1300 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1710841341
transform 1 0 1300 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1710841341
transform 1 0 1252 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1710841341
transform 1 0 924 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1710841341
transform 1 0 892 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1710841341
transform 1 0 892 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1710841341
transform 1 0 764 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1710841341
transform 1 0 756 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1710841341
transform 1 0 1076 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1710841341
transform 1 0 828 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1710841341
transform 1 0 596 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1710841341
transform 1 0 2116 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1710841341
transform 1 0 2052 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1710841341
transform 1 0 2052 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1710841341
transform 1 0 1996 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1710841341
transform 1 0 1732 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1710841341
transform 1 0 1732 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1710841341
transform 1 0 1620 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1710841341
transform 1 0 2516 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1710841341
transform 1 0 2204 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1710841341
transform 1 0 2204 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1710841341
transform 1 0 2100 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1710841341
transform 1 0 1956 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1710841341
transform 1 0 1876 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1710841341
transform 1 0 1532 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1710841341
transform 1 0 1508 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1710841341
transform 1 0 1220 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1710841341
transform 1 0 1580 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1710841341
transform 1 0 1420 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1710841341
transform 1 0 1420 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1710841341
transform 1 0 1348 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1710841341
transform 1 0 964 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1710841341
transform 1 0 740 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1710841341
transform 1 0 2028 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1710841341
transform 1 0 1964 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1710841341
transform 1 0 2156 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1710841341
transform 1 0 2020 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1710841341
transform 1 0 2020 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1710841341
transform 1 0 1676 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1710841341
transform 1 0 1588 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1710841341
transform 1 0 1452 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1710841341
transform 1 0 236 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1710841341
transform 1 0 204 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1710841341
transform 1 0 308 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1710841341
transform 1 0 236 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1710841341
transform 1 0 196 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1710841341
transform 1 0 260 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1710841341
transform 1 0 188 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1710841341
transform 1 0 188 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1710841341
transform 1 0 164 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1710841341
transform 1 0 660 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1710841341
transform 1 0 452 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1710841341
transform 1 0 708 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1710841341
transform 1 0 548 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1710841341
transform 1 0 636 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1710841341
transform 1 0 484 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1710841341
transform 1 0 1124 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1710841341
transform 1 0 1060 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1710841341
transform 1 0 1060 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1710841341
transform 1 0 900 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1710841341
transform 1 0 892 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1710841341
transform 1 0 764 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1710841341
transform 1 0 788 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1710841341
transform 1 0 700 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1710841341
transform 1 0 940 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1710841341
transform 1 0 892 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1710841341
transform 1 0 1340 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1710841341
transform 1 0 1268 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1710841341
transform 1 0 588 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1710841341
transform 1 0 532 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1710841341
transform 1 0 1116 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1710841341
transform 1 0 1052 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1710841341
transform 1 0 1220 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1710841341
transform 1 0 1140 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1710841341
transform 1 0 1700 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1710841341
transform 1 0 1612 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1710841341
transform 1 0 1556 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1710841341
transform 1 0 1556 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1710841341
transform 1 0 1524 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1710841341
transform 1 0 1796 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1710841341
transform 1 0 1692 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1710841341
transform 1 0 1684 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1710841341
transform 1 0 1548 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1710841341
transform 1 0 1932 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1710841341
transform 1 0 1892 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1710841341
transform 1 0 1956 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1710841341
transform 1 0 1892 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1710841341
transform 1 0 1484 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1710841341
transform 1 0 1452 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1710841341
transform 1 0 1916 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1710841341
transform 1 0 1876 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1710841341
transform 1 0 1940 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1710841341
transform 1 0 1516 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1710841341
transform 1 0 1428 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1710841341
transform 1 0 2348 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1710841341
transform 1 0 2172 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1710841341
transform 1 0 2404 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1710841341
transform 1 0 2372 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1710841341
transform 1 0 2340 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1710841341
transform 1 0 2308 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1710841341
transform 1 0 2164 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1710841341
transform 1 0 2124 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1710841341
transform 1 0 2252 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1710841341
transform 1 0 2092 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1710841341
transform 1 0 2148 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1710841341
transform 1 0 2060 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1710841341
transform 1 0 2172 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1710841341
transform 1 0 2140 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1710841341
transform 1 0 2596 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1710841341
transform 1 0 2540 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1710841341
transform 1 0 2444 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1710841341
transform 1 0 2316 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1710841341
transform 1 0 2220 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1710841341
transform 1 0 2156 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1710841341
transform 1 0 2436 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1710841341
transform 1 0 2396 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1710841341
transform 1 0 2308 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1710841341
transform 1 0 2284 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1710841341
transform 1 0 2228 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1710841341
transform 1 0 2172 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1710841341
transform 1 0 2020 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1710841341
transform 1 0 2324 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1710841341
transform 1 0 2308 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1710841341
transform 1 0 2516 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1710841341
transform 1 0 2484 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1710841341
transform 1 0 2300 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1710841341
transform 1 0 2292 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1710841341
transform 1 0 2148 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1710841341
transform 1 0 1756 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1710841341
transform 1 0 1716 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1710841341
transform 1 0 2084 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1710841341
transform 1 0 1724 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1710841341
transform 1 0 2452 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1710841341
transform 1 0 2388 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1710841341
transform 1 0 2596 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1710841341
transform 1 0 2564 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1710841341
transform 1 0 2268 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1710841341
transform 1 0 2228 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1710841341
transform 1 0 1844 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1710841341
transform 1 0 1828 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1710841341
transform 1 0 1988 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1710841341
transform 1 0 1948 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1710841341
transform 1 0 2116 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1710841341
transform 1 0 1988 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1710841341
transform 1 0 2044 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1710841341
transform 1 0 1940 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1710841341
transform 1 0 1684 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1710841341
transform 1 0 1652 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1710841341
transform 1 0 1748 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1710841341
transform 1 0 1660 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1710841341
transform 1 0 1796 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1710841341
transform 1 0 1756 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1710841341
transform 1 0 1164 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1710841341
transform 1 0 1124 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1710841341
transform 1 0 1084 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1710841341
transform 1 0 700 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1710841341
transform 1 0 700 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1710841341
transform 1 0 660 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1710841341
transform 1 0 564 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1710841341
transform 1 0 476 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1710841341
transform 1 0 1468 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1710841341
transform 1 0 1340 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1710841341
transform 1 0 1340 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1710841341
transform 1 0 1340 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1710841341
transform 1 0 1332 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1710841341
transform 1 0 1300 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1710841341
transform 1 0 1284 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1710841341
transform 1 0 1268 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1710841341
transform 1 0 1212 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1710841341
transform 1 0 1108 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1710841341
transform 1 0 908 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1710841341
transform 1 0 892 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1710841341
transform 1 0 892 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1710841341
transform 1 0 412 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1710841341
transform 1 0 396 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1710841341
transform 1 0 396 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1710841341
transform 1 0 372 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1710841341
transform 1 0 332 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1710841341
transform 1 0 172 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1710841341
transform 1 0 164 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1710841341
transform 1 0 108 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1710841341
transform 1 0 1004 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1710841341
transform 1 0 964 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1710841341
transform 1 0 2380 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1710841341
transform 1 0 2300 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1710841341
transform 1 0 2332 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1710841341
transform 1 0 2284 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1710841341
transform 1 0 1484 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1710841341
transform 1 0 1484 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1710841341
transform 1 0 1020 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1710841341
transform 1 0 1020 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1710841341
transform 1 0 772 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1710841341
transform 1 0 2172 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1710841341
transform 1 0 1508 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1710841341
transform 1 0 1508 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1710841341
transform 1 0 1380 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1710841341
transform 1 0 1356 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1710841341
transform 1 0 1356 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1710841341
transform 1 0 1004 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1710841341
transform 1 0 1540 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1710841341
transform 1 0 1468 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1710841341
transform 1 0 1468 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1710841341
transform 1 0 1396 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1710841341
transform 1 0 1220 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1710841341
transform 1 0 1156 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1710841341
transform 1 0 164 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1710841341
transform 1 0 84 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1710841341
transform 1 0 308 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1710841341
transform 1 0 244 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1710841341
transform 1 0 188 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1710841341
transform 1 0 140 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1710841341
transform 1 0 116 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1710841341
transform 1 0 76 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1710841341
transform 1 0 460 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1710841341
transform 1 0 364 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1710841341
transform 1 0 372 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1710841341
transform 1 0 332 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1710841341
transform 1 0 2620 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1710841341
transform 1 0 2556 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1710841341
transform 1 0 2548 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1710841341
transform 1 0 2540 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1710841341
transform 1 0 2500 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1710841341
transform 1 0 2476 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1710841341
transform 1 0 2380 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1710841341
transform 1 0 2380 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1710841341
transform 1 0 2356 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1710841341
transform 1 0 2284 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1710841341
transform 1 0 2244 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1710841341
transform 1 0 2076 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1710841341
transform 1 0 1900 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1710841341
transform 1 0 1884 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1710841341
transform 1 0 1884 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1710841341
transform 1 0 1812 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1710841341
transform 1 0 1756 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1710841341
transform 1 0 1756 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1710841341
transform 1 0 1444 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1710841341
transform 1 0 1444 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1710841341
transform 1 0 1332 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1710841341
transform 1 0 1284 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1710841341
transform 1 0 908 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1710841341
transform 1 0 668 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1710841341
transform 1 0 636 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1710841341
transform 1 0 524 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1710841341
transform 1 0 500 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1710841341
transform 1 0 316 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1710841341
transform 1 0 316 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1710841341
transform 1 0 92 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1710841341
transform 1 0 68 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1710841341
transform 1 0 68 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1710841341
transform 1 0 2108 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1710841341
transform 1 0 2076 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1710841341
transform 1 0 2076 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1710841341
transform 1 0 1996 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1710841341
transform 1 0 1900 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1710841341
transform 1 0 1892 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1710841341
transform 1 0 1596 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1710841341
transform 1 0 1500 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1710841341
transform 1 0 1212 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1710841341
transform 1 0 1148 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1710841341
transform 1 0 1140 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1710841341
transform 1 0 1084 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1710841341
transform 1 0 868 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1710841341
transform 1 0 852 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1710841341
transform 1 0 756 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1710841341
transform 1 0 716 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1710841341
transform 1 0 684 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1710841341
transform 1 0 676 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1710841341
transform 1 0 636 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1710841341
transform 1 0 628 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1710841341
transform 1 0 628 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1710841341
transform 1 0 620 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1710841341
transform 1 0 2620 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1710841341
transform 1 0 2572 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1710841341
transform 1 0 2540 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1710841341
transform 1 0 2516 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1710841341
transform 1 0 2252 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1710841341
transform 1 0 2220 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1710841341
transform 1 0 2220 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1710841341
transform 1 0 2220 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1710841341
transform 1 0 2036 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1710841341
transform 1 0 2036 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1710841341
transform 1 0 2036 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1710841341
transform 1 0 2004 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1710841341
transform 1 0 1980 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1710841341
transform 1 0 1964 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1710841341
transform 1 0 1948 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1710841341
transform 1 0 1932 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1710841341
transform 1 0 1908 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1710841341
transform 1 0 1908 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1710841341
transform 1 0 1884 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1710841341
transform 1 0 1884 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1710841341
transform 1 0 1580 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1710841341
transform 1 0 1556 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1710841341
transform 1 0 1516 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1710841341
transform 1 0 1516 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1710841341
transform 1 0 1476 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1710841341
transform 1 0 1252 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1710841341
transform 1 0 1172 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1710841341
transform 1 0 1084 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1710841341
transform 1 0 1084 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1710841341
transform 1 0 1052 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1710841341
transform 1 0 852 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1710841341
transform 1 0 2476 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1710841341
transform 1 0 2452 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1710841341
transform 1 0 2244 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1710841341
transform 1 0 2172 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1710841341
transform 1 0 2172 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1710841341
transform 1 0 2092 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1710841341
transform 1 0 2044 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1710841341
transform 1 0 1924 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1710841341
transform 1 0 1924 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1710841341
transform 1 0 1588 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1710841341
transform 1 0 1588 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1710841341
transform 1 0 1500 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1710841341
transform 1 0 996 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1710841341
transform 1 0 820 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1710841341
transform 1 0 692 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1710841341
transform 1 0 524 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1710841341
transform 1 0 516 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1710841341
transform 1 0 476 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1710841341
transform 1 0 428 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1710841341
transform 1 0 428 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1710841341
transform 1 0 420 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1710841341
transform 1 0 388 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1710841341
transform 1 0 356 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1710841341
transform 1 0 316 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1710841341
transform 1 0 316 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1710841341
transform 1 0 308 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1710841341
transform 1 0 2628 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1710841341
transform 1 0 2596 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1710841341
transform 1 0 2572 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1710841341
transform 1 0 2420 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1710841341
transform 1 0 2420 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1710841341
transform 1 0 2380 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1710841341
transform 1 0 2372 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1710841341
transform 1 0 2364 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1710841341
transform 1 0 2332 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1710841341
transform 1 0 2020 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1710841341
transform 1 0 1804 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1710841341
transform 1 0 1804 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1710841341
transform 1 0 1796 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1710841341
transform 1 0 1764 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1710841341
transform 1 0 1764 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1710841341
transform 1 0 1660 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1710841341
transform 1 0 1652 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1710841341
transform 1 0 1356 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1710841341
transform 1 0 1348 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1710841341
transform 1 0 1204 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1710841341
transform 1 0 1156 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1710841341
transform 1 0 1116 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1710841341
transform 1 0 1004 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1710841341
transform 1 0 1004 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1710841341
transform 1 0 932 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1710841341
transform 1 0 932 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1710841341
transform 1 0 644 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1710841341
transform 1 0 644 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1710841341
transform 1 0 548 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1710841341
transform 1 0 548 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1710841341
transform 1 0 412 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1710841341
transform 1 0 332 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1710841341
transform 1 0 332 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1710841341
transform 1 0 212 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1710841341
transform 1 0 196 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1710841341
transform 1 0 196 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1710841341
transform 1 0 2668 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1710841341
transform 1 0 2644 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1710841341
transform 1 0 2572 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1710841341
transform 1 0 2516 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1710841341
transform 1 0 2508 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1710841341
transform 1 0 2484 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1710841341
transform 1 0 2332 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1710841341
transform 1 0 2300 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1710841341
transform 1 0 2204 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1710841341
transform 1 0 1852 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1710841341
transform 1 0 1732 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1710841341
transform 1 0 1396 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1710841341
transform 1 0 1340 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1710841341
transform 1 0 1284 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1710841341
transform 1 0 1204 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1710841341
transform 1 0 1004 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1710841341
transform 1 0 908 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1710841341
transform 1 0 868 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1710841341
transform 1 0 484 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1710841341
transform 1 0 2676 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1710841341
transform 1 0 2676 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1710841341
transform 1 0 2564 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1710841341
transform 1 0 2468 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1710841341
transform 1 0 2428 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1710841341
transform 1 0 2428 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1710841341
transform 1 0 2372 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1710841341
transform 1 0 2052 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1710841341
transform 1 0 1988 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1710841341
transform 1 0 1652 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1710841341
transform 1 0 1644 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1710841341
transform 1 0 1644 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1710841341
transform 1 0 1612 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1710841341
transform 1 0 1612 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1710841341
transform 1 0 1612 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1710841341
transform 1 0 1564 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1710841341
transform 1 0 1540 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1710841341
transform 1 0 1476 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1710841341
transform 1 0 1468 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1710841341
transform 1 0 1444 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1710841341
transform 1 0 1444 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1710841341
transform 1 0 1252 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1710841341
transform 1 0 1252 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1710841341
transform 1 0 1228 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1710841341
transform 1 0 1212 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1710841341
transform 1 0 1140 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1710841341
transform 1 0 916 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1710841341
transform 1 0 916 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1710841341
transform 1 0 708 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1710841341
transform 1 0 1668 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1710841341
transform 1 0 1612 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1710841341
transform 1 0 1604 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1710841341
transform 1 0 1372 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1710841341
transform 1 0 1156 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1710841341
transform 1 0 932 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1710841341
transform 1 0 932 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1710841341
transform 1 0 836 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1710841341
transform 1 0 812 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1710841341
transform 1 0 812 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1710841341
transform 1 0 764 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1710841341
transform 1 0 764 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1710841341
transform 1 0 2100 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1710841341
transform 1 0 2092 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1710841341
transform 1 0 2060 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1710841341
transform 1 0 2060 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1710841341
transform 1 0 2052 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1710841341
transform 1 0 2052 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1710841341
transform 1 0 2044 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1710841341
transform 1 0 2044 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1710841341
transform 1 0 2020 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1710841341
transform 1 0 2020 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1710841341
transform 1 0 2012 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1710841341
transform 1 0 1636 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1710841341
transform 1 0 1436 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1710841341
transform 1 0 1244 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1710841341
transform 1 0 1060 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1710841341
transform 1 0 988 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1710841341
transform 1 0 956 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1710841341
transform 1 0 940 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1710841341
transform 1 0 940 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1710841341
transform 1 0 932 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1710841341
transform 1 0 876 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1710841341
transform 1 0 852 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1710841341
transform 1 0 852 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1710841341
transform 1 0 820 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1710841341
transform 1 0 812 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1710841341
transform 1 0 796 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1710841341
transform 1 0 788 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1710841341
transform 1 0 2244 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1710841341
transform 1 0 2164 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1710841341
transform 1 0 2124 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1710841341
transform 1 0 2100 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1710841341
transform 1 0 1492 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1710841341
transform 1 0 1236 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1710841341
transform 1 0 1196 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1710841341
transform 1 0 948 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1710841341
transform 1 0 860 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1710841341
transform 1 0 2132 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1710841341
transform 1 0 2100 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1710841341
transform 1 0 2084 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1710841341
transform 1 0 2084 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1710841341
transform 1 0 2084 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1710841341
transform 1 0 2036 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1710841341
transform 1 0 2036 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1710841341
transform 1 0 2028 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1710841341
transform 1 0 1980 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1710841341
transform 1 0 1980 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1710841341
transform 1 0 1940 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1710841341
transform 1 0 1940 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1710841341
transform 1 0 1924 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1710841341
transform 1 0 1916 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1710841341
transform 1 0 1604 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1710841341
transform 1 0 1364 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1710841341
transform 1 0 1364 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1710841341
transform 1 0 1220 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1710841341
transform 1 0 972 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1710841341
transform 1 0 956 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1710841341
transform 1 0 900 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1710841341
transform 1 0 868 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1710841341
transform 1 0 836 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1710841341
transform 1 0 836 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1710841341
transform 1 0 764 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1710841341
transform 1 0 764 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1710841341
transform 1 0 708 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1710841341
transform 1 0 692 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1710841341
transform 1 0 692 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1710841341
transform 1 0 2604 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1710841341
transform 1 0 2468 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1710841341
transform 1 0 2460 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1710841341
transform 1 0 2436 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1710841341
transform 1 0 2412 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1710841341
transform 1 0 2100 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1710841341
transform 1 0 1380 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1710841341
transform 1 0 1380 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1710841341
transform 1 0 1236 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1710841341
transform 1 0 1908 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1710841341
transform 1 0 1820 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1710841341
transform 1 0 1780 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1710841341
transform 1 0 1756 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1710841341
transform 1 0 1692 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1710841341
transform 1 0 2092 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1710841341
transform 1 0 1948 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1710841341
transform 1 0 1364 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1710841341
transform 1 0 1364 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1710841341
transform 1 0 1220 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1710841341
transform 1 0 1212 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1710841341
transform 1 0 1180 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1710841341
transform 1 0 2300 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1710841341
transform 1 0 2252 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1710841341
transform 1 0 2252 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1710841341
transform 1 0 1916 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1710841341
transform 1 0 1860 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1710841341
transform 1 0 1860 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1710841341
transform 1 0 1380 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1710841341
transform 1 0 2508 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1710841341
transform 1 0 2460 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1710841341
transform 1 0 2460 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1710841341
transform 1 0 1228 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1710841341
transform 1 0 1212 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1710841341
transform 1 0 636 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1710841341
transform 1 0 2468 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1710841341
transform 1 0 1796 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1710841341
transform 1 0 1740 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1710841341
transform 1 0 1732 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1710841341
transform 1 0 1308 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1710841341
transform 1 0 2500 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1710841341
transform 1 0 2500 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1710841341
transform 1 0 2452 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1710841341
transform 1 0 2428 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1710841341
transform 1 0 2324 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1710841341
transform 1 0 2324 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1710841341
transform 1 0 2252 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1710841341
transform 1 0 1316 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1710841341
transform 1 0 412 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1710841341
transform 1 0 364 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1710841341
transform 1 0 2052 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1710841341
transform 1 0 1924 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1710841341
transform 1 0 1772 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1710841341
transform 1 0 1748 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1710841341
transform 1 0 1732 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1710841341
transform 1 0 1724 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1710841341
transform 1 0 1668 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1710841341
transform 1 0 1668 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1710841341
transform 1 0 1556 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1710841341
transform 1 0 1548 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1710841341
transform 1 0 1388 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1710841341
transform 1 0 1388 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1710841341
transform 1 0 612 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1710841341
transform 1 0 1348 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1710841341
transform 1 0 1292 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1710841341
transform 1 0 2396 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1710841341
transform 1 0 2396 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1710841341
transform 1 0 2324 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1710841341
transform 1 0 2300 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1710841341
transform 1 0 2172 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1710841341
transform 1 0 2164 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1710841341
transform 1 0 2164 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1710841341
transform 1 0 2132 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1710841341
transform 1 0 2108 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1710841341
transform 1 0 2028 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1710841341
transform 1 0 1772 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1710841341
transform 1 0 1548 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1710841341
transform 1 0 1516 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1710841341
transform 1 0 1492 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1710841341
transform 1 0 1476 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1710841341
transform 1 0 1116 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1710841341
transform 1 0 1116 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1710841341
transform 1 0 540 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1710841341
transform 1 0 420 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1710841341
transform 1 0 2428 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1710841341
transform 1 0 2364 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1710841341
transform 1 0 2356 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1710841341
transform 1 0 2164 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1710841341
transform 1 0 1844 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1710841341
transform 1 0 1180 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1710841341
transform 1 0 1108 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1710841341
transform 1 0 1108 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1710841341
transform 1 0 1484 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1710841341
transform 1 0 1220 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1710841341
transform 1 0 1204 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1710841341
transform 1 0 1124 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1710841341
transform 1 0 1108 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1710841341
transform 1 0 708 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1710841341
transform 1 0 356 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1710841341
transform 1 0 2372 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1710841341
transform 1 0 2356 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1710841341
transform 1 0 2284 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1710841341
transform 1 0 2276 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1710841341
transform 1 0 2140 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1710841341
transform 1 0 1260 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1710841341
transform 1 0 1260 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1710841341
transform 1 0 1164 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1710841341
transform 1 0 1148 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1710841341
transform 1 0 1100 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1710841341
transform 1 0 1092 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1710841341
transform 1 0 956 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1710841341
transform 1 0 2452 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1710841341
transform 1 0 2444 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1710841341
transform 1 0 2444 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1710841341
transform 1 0 2420 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1710841341
transform 1 0 2404 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1710841341
transform 1 0 2404 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1710841341
transform 1 0 2348 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1710841341
transform 1 0 2332 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1710841341
transform 1 0 2332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1710841341
transform 1 0 2308 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1710841341
transform 1 0 2300 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1710841341
transform 1 0 2260 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1710841341
transform 1 0 2148 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1710841341
transform 1 0 2068 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1710841341
transform 1 0 2012 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1710841341
transform 1 0 1868 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1710841341
transform 1 0 1868 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1710841341
transform 1 0 1828 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1710841341
transform 1 0 1828 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1710841341
transform 1 0 1828 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1710841341
transform 1 0 1820 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1710841341
transform 1 0 1780 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1710841341
transform 1 0 1652 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1710841341
transform 1 0 1636 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1710841341
transform 1 0 1572 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1710841341
transform 1 0 1556 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1710841341
transform 1 0 1476 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1710841341
transform 1 0 1196 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1710841341
transform 1 0 1196 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1710841341
transform 1 0 1132 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1710841341
transform 1 0 1132 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1710841341
transform 1 0 1076 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1710841341
transform 1 0 564 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1710841341
transform 1 0 1884 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1710841341
transform 1 0 1788 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1710841341
transform 1 0 1708 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1710841341
transform 1 0 1668 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1710841341
transform 1 0 1668 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1710841341
transform 1 0 1620 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1710841341
transform 1 0 1164 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1710841341
transform 1 0 1068 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1710841341
transform 1 0 1004 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1710841341
transform 1 0 940 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1710841341
transform 1 0 692 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1710841341
transform 1 0 572 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1710841341
transform 1 0 2476 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1710841341
transform 1 0 2476 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1710841341
transform 1 0 2436 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1710841341
transform 1 0 2436 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1710841341
transform 1 0 2388 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1710841341
transform 1 0 2380 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1710841341
transform 1 0 2340 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1710841341
transform 1 0 2332 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1710841341
transform 1 0 2316 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1710841341
transform 1 0 2268 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1710841341
transform 1 0 2260 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1710841341
transform 1 0 2116 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1710841341
transform 1 0 2116 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1710841341
transform 1 0 2108 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1710841341
transform 1 0 2108 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1710841341
transform 1 0 2068 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1710841341
transform 1 0 2012 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1710841341
transform 1 0 1980 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1710841341
transform 1 0 1972 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1710841341
transform 1 0 1972 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1710841341
transform 1 0 1972 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1710841341
transform 1 0 1804 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1710841341
transform 1 0 1796 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1710841341
transform 1 0 1780 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1710841341
transform 1 0 1772 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1710841341
transform 1 0 1764 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1710841341
transform 1 0 1620 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1710841341
transform 1 0 1388 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1710841341
transform 1 0 1196 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1710841341
transform 1 0 1196 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1710841341
transform 1 0 628 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1710841341
transform 1 0 572 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1710841341
transform 1 0 564 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1710841341
transform 1 0 540 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1710841341
transform 1 0 524 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1710841341
transform 1 0 516 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1710841341
transform 1 0 1692 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1710841341
transform 1 0 1684 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1710841341
transform 1 0 1620 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1710841341
transform 1 0 1580 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1710841341
transform 1 0 1356 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1710841341
transform 1 0 876 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1710841341
transform 1 0 876 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1710841341
transform 1 0 836 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1710841341
transform 1 0 804 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1710841341
transform 1 0 2644 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1710841341
transform 1 0 2612 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1710841341
transform 1 0 2588 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1710841341
transform 1 0 2420 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1710841341
transform 1 0 2380 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1710841341
transform 1 0 2364 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1710841341
transform 1 0 2036 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1710841341
transform 1 0 1820 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1710841341
transform 1 0 1812 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1710841341
transform 1 0 1812 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1710841341
transform 1 0 1732 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1710841341
transform 1 0 1724 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1710841341
transform 1 0 1684 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1710841341
transform 1 0 1684 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1710841341
transform 1 0 1676 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1710841341
transform 1 0 1468 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1710841341
transform 1 0 1284 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1710841341
transform 1 0 1236 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1710841341
transform 1 0 1172 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1710841341
transform 1 0 948 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1710841341
transform 1 0 924 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1710841341
transform 1 0 916 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1710841341
transform 1 0 524 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1710841341
transform 1 0 516 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1710841341
transform 1 0 516 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1710841341
transform 1 0 436 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1710841341
transform 1 0 436 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1710841341
transform 1 0 404 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1710841341
transform 1 0 372 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1710841341
transform 1 0 372 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1710841341
transform 1 0 324 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1710841341
transform 1 0 316 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1710841341
transform 1 0 1636 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1710841341
transform 1 0 1540 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1710841341
transform 1 0 1484 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1710841341
transform 1 0 1276 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1710841341
transform 1 0 908 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1710841341
transform 1 0 796 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1710841341
transform 1 0 756 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1710841341
transform 1 0 716 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1710841341
transform 1 0 2204 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1710841341
transform 1 0 1660 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1710841341
transform 1 0 1012 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1710841341
transform 1 0 964 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1710841341
transform 1 0 748 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1710841341
transform 1 0 748 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1710841341
transform 1 0 740 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1710841341
transform 1 0 740 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1710841341
transform 1 0 732 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1710841341
transform 1 0 708 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1710841341
transform 1 0 660 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1710841341
transform 1 0 548 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1710841341
transform 1 0 2364 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1710841341
transform 1 0 2364 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1710841341
transform 1 0 2308 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1710841341
transform 1 0 2236 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1710841341
transform 1 0 1828 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1710841341
transform 1 0 1820 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1710841341
transform 1 0 892 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1710841341
transform 1 0 892 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1710841341
transform 1 0 868 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1710841341
transform 1 0 740 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1710841341
transform 1 0 2372 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1710841341
transform 1 0 2332 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1710841341
transform 1 0 2324 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1710841341
transform 1 0 2300 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1710841341
transform 1 0 2292 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1710841341
transform 1 0 2292 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1710841341
transform 1 0 2260 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1710841341
transform 1 0 2260 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1710841341
transform 1 0 2212 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1710841341
transform 1 0 2172 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1710841341
transform 1 0 2124 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1710841341
transform 1 0 1916 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1710841341
transform 1 0 1916 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1710841341
transform 1 0 1564 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1710841341
transform 1 0 1444 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1710841341
transform 1 0 1052 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1710841341
transform 1 0 1052 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1710841341
transform 1 0 780 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1710841341
transform 1 0 780 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1710841341
transform 1 0 732 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1710841341
transform 1 0 708 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1710841341
transform 1 0 516 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1710841341
transform 1 0 516 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1710841341
transform 1 0 508 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1710841341
transform 1 0 460 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1710841341
transform 1 0 460 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1710841341
transform 1 0 340 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1710841341
transform 1 0 292 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1710841341
transform 1 0 292 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1710841341
transform 1 0 284 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1710841341
transform 1 0 276 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1710841341
transform 1 0 276 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1710841341
transform 1 0 252 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1710841341
transform 1 0 2620 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1710841341
transform 1 0 2588 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1710841341
transform 1 0 2588 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1710841341
transform 1 0 2588 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1710841341
transform 1 0 2580 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1710841341
transform 1 0 2484 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1710841341
transform 1 0 2468 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1710841341
transform 1 0 2452 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1710841341
transform 1 0 2436 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1710841341
transform 1 0 2420 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1710841341
transform 1 0 2420 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1710841341
transform 1 0 2068 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1710841341
transform 1 0 2052 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1710841341
transform 1 0 2004 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1710841341
transform 1 0 1932 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1710841341
transform 1 0 1844 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1710841341
transform 1 0 1636 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1710841341
transform 1 0 1628 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1710841341
transform 1 0 1628 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1710841341
transform 1 0 1444 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1710841341
transform 1 0 1108 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1710841341
transform 1 0 1068 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1710841341
transform 1 0 996 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1710841341
transform 1 0 980 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1710841341
transform 1 0 828 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1710841341
transform 1 0 740 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1710841341
transform 1 0 668 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1710841341
transform 1 0 660 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1710841341
transform 1 0 652 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1710841341
transform 1 0 540 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1710841341
transform 1 0 484 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1710841341
transform 1 0 412 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1710841341
transform 1 0 380 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1710841341
transform 1 0 340 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1710841341
transform 1 0 292 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1710841341
transform 1 0 252 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1710841341
transform 1 0 172 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1710841341
transform 1 0 172 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1710841341
transform 1 0 132 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1710841341
transform 1 0 124 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1710841341
transform 1 0 100 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1710841341
transform 1 0 84 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1710841341
transform 1 0 76 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1710841341
transform 1 0 76 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1710841341
transform 1 0 2660 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1710841341
transform 1 0 2660 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1710841341
transform 1 0 2612 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1710841341
transform 1 0 2588 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1710841341
transform 1 0 2548 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1710841341
transform 1 0 2524 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1710841341
transform 1 0 2500 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1710841341
transform 1 0 2468 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1710841341
transform 1 0 2428 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1710841341
transform 1 0 2388 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1710841341
transform 1 0 2036 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1710841341
transform 1 0 1940 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1710841341
transform 1 0 1916 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1710841341
transform 1 0 1900 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1710841341
transform 1 0 1804 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1710841341
transform 1 0 1788 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1710841341
transform 1 0 1772 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1710841341
transform 1 0 1596 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1710841341
transform 1 0 1196 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1710841341
transform 1 0 1060 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1710841341
transform 1 0 1044 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1710841341
transform 1 0 780 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1710841341
transform 1 0 764 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1710841341
transform 1 0 636 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1710841341
transform 1 0 636 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1710841341
transform 1 0 540 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1710841341
transform 1 0 540 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1710841341
transform 1 0 524 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1710841341
transform 1 0 516 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1710841341
transform 1 0 476 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1710841341
transform 1 0 476 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1710841341
transform 1 0 468 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1710841341
transform 1 0 460 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1710841341
transform 1 0 404 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1710841341
transform 1 0 404 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1710841341
transform 1 0 404 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1710841341
transform 1 0 380 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1710841341
transform 1 0 380 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1710841341
transform 1 0 252 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1710841341
transform 1 0 220 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1710841341
transform 1 0 212 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1710841341
transform 1 0 204 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1710841341
transform 1 0 204 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1710841341
transform 1 0 196 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1710841341
transform 1 0 1300 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1710841341
transform 1 0 1172 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1710841341
transform 1 0 988 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1710841341
transform 1 0 980 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1710841341
transform 1 0 900 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1710841341
transform 1 0 476 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1710841341
transform 1 0 476 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1710841341
transform 1 0 436 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1710841341
transform 1 0 228 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1710841341
transform 1 0 172 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1710841341
transform 1 0 124 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1710841341
transform 1 0 116 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1710841341
transform 1 0 116 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1710841341
transform 1 0 668 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1710841341
transform 1 0 572 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1710841341
transform 1 0 564 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1710841341
transform 1 0 516 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1710841341
transform 1 0 468 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1710841341
transform 1 0 452 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1710841341
transform 1 0 420 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1710841341
transform 1 0 404 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1710841341
transform 1 0 364 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1710841341
transform 1 0 308 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1710841341
transform 1 0 268 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1710841341
transform 1 0 372 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1710841341
transform 1 0 252 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1710841341
transform 1 0 1764 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1710841341
transform 1 0 1732 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1710841341
transform 1 0 1828 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1710841341
transform 1 0 1796 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1710841341
transform 1 0 2468 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1710841341
transform 1 0 2420 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1710841341
transform 1 0 996 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1710841341
transform 1 0 932 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1710841341
transform 1 0 828 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1710841341
transform 1 0 2188 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1710841341
transform 1 0 2164 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1710841341
transform 1 0 2124 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1710841341
transform 1 0 2124 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1710841341
transform 1 0 1668 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1710841341
transform 1 0 1636 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1710841341
transform 1 0 1572 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1710841341
transform 1 0 332 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1710841341
transform 1 0 300 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1710841341
transform 1 0 2284 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1710841341
transform 1 0 2220 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1710841341
transform 1 0 2076 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1710841341
transform 1 0 1964 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1710841341
transform 1 0 1844 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1710841341
transform 1 0 1844 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1710841341
transform 1 0 1532 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1710841341
transform 1 0 1532 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1710841341
transform 1 0 1428 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1710841341
transform 1 0 2092 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1710841341
transform 1 0 1988 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1710841341
transform 1 0 1892 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1710841341
transform 1 0 1884 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1710841341
transform 1 0 1548 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1710841341
transform 1 0 1428 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1710841341
transform 1 0 1428 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1710841341
transform 1 0 1428 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1710841341
transform 1 0 1316 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1710841341
transform 1 0 1212 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1710841341
transform 1 0 1204 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1710841341
transform 1 0 1188 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1710841341
transform 1 0 1140 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1710841341
transform 1 0 868 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1710841341
transform 1 0 1660 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1710841341
transform 1 0 1652 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1710841341
transform 1 0 1476 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1710841341
transform 1 0 1252 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1710841341
transform 1 0 996 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1710841341
transform 1 0 1220 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1710841341
transform 1 0 1164 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1710841341
transform 1 0 964 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1710841341
transform 1 0 916 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1710841341
transform 1 0 804 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1710841341
transform 1 0 724 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1710841341
transform 1 0 724 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1710841341
transform 1 0 716 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1710841341
transform 1 0 660 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1710841341
transform 1 0 588 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1710841341
transform 1 0 564 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1710841341
transform 1 0 1972 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1710841341
transform 1 0 1924 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1710841341
transform 1 0 1924 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1710841341
transform 1 0 1788 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1710841341
transform 1 0 1788 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1710841341
transform 1 0 1572 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1710841341
transform 1 0 1524 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1710841341
transform 1 0 1524 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1710841341
transform 1 0 1500 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1710841341
transform 1 0 1428 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1710841341
transform 1 0 1420 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1710841341
transform 1 0 1308 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1710841341
transform 1 0 1260 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1710841341
transform 1 0 1244 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1710841341
transform 1 0 1228 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1710841341
transform 1 0 1228 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1710841341
transform 1 0 1172 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1710841341
transform 1 0 1036 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1710841341
transform 1 0 1036 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1710841341
transform 1 0 660 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1710841341
transform 1 0 1964 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1710841341
transform 1 0 1956 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1710841341
transform 1 0 1876 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1710841341
transform 1 0 1788 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1710841341
transform 1 0 1788 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1710841341
transform 1 0 1756 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1710841341
transform 1 0 1660 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1710841341
transform 1 0 1612 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1710841341
transform 1 0 1556 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1710841341
transform 1 0 724 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1710841341
transform 1 0 1836 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1710841341
transform 1 0 1772 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1710841341
transform 1 0 1772 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1710841341
transform 1 0 1644 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1710841341
transform 1 0 1548 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1710841341
transform 1 0 1428 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1710841341
transform 1 0 1428 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1710841341
transform 1 0 916 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1710841341
transform 1 0 908 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1710841341
transform 1 0 852 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1710841341
transform 1 0 852 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1710841341
transform 1 0 828 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1710841341
transform 1 0 820 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1710841341
transform 1 0 820 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1710841341
transform 1 0 748 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1710841341
transform 1 0 748 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1710841341
transform 1 0 724 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1710841341
transform 1 0 692 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1710841341
transform 1 0 676 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1710841341
transform 1 0 676 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1710841341
transform 1 0 292 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1710841341
transform 1 0 212 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1710841341
transform 1 0 220 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1710841341
transform 1 0 148 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1710841341
transform 1 0 276 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1710841341
transform 1 0 188 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1710841341
transform 1 0 196 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1710841341
transform 1 0 156 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1710841341
transform 1 0 180 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1710841341
transform 1 0 148 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1710841341
transform 1 0 220 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1710841341
transform 1 0 140 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1710841341
transform 1 0 220 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1710841341
transform 1 0 132 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1710841341
transform 1 0 612 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1710841341
transform 1 0 260 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1710841341
transform 1 0 596 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1710841341
transform 1 0 500 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1710841341
transform 1 0 1436 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1710841341
transform 1 0 1428 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1710841341
transform 1 0 1364 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1710841341
transform 1 0 652 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1710841341
transform 1 0 652 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1710841341
transform 1 0 532 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1710841341
transform 1 0 172 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1710841341
transform 1 0 132 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1710841341
transform 1 0 1756 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1710841341
transform 1 0 1676 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1710841341
transform 1 0 2660 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1710841341
transform 1 0 2636 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1710841341
transform 1 0 2676 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1710841341
transform 1 0 2636 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1710841341
transform 1 0 2668 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1710841341
transform 1 0 2636 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1710841341
transform 1 0 2612 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1710841341
transform 1 0 2556 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1710841341
transform 1 0 2612 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1710841341
transform 1 0 2564 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1710841341
transform 1 0 2484 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1710841341
transform 1 0 2444 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1710841341
transform 1 0 1868 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1710841341
transform 1 0 1796 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1710841341
transform 1 0 1196 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1710841341
transform 1 0 1116 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1710841341
transform 1 0 1044 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1710841341
transform 1 0 788 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1710841341
transform 1 0 380 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1710841341
transform 1 0 300 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1710841341
transform 1 0 316 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1710841341
transform 1 0 220 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1710841341
transform 1 0 524 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1710841341
transform 1 0 388 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1710841341
transform 1 0 388 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1710841341
transform 1 0 340 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1710841341
transform 1 0 732 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1710841341
transform 1 0 260 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1710841341
transform 1 0 2564 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1710841341
transform 1 0 2092 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1710841341
transform 1 0 2524 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1710841341
transform 1 0 2164 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1710841341
transform 1 0 2580 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1710841341
transform 1 0 2164 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1710841341
transform 1 0 556 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1710841341
transform 1 0 492 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1710841341
transform 1 0 380 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1710841341
transform 1 0 348 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1710841341
transform 1 0 2116 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1710841341
transform 1 0 2068 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1710841341
transform 1 0 212 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1710841341
transform 1 0 84 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1710841341
transform 1 0 1876 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1710841341
transform 1 0 1780 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1710841341
transform 1 0 1588 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1710841341
transform 1 0 1580 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1710841341
transform 1 0 1524 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1710841341
transform 1 0 1788 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1710841341
transform 1 0 1764 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1710841341
transform 1 0 1740 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1710841341
transform 1 0 1740 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1710841341
transform 1 0 1548 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1710841341
transform 1 0 1548 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1710841341
transform 1 0 1452 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1710841341
transform 1 0 1452 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1710841341
transform 1 0 1404 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1710841341
transform 1 0 1404 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1710841341
transform 1 0 1244 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1710841341
transform 1 0 1196 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1710841341
transform 1 0 1092 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1710841341
transform 1 0 1076 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1710841341
transform 1 0 156 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1710841341
transform 1 0 92 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1710841341
transform 1 0 164 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1710841341
transform 1 0 84 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1710841341
transform 1 0 1300 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1710841341
transform 1 0 1076 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1710841341
transform 1 0 964 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1710841341
transform 1 0 956 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1710841341
transform 1 0 2636 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1710841341
transform 1 0 2540 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1710841341
transform 1 0 1908 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1710841341
transform 1 0 1860 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1710841341
transform 1 0 1572 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1710841341
transform 1 0 1444 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1710841341
transform 1 0 1444 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1710841341
transform 1 0 1380 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1710841341
transform 1 0 1340 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1710841341
transform 1 0 1044 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1710841341
transform 1 0 948 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1710841341
transform 1 0 2364 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1710841341
transform 1 0 2284 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1710841341
transform 1 0 2452 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1710841341
transform 1 0 2340 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1710841341
transform 1 0 2212 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1710841341
transform 1 0 2116 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1710841341
transform 1 0 2556 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1710841341
transform 1 0 2516 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1710841341
transform 1 0 1860 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1710841341
transform 1 0 1828 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1710841341
transform 1 0 1772 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1710841341
transform 1 0 1708 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1710841341
transform 1 0 1644 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1710841341
transform 1 0 1644 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1710841341
transform 1 0 1172 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1710841341
transform 1 0 556 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1710841341
transform 1 0 508 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1710841341
transform 1 0 1932 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1710841341
transform 1 0 1892 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1710841341
transform 1 0 1940 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1710841341
transform 1 0 1900 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1710841341
transform 1 0 1844 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1710841341
transform 1 0 1748 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1710841341
transform 1 0 1780 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1710841341
transform 1 0 1732 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1710841341
transform 1 0 1500 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1710841341
transform 1 0 1500 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1710841341
transform 1 0 1500 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1710841341
transform 1 0 1484 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1710841341
transform 1 0 1092 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1710841341
transform 1 0 1076 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1710841341
transform 1 0 1060 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1710841341
transform 1 0 1028 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1710841341
transform 1 0 956 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1710841341
transform 1 0 1844 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1710841341
transform 1 0 1804 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1710841341
transform 1 0 1804 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1710841341
transform 1 0 1668 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1710841341
transform 1 0 1892 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1710841341
transform 1 0 1852 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1710841341
transform 1 0 2436 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1710841341
transform 1 0 2268 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1710841341
transform 1 0 2268 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1710841341
transform 1 0 2244 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1710841341
transform 1 0 1996 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1710841341
transform 1 0 1900 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1710841341
transform 1 0 660 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1710841341
transform 1 0 628 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1710841341
transform 1 0 500 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1710841341
transform 1 0 444 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1710841341
transform 1 0 2268 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1710841341
transform 1 0 2140 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1710841341
transform 1 0 2388 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1710841341
transform 1 0 2364 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1710841341
transform 1 0 420 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1710841341
transform 1 0 356 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1710841341
transform 1 0 2316 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1710841341
transform 1 0 2268 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1710841341
transform 1 0 964 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1710841341
transform 1 0 940 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1710841341
transform 1 0 2060 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1710841341
transform 1 0 1988 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1710841341
transform 1 0 1700 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1710841341
transform 1 0 1684 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1710841341
transform 1 0 1628 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1710841341
transform 1 0 1628 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1710841341
transform 1 0 1556 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1710841341
transform 1 0 1500 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1710841341
transform 1 0 1324 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1710841341
transform 1 0 1324 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1710841341
transform 1 0 1260 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1710841341
transform 1 0 1196 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1710841341
transform 1 0 2332 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1710841341
transform 1 0 2188 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1710841341
transform 1 0 2068 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1710841341
transform 1 0 2004 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1710841341
transform 1 0 2636 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1710841341
transform 1 0 2612 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1710841341
transform 1 0 660 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1710841341
transform 1 0 444 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1710841341
transform 1 0 1932 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1710841341
transform 1 0 1900 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1710841341
transform 1 0 1324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1710841341
transform 1 0 1212 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1710841341
transform 1 0 1044 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1710841341
transform 1 0 988 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1710841341
transform 1 0 388 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1710841341
transform 1 0 364 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1710841341
transform 1 0 1204 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1710841341
transform 1 0 1116 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1710841341
transform 1 0 2236 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1710841341
transform 1 0 2188 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1710841341
transform 1 0 2188 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1710841341
transform 1 0 2188 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1710841341
transform 1 0 2156 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1710841341
transform 1 0 2036 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1710841341
transform 1 0 2020 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1710841341
transform 1 0 1916 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1710841341
transform 1 0 1884 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1710841341
transform 1 0 1484 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1710841341
transform 1 0 780 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1710841341
transform 1 0 540 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1710841341
transform 1 0 532 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1710841341
transform 1 0 500 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1710841341
transform 1 0 476 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1710841341
transform 1 0 460 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1710841341
transform 1 0 460 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1710841341
transform 1 0 412 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1710841341
transform 1 0 2396 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1710841341
transform 1 0 2316 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1710841341
transform 1 0 2476 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1710841341
transform 1 0 2404 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1710841341
transform 1 0 2404 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1710841341
transform 1 0 2404 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1710841341
transform 1 0 2388 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1710841341
transform 1 0 2364 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1710841341
transform 1 0 2316 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1710841341
transform 1 0 2140 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1710841341
transform 1 0 2132 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1710841341
transform 1 0 2116 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1710841341
transform 1 0 2116 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1710841341
transform 1 0 2108 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1710841341
transform 1 0 1596 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1710841341
transform 1 0 2116 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1710841341
transform 1 0 2028 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1710841341
transform 1 0 1908 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1710841341
transform 1 0 1828 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1710841341
transform 1 0 1780 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1710841341
transform 1 0 2380 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1710841341
transform 1 0 2300 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1710841341
transform 1 0 2300 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1710841341
transform 1 0 2268 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1710841341
transform 1 0 2268 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1710841341
transform 1 0 2236 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1710841341
transform 1 0 2236 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1710841341
transform 1 0 2188 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1710841341
transform 1 0 2148 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1710841341
transform 1 0 1940 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1710841341
transform 1 0 1740 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1710841341
transform 1 0 1580 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1710841341
transform 1 0 1580 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1710841341
transform 1 0 748 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1710841341
transform 1 0 748 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1710841341
transform 1 0 684 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1710841341
transform 1 0 660 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1710841341
transform 1 0 2180 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1710841341
transform 1 0 2012 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1710841341
transform 1 0 2012 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1710841341
transform 1 0 1964 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1710841341
transform 1 0 1908 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1710841341
transform 1 0 1892 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1710841341
transform 1 0 2012 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1710841341
transform 1 0 1924 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1710841341
transform 1 0 1860 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1710841341
transform 1 0 1740 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1710841341
transform 1 0 1556 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1710841341
transform 1 0 1516 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1710841341
transform 1 0 2156 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1710841341
transform 1 0 1956 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1710841341
transform 1 0 1956 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1710841341
transform 1 0 1484 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1710841341
transform 1 0 1476 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1710841341
transform 1 0 1412 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1710841341
transform 1 0 1356 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1710841341
transform 1 0 772 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1710841341
transform 1 0 604 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1710841341
transform 1 0 564 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1710841341
transform 1 0 532 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1710841341
transform 1 0 404 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1710841341
transform 1 0 2428 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1710841341
transform 1 0 2348 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1710841341
transform 1 0 2244 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1710841341
transform 1 0 2036 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1710841341
transform 1 0 2020 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1710841341
transform 1 0 1988 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1710841341
transform 1 0 1980 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1710841341
transform 1 0 1948 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1710841341
transform 1 0 1948 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1710841341
transform 1 0 1924 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1710841341
transform 1 0 1924 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1710841341
transform 1 0 1900 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1710841341
transform 1 0 1844 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1710841341
transform 1 0 1764 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1710841341
transform 1 0 1588 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1710841341
transform 1 0 1588 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1710841341
transform 1 0 1476 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1710841341
transform 1 0 1164 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1710841341
transform 1 0 1108 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1710841341
transform 1 0 2124 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1710841341
transform 1 0 2068 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1710841341
transform 1 0 2028 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1710841341
transform 1 0 2020 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1710841341
transform 1 0 1852 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1710841341
transform 1 0 1764 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1710841341
transform 1 0 1684 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1710841341
transform 1 0 2436 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1710841341
transform 1 0 2316 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1710841341
transform 1 0 1972 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1710841341
transform 1 0 1652 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1710841341
transform 1 0 1572 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1710841341
transform 1 0 1508 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1710841341
transform 1 0 1468 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1710841341
transform 1 0 1524 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1710841341
transform 1 0 1476 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1710841341
transform 1 0 2540 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1710841341
transform 1 0 2228 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1710841341
transform 1 0 2140 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1710841341
transform 1 0 2604 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1710841341
transform 1 0 2596 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1710841341
transform 1 0 2540 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1710841341
transform 1 0 2540 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1710841341
transform 1 0 1932 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1710841341
transform 1 0 1564 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1710841341
transform 1 0 1564 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1710841341
transform 1 0 1500 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1710841341
transform 1 0 1428 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1710841341
transform 1 0 1740 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1710841341
transform 1 0 1716 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1710841341
transform 1 0 1708 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1710841341
transform 1 0 1684 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1710841341
transform 1 0 1468 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1710841341
transform 1 0 1468 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1710841341
transform 1 0 1308 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1710841341
transform 1 0 1308 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1710841341
transform 1 0 1124 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1710841341
transform 1 0 1076 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1710841341
transform 1 0 1068 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1710841341
transform 1 0 332 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1710841341
transform 1 0 300 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1710841341
transform 1 0 220 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1710841341
transform 1 0 1228 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1710841341
transform 1 0 644 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1710841341
transform 1 0 588 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1710841341
transform 1 0 580 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1710841341
transform 1 0 508 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1710841341
transform 1 0 492 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1710841341
transform 1 0 492 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1710841341
transform 1 0 460 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1710841341
transform 1 0 772 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1710841341
transform 1 0 692 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1710841341
transform 1 0 1652 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1710841341
transform 1 0 1492 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1710841341
transform 1 0 1812 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1710841341
transform 1 0 1772 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1710841341
transform 1 0 1276 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1710841341
transform 1 0 1212 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1710841341
transform 1 0 2340 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1710841341
transform 1 0 2244 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1710841341
transform 1 0 2348 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1710841341
transform 1 0 2316 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1710841341
transform 1 0 1980 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1710841341
transform 1 0 1860 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1710841341
transform 1 0 2284 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1710841341
transform 1 0 2172 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1710841341
transform 1 0 468 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1710841341
transform 1 0 364 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1710841341
transform 1 0 1372 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1710841341
transform 1 0 1340 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1710841341
transform 1 0 1292 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1710841341
transform 1 0 1284 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1710841341
transform 1 0 1132 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1710841341
transform 1 0 196 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1710841341
transform 1 0 132 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1710841341
transform 1 0 188 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1710841341
transform 1 0 100 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1710841341
transform 1 0 148 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1710841341
transform 1 0 100 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1710841341
transform 1 0 1172 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1710841341
transform 1 0 1116 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1710841341
transform 1 0 996 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1710841341
transform 1 0 324 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1710841341
transform 1 0 252 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1710841341
transform 1 0 252 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1710841341
transform 1 0 204 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1710841341
transform 1 0 2332 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1710841341
transform 1 0 2316 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1710841341
transform 1 0 2292 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1710841341
transform 1 0 2220 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1710841341
transform 1 0 2220 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1710841341
transform 1 0 2180 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1710841341
transform 1 0 2180 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1710841341
transform 1 0 1956 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1710841341
transform 1 0 1676 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1710841341
transform 1 0 2620 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1710841341
transform 1 0 2532 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1710841341
transform 1 0 2196 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1710841341
transform 1 0 1988 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1710841341
transform 1 0 1988 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1710841341
transform 1 0 1708 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1710841341
transform 1 0 1596 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1710841341
transform 1 0 2228 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1710841341
transform 1 0 2140 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1710841341
transform 1 0 2132 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1710841341
transform 1 0 2108 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1710841341
transform 1 0 2084 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1710841341
transform 1 0 1988 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1710841341
transform 1 0 1988 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1710841341
transform 1 0 1868 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1710841341
transform 1 0 1716 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1710841341
transform 1 0 1436 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1710841341
transform 1 0 1412 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1710841341
transform 1 0 228 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1710841341
transform 1 0 148 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1710841341
transform 1 0 284 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1710841341
transform 1 0 172 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1710841341
transform 1 0 1612 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1710841341
transform 1 0 1596 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1710841341
transform 1 0 1476 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1710841341
transform 1 0 1364 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1710841341
transform 1 0 2268 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1710841341
transform 1 0 2220 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1710841341
transform 1 0 2292 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1710841341
transform 1 0 2260 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1710841341
transform 1 0 1132 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1710841341
transform 1 0 940 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1710841341
transform 1 0 764 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1710841341
transform 1 0 556 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1710841341
transform 1 0 396 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1710841341
transform 1 0 324 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1710841341
transform 1 0 2540 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1710841341
transform 1 0 2308 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1710841341
transform 1 0 2228 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1710841341
transform 1 0 2356 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1710841341
transform 1 0 2324 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1710841341
transform 1 0 1644 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1710841341
transform 1 0 1588 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1710841341
transform 1 0 1620 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1710841341
transform 1 0 1452 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1710841341
transform 1 0 1316 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1710841341
transform 1 0 484 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1710841341
transform 1 0 428 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1710841341
transform 1 0 428 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1710841341
transform 1 0 428 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1710841341
transform 1 0 396 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1710841341
transform 1 0 716 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1710841341
transform 1 0 644 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1710841341
transform 1 0 596 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1710841341
transform 1 0 556 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1710841341
transform 1 0 2516 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1710841341
transform 1 0 2412 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1710841341
transform 1 0 1940 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1710841341
transform 1 0 2244 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1710841341
transform 1 0 2148 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1710841341
transform 1 0 2180 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1710841341
transform 1 0 2132 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1710841341
transform 1 0 2492 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1710841341
transform 1 0 2404 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1710841341
transform 1 0 1244 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1710841341
transform 1 0 1196 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1710841341
transform 1 0 2356 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1710841341
transform 1 0 2260 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1710841341
transform 1 0 2388 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1710841341
transform 1 0 2348 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1710841341
transform 1 0 1836 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1710841341
transform 1 0 1740 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1710841341
transform 1 0 2252 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1710841341
transform 1 0 2220 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1710841341
transform 1 0 2204 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1710841341
transform 1 0 1756 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1710841341
transform 1 0 1820 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1710841341
transform 1 0 1788 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1710841341
transform 1 0 2148 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1710841341
transform 1 0 2124 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1710841341
transform 1 0 2100 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1710841341
transform 1 0 2092 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1710841341
transform 1 0 2036 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1710841341
transform 1 0 1804 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1710841341
transform 1 0 1772 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1710841341
transform 1 0 1772 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1710841341
transform 1 0 1068 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1710841341
transform 1 0 1012 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1710841341
transform 1 0 2132 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1710841341
transform 1 0 2076 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1710841341
transform 1 0 2076 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1710841341
transform 1 0 1412 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1710841341
transform 1 0 1020 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1710841341
transform 1 0 2228 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1710841341
transform 1 0 1988 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1710841341
transform 1 0 1988 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1710841341
transform 1 0 1540 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1710841341
transform 1 0 1540 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1710841341
transform 1 0 1444 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1710841341
transform 1 0 868 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1710841341
transform 1 0 1684 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1710841341
transform 1 0 1604 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1710841341
transform 1 0 2348 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1710841341
transform 1 0 2236 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1710841341
transform 1 0 2508 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1710841341
transform 1 0 2404 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1710841341
transform 1 0 2268 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1710841341
transform 1 0 1692 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1710841341
transform 1 0 1420 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1710841341
transform 1 0 1420 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1710841341
transform 1 0 1420 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1710841341
transform 1 0 1332 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1710841341
transform 1 0 956 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1710841341
transform 1 0 852 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1710841341
transform 1 0 628 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1710841341
transform 1 0 524 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1710841341
transform 1 0 284 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1710841341
transform 1 0 196 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1710841341
transform 1 0 292 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1710841341
transform 1 0 164 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1710841341
transform 1 0 1956 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1710841341
transform 1 0 1820 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1710841341
transform 1 0 1636 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1710841341
transform 1 0 1636 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1710841341
transform 1 0 1468 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1710841341
transform 1 0 660 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1710841341
transform 1 0 548 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1710841341
transform 1 0 484 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1710841341
transform 1 0 2484 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1710841341
transform 1 0 2452 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1710841341
transform 1 0 2180 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1710841341
transform 1 0 2020 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1710841341
transform 1 0 1828 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1710841341
transform 1 0 1796 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1710841341
transform 1 0 1780 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1710841341
transform 1 0 1620 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1710841341
transform 1 0 1580 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1710841341
transform 1 0 1980 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1710841341
transform 1 0 1908 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1710841341
transform 1 0 2420 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1710841341
transform 1 0 2108 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1710841341
transform 1 0 2388 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1710841341
transform 1 0 1436 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1710841341
transform 1 0 1380 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1710841341
transform 1 0 1212 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1710841341
transform 1 0 2028 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1710841341
transform 1 0 1988 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1710841341
transform 1 0 2180 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1710841341
transform 1 0 2100 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1710841341
transform 1 0 1212 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1710841341
transform 1 0 1020 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1710841341
transform 1 0 228 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1710841341
transform 1 0 116 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1710841341
transform 1 0 1052 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1710841341
transform 1 0 876 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1710841341
transform 1 0 628 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1710841341
transform 1 0 500 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1710841341
transform 1 0 484 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1710841341
transform 1 0 380 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1710841341
transform 1 0 268 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1710841341
transform 1 0 380 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1710841341
transform 1 0 324 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1710841341
transform 1 0 284 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1710841341
transform 1 0 140 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1710841341
transform 1 0 116 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1710841341
transform 1 0 452 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1710841341
transform 1 0 84 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1710841341
transform 1 0 1996 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1710841341
transform 1 0 1996 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1710841341
transform 1 0 1924 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1710841341
transform 1 0 1900 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1710841341
transform 1 0 860 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1710841341
transform 1 0 860 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1710841341
transform 1 0 580 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1710841341
transform 1 0 476 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1710841341
transform 1 0 476 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1710841341
transform 1 0 276 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1710841341
transform 1 0 260 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1710841341
transform 1 0 564 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1710841341
transform 1 0 348 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1710841341
transform 1 0 284 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1710841341
transform 1 0 236 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1710841341
transform 1 0 684 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1710841341
transform 1 0 604 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1710841341
transform 1 0 324 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1710841341
transform 1 0 140 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1710841341
transform 1 0 84 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1710841341
transform 1 0 228 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1710841341
transform 1 0 116 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1710841341
transform 1 0 308 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1710841341
transform 1 0 244 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1710841341
transform 1 0 1156 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1710841341
transform 1 0 836 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1710841341
transform 1 0 836 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1710841341
transform 1 0 364 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1710841341
transform 1 0 364 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1710841341
transform 1 0 300 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1710841341
transform 1 0 284 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1710841341
transform 1 0 116 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1710841341
transform 1 0 100 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1710841341
transform 1 0 908 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1710841341
transform 1 0 268 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1710841341
transform 1 0 204 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1710841341
transform 1 0 116 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1710841341
transform 1 0 92 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1710841341
transform 1 0 212 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1710841341
transform 1 0 100 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1710841341
transform 1 0 276 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1710841341
transform 1 0 212 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1710841341
transform 1 0 332 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1710841341
transform 1 0 268 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1710841341
transform 1 0 268 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1710841341
transform 1 0 188 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1710841341
transform 1 0 156 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1710841341
transform 1 0 860 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1710841341
transform 1 0 556 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1710841341
transform 1 0 532 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1710841341
transform 1 0 444 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1710841341
transform 1 0 1356 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1710841341
transform 1 0 1308 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1710841341
transform 1 0 1196 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1710841341
transform 1 0 1092 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1710841341
transform 1 0 1092 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1710841341
transform 1 0 500 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1710841341
transform 1 0 932 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1710841341
transform 1 0 460 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1710841341
transform 1 0 428 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1710841341
transform 1 0 428 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1710841341
transform 1 0 388 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1710841341
transform 1 0 324 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1710841341
transform 1 0 316 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1710841341
transform 1 0 276 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1710841341
transform 1 0 180 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1710841341
transform 1 0 724 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1710841341
transform 1 0 620 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1710841341
transform 1 0 620 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1710841341
transform 1 0 404 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1710841341
transform 1 0 364 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1710841341
transform 1 0 436 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1710841341
transform 1 0 356 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1710841341
transform 1 0 540 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1710841341
transform 1 0 348 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1710841341
transform 1 0 412 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1710841341
transform 1 0 396 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1710841341
transform 1 0 1364 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1710841341
transform 1 0 1332 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1710841341
transform 1 0 2140 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1710841341
transform 1 0 1988 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1710841341
transform 1 0 1988 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1710841341
transform 1 0 1460 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1710841341
transform 1 0 1060 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1710841341
transform 1 0 572 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1710841341
transform 1 0 524 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1710841341
transform 1 0 524 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1710841341
transform 1 0 524 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1710841341
transform 1 0 452 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1710841341
transform 1 0 724 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1710841341
transform 1 0 644 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1710841341
transform 1 0 716 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1710841341
transform 1 0 652 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1710841341
transform 1 0 884 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1710841341
transform 1 0 692 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1710841341
transform 1 0 644 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1710841341
transform 1 0 628 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1710841341
transform 1 0 612 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1710841341
transform 1 0 596 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1710841341
transform 1 0 812 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1710841341
transform 1 0 772 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1710841341
transform 1 0 860 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1710841341
transform 1 0 788 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1710841341
transform 1 0 628 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1710841341
transform 1 0 620 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1710841341
transform 1 0 604 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1710841341
transform 1 0 508 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1710841341
transform 1 0 412 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1710841341
transform 1 0 468 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1710841341
transform 1 0 420 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1710841341
transform 1 0 628 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1710841341
transform 1 0 444 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1710841341
transform 1 0 1772 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1710841341
transform 1 0 1724 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1710841341
transform 1 0 1724 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1710841341
transform 1 0 892 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1710841341
transform 1 0 796 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1710841341
transform 1 0 788 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1710841341
transform 1 0 580 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1710841341
transform 1 0 564 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1710841341
transform 1 0 660 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1710841341
transform 1 0 548 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1710841341
transform 1 0 556 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1710841341
transform 1 0 516 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1710841341
transform 1 0 660 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1710841341
transform 1 0 556 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1710841341
transform 1 0 1220 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1710841341
transform 1 0 1092 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1710841341
transform 1 0 660 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1710841341
transform 1 0 636 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1710841341
transform 1 0 636 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1710841341
transform 1 0 636 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1710841341
transform 1 0 636 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1710841341
transform 1 0 612 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1710841341
transform 1 0 612 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1710841341
transform 1 0 596 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1710841341
transform 1 0 1100 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1710841341
transform 1 0 964 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1710841341
transform 1 0 964 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1710841341
transform 1 0 604 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1710841341
transform 1 0 596 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1710841341
transform 1 0 588 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1710841341
transform 1 0 572 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1710841341
transform 1 0 540 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1710841341
transform 1 0 556 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1710841341
transform 1 0 500 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1710841341
transform 1 0 636 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1710841341
transform 1 0 468 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1710841341
transform 1 0 484 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1710841341
transform 1 0 436 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1710841341
transform 1 0 516 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1710841341
transform 1 0 484 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1710841341
transform 1 0 388 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1710841341
transform 1 0 380 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1710841341
transform 1 0 628 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1710841341
transform 1 0 396 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1710841341
transform 1 0 588 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1710841341
transform 1 0 388 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1710841341
transform 1 0 716 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1710841341
transform 1 0 716 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1710841341
transform 1 0 660 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1710841341
transform 1 0 580 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1710841341
transform 1 0 1700 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1710841341
transform 1 0 1572 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1710841341
transform 1 0 788 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1710841341
transform 1 0 692 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1710841341
transform 1 0 812 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1710841341
transform 1 0 700 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1710841341
transform 1 0 708 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1710841341
transform 1 0 668 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1710841341
transform 1 0 1804 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1710841341
transform 1 0 1652 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1710841341
transform 1 0 1596 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1710841341
transform 1 0 1588 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1710841341
transform 1 0 1572 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1710841341
transform 1 0 1572 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1710841341
transform 1 0 1476 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1710841341
transform 1 0 1468 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1710841341
transform 1 0 1396 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1710841341
transform 1 0 1396 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1710841341
transform 1 0 1132 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1710841341
transform 1 0 1124 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1710841341
transform 1 0 1108 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1710841341
transform 1 0 1076 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1710841341
transform 1 0 1052 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1710841341
transform 1 0 804 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1710841341
transform 1 0 804 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1710841341
transform 1 0 700 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1710841341
transform 1 0 820 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1710841341
transform 1 0 748 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1710841341
transform 1 0 868 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1710841341
transform 1 0 748 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1710841341
transform 1 0 1068 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1710841341
transform 1 0 956 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1710841341
transform 1 0 956 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1710841341
transform 1 0 916 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1710841341
transform 1 0 852 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1710841341
transform 1 0 1004 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1710841341
transform 1 0 884 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1710841341
transform 1 0 868 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1710841341
transform 1 0 788 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1710841341
transform 1 0 1284 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1710841341
transform 1 0 1172 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1710841341
transform 1 0 1116 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1710841341
transform 1 0 1116 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1710841341
transform 1 0 1092 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1710841341
transform 1 0 1076 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1710841341
transform 1 0 1076 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1710841341
transform 1 0 1012 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1710841341
transform 1 0 892 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1710841341
transform 1 0 884 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1710841341
transform 1 0 844 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1710841341
transform 1 0 844 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1710841341
transform 1 0 964 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1710841341
transform 1 0 788 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1710841341
transform 1 0 1852 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1710841341
transform 1 0 1796 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1710841341
transform 1 0 1780 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1710841341
transform 1 0 1364 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1710841341
transform 1 0 1308 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1710841341
transform 1 0 964 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1710841341
transform 1 0 964 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1710841341
transform 1 0 932 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1710841341
transform 1 0 956 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1710841341
transform 1 0 932 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1710841341
transform 1 0 1876 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1710841341
transform 1 0 1852 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1710841341
transform 1 0 1844 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1710841341
transform 1 0 1100 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1710841341
transform 1 0 1100 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1710841341
transform 1 0 1044 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1710841341
transform 1 0 1908 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1710841341
transform 1 0 1876 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1710841341
transform 1 0 1156 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1710841341
transform 1 0 1132 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1710841341
transform 1 0 1132 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1710841341
transform 1 0 1084 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1710841341
transform 1 0 1068 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1710841341
transform 1 0 1036 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1710841341
transform 1 0 1036 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1710841341
transform 1 0 1012 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1710841341
transform 1 0 1004 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1710841341
transform 1 0 908 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1710841341
transform 1 0 828 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1710841341
transform 1 0 740 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1710841341
transform 1 0 724 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1710841341
transform 1 0 684 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1710841341
transform 1 0 1244 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1710841341
transform 1 0 1044 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1710841341
transform 1 0 884 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1710841341
transform 1 0 868 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1710841341
transform 1 0 1148 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1710841341
transform 1 0 1060 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1710841341
transform 1 0 828 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1710841341
transform 1 0 1044 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1710841341
transform 1 0 1044 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1710841341
transform 1 0 1028 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1710841341
transform 1 0 844 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1710841341
transform 1 0 844 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1710841341
transform 1 0 532 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1710841341
transform 1 0 1036 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1710841341
transform 1 0 1004 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1710841341
transform 1 0 1388 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1710841341
transform 1 0 1380 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1710841341
transform 1 0 1236 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1710841341
transform 1 0 1204 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1710841341
transform 1 0 1140 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1710841341
transform 1 0 1132 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1710841341
transform 1 0 1084 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1710841341
transform 1 0 1076 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1710841341
transform 1 0 820 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1710841341
transform 1 0 780 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1710841341
transform 1 0 1292 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1710841341
transform 1 0 1220 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1710841341
transform 1 0 1188 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1710841341
transform 1 0 1084 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1710841341
transform 1 0 1764 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1710841341
transform 1 0 1732 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1710841341
transform 1 0 1652 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1710841341
transform 1 0 1652 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1710841341
transform 1 0 1196 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1710841341
transform 1 0 1188 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1710841341
transform 1 0 1156 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1710841341
transform 1 0 1196 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1710841341
transform 1 0 1140 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1710841341
transform 1 0 1660 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1710841341
transform 1 0 1636 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1710841341
transform 1 0 1028 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1710841341
transform 1 0 1012 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1710841341
transform 1 0 1012 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1710841341
transform 1 0 956 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1710841341
transform 1 0 1668 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1710841341
transform 1 0 1580 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1710841341
transform 1 0 1196 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1710841341
transform 1 0 1156 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1710841341
transform 1 0 1140 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1710841341
transform 1 0 1100 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1710841341
transform 1 0 1092 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1710841341
transform 1 0 1092 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1710841341
transform 1 0 1084 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1710841341
transform 1 0 1052 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1710841341
transform 1 0 1164 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1710841341
transform 1 0 1132 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1710841341
transform 1 0 1100 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1710841341
transform 1 0 1100 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1710841341
transform 1 0 1020 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1710841341
transform 1 0 1020 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1710841341
transform 1 0 948 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1710841341
transform 1 0 940 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1710841341
transform 1 0 364 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1710841341
transform 1 0 300 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1710841341
transform 1 0 540 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1710841341
transform 1 0 324 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1710841341
transform 1 0 604 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1710841341
transform 1 0 524 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1710841341
transform 1 0 492 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1710841341
transform 1 0 444 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1710841341
transform 1 0 404 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1710841341
transform 1 0 620 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1710841341
transform 1 0 452 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1710841341
transform 1 0 348 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1710841341
transform 1 0 284 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1710841341
transform 1 0 420 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1710841341
transform 1 0 268 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1710841341
transform 1 0 588 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1710841341
transform 1 0 484 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1710841341
transform 1 0 1364 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1710841341
transform 1 0 1340 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1710841341
transform 1 0 1292 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1710841341
transform 1 0 1260 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1710841341
transform 1 0 1260 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1710841341
transform 1 0 1252 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1710841341
transform 1 0 1252 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1710841341
transform 1 0 1212 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1710841341
transform 1 0 1196 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1710841341
transform 1 0 804 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1710841341
transform 1 0 804 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1710841341
transform 1 0 572 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1710841341
transform 1 0 572 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1710841341
transform 1 0 444 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1710841341
transform 1 0 780 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1710841341
transform 1 0 588 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1710841341
transform 1 0 2004 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1710841341
transform 1 0 2004 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1710841341
transform 1 0 1948 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1710841341
transform 1 0 788 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1710841341
transform 1 0 860 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1710841341
transform 1 0 524 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1710841341
transform 1 0 452 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1710841341
transform 1 0 356 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1710841341
transform 1 0 612 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1710841341
transform 1 0 500 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1710841341
transform 1 0 740 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1710841341
transform 1 0 684 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1710841341
transform 1 0 1268 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1710841341
transform 1 0 1012 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1710841341
transform 1 0 996 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1710841341
transform 1 0 700 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1710841341
transform 1 0 748 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1710841341
transform 1 0 516 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1710841341
transform 1 0 828 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1710841341
transform 1 0 716 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1710841341
transform 1 0 692 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1710841341
transform 1 0 596 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1710841341
transform 1 0 540 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1710841341
transform 1 0 1508 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1710841341
transform 1 0 1340 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1710841341
transform 1 0 1340 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1710841341
transform 1 0 796 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1710841341
transform 1 0 780 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1710841341
transform 1 0 780 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1710841341
transform 1 0 732 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1710841341
transform 1 0 620 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1710841341
transform 1 0 668 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1710841341
transform 1 0 468 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1710841341
transform 1 0 372 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1710841341
transform 1 0 1892 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1710841341
transform 1 0 1468 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1710841341
transform 1 0 1364 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1710841341
transform 1 0 1364 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1710841341
transform 1 0 1356 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1710841341
transform 1 0 1292 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1710841341
transform 1 0 1292 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1710841341
transform 1 0 948 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1710841341
transform 1 0 492 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1710841341
transform 1 0 396 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1710841341
transform 1 0 556 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1710841341
transform 1 0 540 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1710841341
transform 1 0 1188 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1710841341
transform 1 0 1132 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1710841341
transform 1 0 1388 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1710841341
transform 1 0 1284 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1710841341
transform 1 0 1260 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1710841341
transform 1 0 1060 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1710841341
transform 1 0 996 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1710841341
transform 1 0 924 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1710841341
transform 1 0 852 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1710841341
transform 1 0 1724 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1710841341
transform 1 0 1204 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1710841341
transform 1 0 1204 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1710841341
transform 1 0 1084 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1710841341
transform 1 0 1012 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1710841341
transform 1 0 940 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1710841341
transform 1 0 868 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1710841341
transform 1 0 892 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1710841341
transform 1 0 828 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1710841341
transform 1 0 972 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1710841341
transform 1 0 900 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1710841341
transform 1 0 996 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1710841341
transform 1 0 940 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1710841341
transform 1 0 924 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1710841341
transform 1 0 876 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1710841341
transform 1 0 836 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1710841341
transform 1 0 1220 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1710841341
transform 1 0 1172 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1710841341
transform 1 0 1380 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1710841341
transform 1 0 1188 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1710841341
transform 1 0 1412 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1710841341
transform 1 0 1300 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1710841341
transform 1 0 1268 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1710841341
transform 1 0 1436 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1710841341
transform 1 0 1436 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1710841341
transform 1 0 1436 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1710841341
transform 1 0 1412 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1710841341
transform 1 0 1412 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1710841341
transform 1 0 1412 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1710841341
transform 1 0 1388 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1710841341
transform 1 0 1372 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1710841341
transform 1 0 1276 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1710841341
transform 1 0 1228 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1710841341
transform 1 0 1196 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1710841341
transform 1 0 1596 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1710841341
transform 1 0 1340 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1710841341
transform 1 0 1268 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1710841341
transform 1 0 1252 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1710841341
transform 1 0 1396 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1710841341
transform 1 0 1396 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1710841341
transform 1 0 1396 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1710841341
transform 1 0 1380 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1710841341
transform 1 0 1356 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1710841341
transform 1 0 1348 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1710841341
transform 1 0 1308 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1710841341
transform 1 0 1260 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1710841341
transform 1 0 1276 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1710841341
transform 1 0 1228 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1710841341
transform 1 0 1268 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1710841341
transform 1 0 980 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1710841341
transform 1 0 1324 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1710841341
transform 1 0 1220 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1710841341
transform 1 0 1244 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1710841341
transform 1 0 1164 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1710841341
transform 1 0 1348 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1710841341
transform 1 0 1260 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1710841341
transform 1 0 1500 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1710841341
transform 1 0 1484 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1710841341
transform 1 0 1492 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1710841341
transform 1 0 1460 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1710841341
transform 1 0 1452 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1710841341
transform 1 0 1412 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1710841341
transform 1 0 1412 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1710841341
transform 1 0 1396 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1710841341
transform 1 0 1388 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1710841341
transform 1 0 1564 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1710841341
transform 1 0 1564 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1710841341
transform 1 0 1524 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1710841341
transform 1 0 1460 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1710841341
transform 1 0 1492 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1710841341
transform 1 0 1468 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1710841341
transform 1 0 2052 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1710841341
transform 1 0 1444 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1710841341
transform 1 0 1420 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1710841341
transform 1 0 1420 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1710841341
transform 1 0 988 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1710841341
transform 1 0 972 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1710841341
transform 1 0 1388 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1710841341
transform 1 0 940 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1710841341
transform 1 0 1500 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1710841341
transform 1 0 1436 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1710841341
transform 1 0 1444 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1710841341
transform 1 0 1404 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1710841341
transform 1 0 1524 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1710841341
transform 1 0 1476 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1710841341
transform 1 0 1540 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1710841341
transform 1 0 1508 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1710841341
transform 1 0 1548 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1710841341
transform 1 0 1484 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1710841341
transform 1 0 1484 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1710841341
transform 1 0 1404 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1710841341
transform 1 0 1588 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1710841341
transform 1 0 1556 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1710841341
transform 1 0 2100 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1710841341
transform 1 0 2020 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1710841341
transform 1 0 2012 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1710841341
transform 1 0 1660 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1710841341
transform 1 0 1628 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1710841341
transform 1 0 1668 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1710841341
transform 1 0 1596 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1710841341
transform 1 0 1692 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1710841341
transform 1 0 1636 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1710841341
transform 1 0 1652 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1710841341
transform 1 0 1612 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1710841341
transform 1 0 1588 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1710841341
transform 1 0 1556 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1710841341
transform 1 0 1716 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1710841341
transform 1 0 1668 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1710841341
transform 1 0 2012 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1710841341
transform 1 0 1764 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1710841341
transform 1 0 1660 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1710841341
transform 1 0 1572 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1710841341
transform 1 0 1596 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1710841341
transform 1 0 1452 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1710841341
transform 1 0 1716 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1710841341
transform 1 0 1684 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1710841341
transform 1 0 1684 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1710841341
transform 1 0 1660 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1710841341
transform 1 0 1948 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1710841341
transform 1 0 1908 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1710841341
transform 1 0 1900 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1710841341
transform 1 0 1820 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1710841341
transform 1 0 1860 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1710841341
transform 1 0 1772 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2584
timestamp 1710841341
transform 1 0 1756 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1710841341
transform 1 0 1700 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1710841341
transform 1 0 1812 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1710841341
transform 1 0 1740 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1710841341
transform 1 0 1908 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1710841341
transform 1 0 1876 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1710841341
transform 1 0 1948 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1710841341
transform 1 0 1924 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1710841341
transform 1 0 1804 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1710841341
transform 1 0 1772 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1710841341
transform 1 0 1876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1710841341
transform 1 0 1828 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1710841341
transform 1 0 1788 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1710841341
transform 1 0 1516 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1710841341
transform 1 0 1844 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2599
timestamp 1710841341
transform 1 0 1804 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1710841341
transform 1 0 1732 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1710841341
transform 1 0 1668 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1710841341
transform 1 0 2140 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1710841341
transform 1 0 1756 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1710841341
transform 1 0 1708 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1710841341
transform 1 0 1708 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1710841341
transform 1 0 1892 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1710841341
transform 1 0 1820 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1710841341
transform 1 0 1844 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1710841341
transform 1 0 1804 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1710841341
transform 1 0 1980 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1710841341
transform 1 0 1756 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1710841341
transform 1 0 1684 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1710841341
transform 1 0 1596 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1710841341
transform 1 0 1524 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1710841341
transform 1 0 2596 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1710841341
transform 1 0 2580 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1710841341
transform 1 0 2468 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1710841341
transform 1 0 2468 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1710841341
transform 1 0 2412 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1710841341
transform 1 0 2404 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1710841341
transform 1 0 2028 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1710841341
transform 1 0 2020 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1710841341
transform 1 0 1956 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1710841341
transform 1 0 1540 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1710841341
transform 1 0 2260 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1710841341
transform 1 0 2228 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1710841341
transform 1 0 2228 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1710841341
transform 1 0 2140 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1710841341
transform 1 0 2116 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1710841341
transform 1 0 2348 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1710841341
transform 1 0 2212 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1710841341
transform 1 0 2428 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1710841341
transform 1 0 2084 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1710841341
transform 1 0 2444 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1710841341
transform 1 0 2396 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1710841341
transform 1 0 2276 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1710841341
transform 1 0 2236 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1710841341
transform 1 0 2340 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1710841341
transform 1 0 2340 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1710841341
transform 1 0 2204 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1710841341
transform 1 0 2204 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1710841341
transform 1 0 1996 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1710841341
transform 1 0 1996 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1710841341
transform 1 0 1708 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1710841341
transform 1 0 2172 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1710841341
transform 1 0 2036 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1710841341
transform 1 0 2092 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1710841341
transform 1 0 1972 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1710841341
transform 1 0 2076 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1710841341
transform 1 0 2044 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1710841341
transform 1 0 1980 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1710841341
transform 1 0 1932 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1710841341
transform 1 0 1932 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1710841341
transform 1 0 1596 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1710841341
transform 1 0 2148 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1710841341
transform 1 0 2060 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1710841341
transform 1 0 2636 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1710841341
transform 1 0 2380 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1710841341
transform 1 0 2348 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1710841341
transform 1 0 1948 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1710841341
transform 1 0 1716 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1710841341
transform 1 0 1556 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1710841341
transform 1 0 2412 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1710841341
transform 1 0 2340 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1710841341
transform 1 0 2212 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1710841341
transform 1 0 2012 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1710841341
transform 1 0 2372 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1710841341
transform 1 0 2316 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1710841341
transform 1 0 2228 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1710841341
transform 1 0 2140 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1710841341
transform 1 0 2372 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1710841341
transform 1 0 2284 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1710841341
transform 1 0 2372 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1710841341
transform 1 0 2348 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1710841341
transform 1 0 2340 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1710841341
transform 1 0 2284 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1710841341
transform 1 0 2132 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1710841341
transform 1 0 2124 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1710841341
transform 1 0 2116 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1710841341
transform 1 0 1892 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1710841341
transform 1 0 1836 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1710841341
transform 1 0 1836 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1710841341
transform 1 0 2532 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1710841341
transform 1 0 2316 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1710841341
transform 1 0 2316 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1710841341
transform 1 0 2044 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1710841341
transform 1 0 2036 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1710841341
transform 1 0 2004 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1710841341
transform 1 0 2172 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1710841341
transform 1 0 2100 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1710841341
transform 1 0 2436 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1710841341
transform 1 0 2372 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1710841341
transform 1 0 2244 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1710841341
transform 1 0 2220 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1710841341
transform 1 0 2452 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1710841341
transform 1 0 2180 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1710841341
transform 1 0 2132 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1710841341
transform 1 0 2060 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1710841341
transform 1 0 2404 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1710841341
transform 1 0 2172 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1710841341
transform 1 0 2540 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1710841341
transform 1 0 2492 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1710841341
transform 1 0 2180 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1710841341
transform 1 0 2180 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1710841341
transform 1 0 1956 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1710841341
transform 1 0 2340 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1710841341
transform 1 0 2188 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1710841341
transform 1 0 2580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1710841341
transform 1 0 2484 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1710841341
transform 1 0 2380 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1710841341
transform 1 0 2468 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1710841341
transform 1 0 2436 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1710841341
transform 1 0 2556 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1710841341
transform 1 0 2516 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1710841341
transform 1 0 2444 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1710841341
transform 1 0 2156 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1710841341
transform 1 0 2156 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2718
timestamp 1710841341
transform 1 0 1964 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1710841341
transform 1 0 1964 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1710841341
transform 1 0 1900 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1710841341
transform 1 0 1884 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1710841341
transform 1 0 1868 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1710841341
transform 1 0 2556 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1710841341
transform 1 0 2460 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1710841341
transform 1 0 2172 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1710841341
transform 1 0 2084 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1710841341
transform 1 0 2660 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1710841341
transform 1 0 2548 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1710841341
transform 1 0 2660 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1710841341
transform 1 0 2636 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1710841341
transform 1 0 2604 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1710841341
transform 1 0 2660 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1710841341
transform 1 0 2620 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1710841341
transform 1 0 2636 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1710841341
transform 1 0 2580 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1710841341
transform 1 0 2596 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1710841341
transform 1 0 2556 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1710841341
transform 1 0 2540 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1710841341
transform 1 0 2428 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1710841341
transform 1 0 2508 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1710841341
transform 1 0 2204 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1710841341
transform 1 0 2508 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2743
timestamp 1710841341
transform 1 0 2388 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1710841341
transform 1 0 2388 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1710841341
transform 1 0 2260 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1710841341
transform 1 0 2260 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1710841341
transform 1 0 1828 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1710841341
transform 1 0 2612 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1710841341
transform 1 0 2484 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1710841341
transform 1 0 2468 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1710841341
transform 1 0 2564 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1710841341
transform 1 0 2124 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1710841341
transform 1 0 2580 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1710841341
transform 1 0 2524 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1710841341
transform 1 0 2660 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1710841341
transform 1 0 2628 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2757
timestamp 1710841341
transform 1 0 2636 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1710841341
transform 1 0 2636 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1710841341
transform 1 0 2628 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1710841341
transform 1 0 2620 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1710841341
transform 1 0 2612 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1710841341
transform 1 0 2564 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2763
timestamp 1710841341
transform 1 0 2532 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1710841341
transform 1 0 2532 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1710841341
transform 1 0 2092 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1710841341
transform 1 0 1892 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2767
timestamp 1710841341
transform 1 0 1652 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1710841341
transform 1 0 2604 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1710841341
transform 1 0 2556 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1710841341
transform 1 0 2116 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1710841341
transform 1 0 2044 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1710841341
transform 1 0 2644 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1710841341
transform 1 0 2540 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1710841341
transform 1 0 2596 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1710841341
transform 1 0 2524 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1710841341
transform 1 0 2540 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1710841341
transform 1 0 2460 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1710841341
transform 1 0 2580 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1710841341
transform 1 0 2556 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1710841341
transform 1 0 2540 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1710841341
transform 1 0 2244 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1710841341
transform 1 0 2532 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1710841341
transform 1 0 2468 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1710841341
transform 1 0 2372 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1710841341
transform 1 0 2300 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1710841341
transform 1 0 2148 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1710841341
transform 1 0 2420 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1710841341
transform 1 0 2404 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1710841341
transform 1 0 2364 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1710841341
transform 1 0 1908 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1710841341
transform 1 0 2540 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1710841341
transform 1 0 2276 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1710841341
transform 1 0 2068 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1710841341
transform 1 0 2020 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1710841341
transform 1 0 2068 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1710841341
transform 1 0 2052 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1710841341
transform 1 0 2204 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1710841341
transform 1 0 2164 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1710841341
transform 1 0 2316 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1710841341
transform 1 0 2284 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1710841341
transform 1 0 2092 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1710841341
transform 1 0 2060 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1710841341
transform 1 0 2236 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1710841341
transform 1 0 2084 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1710841341
transform 1 0 2060 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1710841341
transform 1 0 1748 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2807
timestamp 1710841341
transform 1 0 2532 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1710841341
transform 1 0 2452 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1710841341
transform 1 0 2436 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1710841341
transform 1 0 2188 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1710841341
transform 1 0 2468 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1710841341
transform 1 0 2396 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1710841341
transform 1 0 2348 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1710841341
transform 1 0 2332 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1710841341
transform 1 0 2228 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2816
timestamp 1710841341
transform 1 0 1772 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1710841341
transform 1 0 2356 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1710841341
transform 1 0 1956 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1710841341
transform 1 0 1716 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1710841341
transform 1 0 2212 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1710841341
transform 1 0 2188 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1710841341
transform 1 0 2260 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1710841341
transform 1 0 2204 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1710841341
transform 1 0 2484 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1710841341
transform 1 0 2324 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1710841341
transform 1 0 2468 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2827
timestamp 1710841341
transform 1 0 2044 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2828
timestamp 1710841341
transform 1 0 1940 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1710841341
transform 1 0 1892 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1710841341
transform 1 0 796 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1710841341
transform 1 0 772 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1710841341
transform 1 0 1036 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1710841341
transform 1 0 980 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1710841341
transform 1 0 740 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1710841341
transform 1 0 740 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2836
timestamp 1710841341
transform 1 0 708 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1710841341
transform 1 0 708 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1710841341
transform 1 0 620 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1710841341
transform 1 0 1916 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2840
timestamp 1710841341
transform 1 0 1748 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1710841341
transform 1 0 1740 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1710841341
transform 1 0 1540 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1710841341
transform 1 0 1412 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1710841341
transform 1 0 1988 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1710841341
transform 1 0 1844 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2846
timestamp 1710841341
transform 1 0 2644 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1710841341
transform 1 0 2524 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1710841341
transform 1 0 2484 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1710841341
transform 1 0 2372 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1710841341
transform 1 0 2508 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1710841341
transform 1 0 2444 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1710841341
transform 1 0 2380 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1710841341
transform 1 0 2228 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1710841341
transform 1 0 2172 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1710841341
transform 1 0 2164 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1710841341
transform 1 0 2068 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1710841341
transform 1 0 1900 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1710841341
transform 1 0 2100 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1710841341
transform 1 0 2028 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1710841341
transform 1 0 1972 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1710841341
transform 1 0 1804 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1710841341
transform 1 0 2580 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1710841341
transform 1 0 2500 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1710841341
transform 1 0 2548 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1710841341
transform 1 0 2060 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1710841341
transform 1 0 1964 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1710841341
transform 1 0 1892 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1710841341
transform 1 0 1100 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1710841341
transform 1 0 1052 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1710841341
transform 1 0 884 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2871
timestamp 1710841341
transform 1 0 1116 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1710841341
transform 1 0 1068 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2873
timestamp 1710841341
transform 1 0 964 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1710841341
transform 1 0 844 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1710841341
transform 1 0 844 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2876
timestamp 1710841341
transform 1 0 740 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1710841341
transform 1 0 2124 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1710841341
transform 1 0 1972 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1710841341
transform 1 0 2148 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1710841341
transform 1 0 1964 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1710841341
transform 1 0 2060 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1710841341
transform 1 0 1988 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1710841341
transform 1 0 1988 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1710841341
transform 1 0 1868 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1710841341
transform 1 0 1868 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1710841341
transform 1 0 1740 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1710841341
transform 1 0 2284 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1710841341
transform 1 0 1996 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1710841341
transform 1 0 1748 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1710841341
transform 1 0 1820 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1710841341
transform 1 0 1796 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1710841341
transform 1 0 1852 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1710841341
transform 1 0 1804 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1710841341
transform 1 0 1932 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1710841341
transform 1 0 1892 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1710841341
transform 1 0 1764 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1710841341
transform 1 0 1820 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1710841341
transform 1 0 1788 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1710841341
transform 1 0 948 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1710841341
transform 1 0 908 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1710841341
transform 1 0 732 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1710841341
transform 1 0 1164 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1710841341
transform 1 0 852 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1710841341
transform 1 0 836 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1710841341
transform 1 0 676 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1710841341
transform 1 0 2140 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1710841341
transform 1 0 2124 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1710841341
transform 1 0 1940 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1710841341
transform 1 0 1908 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1710841341
transform 1 0 1908 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1710841341
transform 1 0 1668 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1710841341
transform 1 0 1588 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1710841341
transform 1 0 2644 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1710841341
transform 1 0 2492 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1710841341
transform 1 0 2476 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1710841341
transform 1 0 2348 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1710841341
transform 1 0 2476 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1710841341
transform 1 0 2436 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1710841341
transform 1 0 2332 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1710841341
transform 1 0 2276 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1710841341
transform 1 0 2212 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1710841341
transform 1 0 2580 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1710841341
transform 1 0 2524 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1710841341
transform 1 0 2556 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1710841341
transform 1 0 2244 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1710841341
transform 1 0 2540 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1710841341
transform 1 0 2244 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1710841341
transform 1 0 1716 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1710841341
transform 1 0 1716 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1710841341
transform 1 0 1596 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1710841341
transform 1 0 1388 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1710841341
transform 1 0 1388 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1710841341
transform 1 0 1268 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1710841341
transform 1 0 2172 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1710841341
transform 1 0 1916 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1710841341
transform 1 0 2156 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1710841341
transform 1 0 1924 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1710841341
transform 1 0 804 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1710841341
transform 1 0 756 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1710841341
transform 1 0 884 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1710841341
transform 1 0 812 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1710841341
transform 1 0 700 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1710841341
transform 1 0 2188 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1710841341
transform 1 0 1988 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1710841341
transform 1 0 2612 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1710841341
transform 1 0 2540 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1710841341
transform 1 0 2508 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1710841341
transform 1 0 2372 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1710841341
transform 1 0 2532 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1710841341
transform 1 0 2468 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1710841341
transform 1 0 2508 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1710841341
transform 1 0 2436 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1710841341
transform 1 0 2452 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1710841341
transform 1 0 2244 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1710841341
transform 1 0 2116 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2956
timestamp 1710841341
transform 1 0 2444 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1710841341
transform 1 0 2188 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1710841341
transform 1 0 2548 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1710841341
transform 1 0 2532 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1710841341
transform 1 0 2492 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2961
timestamp 1710841341
transform 1 0 2492 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1710841341
transform 1 0 2508 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2963
timestamp 1710841341
transform 1 0 2508 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1710841341
transform 1 0 2484 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1710841341
transform 1 0 2308 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1710841341
transform 1 0 2132 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1710841341
transform 1 0 2124 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1710841341
transform 1 0 1956 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1710841341
transform 1 0 2172 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1710841341
transform 1 0 2092 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1710841341
transform 1 0 2652 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1710841341
transform 1 0 2580 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2973
timestamp 1710841341
transform 1 0 2532 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1710841341
transform 1 0 2460 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1710841341
transform 1 0 2628 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1710841341
transform 1 0 2596 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1710841341
transform 1 0 2340 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1710841341
transform 1 0 2252 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1710841341
transform 1 0 2268 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1710841341
transform 1 0 2148 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1710841341
transform 1 0 2060 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1710841341
transform 1 0 2252 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1710841341
transform 1 0 2180 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1710841341
transform 1 0 2340 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1710841341
transform 1 0 2180 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1710841341
transform 1 0 2436 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1710841341
transform 1 0 2324 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1710841341
transform 1 0 2124 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1710841341
transform 1 0 1692 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1710841341
transform 1 0 2308 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1710841341
transform 1 0 2236 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1710841341
transform 1 0 2284 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1710841341
transform 1 0 2244 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1710841341
transform 1 0 2204 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2995
timestamp 1710841341
transform 1 0 2164 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2996
timestamp 1710841341
transform 1 0 2268 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2997
timestamp 1710841341
transform 1 0 2180 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1710841341
transform 1 0 2092 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1710841341
transform 1 0 2004 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1710841341
transform 1 0 2012 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1710841341
transform 1 0 1964 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1710841341
transform 1 0 1972 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1710841341
transform 1 0 1876 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1710841341
transform 1 0 2068 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1710841341
transform 1 0 1932 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1710841341
transform 1 0 2036 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1710841341
transform 1 0 1972 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1710841341
transform 1 0 1964 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3009
timestamp 1710841341
transform 1 0 1844 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1710841341
transform 1 0 1844 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1710841341
transform 1 0 1820 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1710841341
transform 1 0 1780 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3013
timestamp 1710841341
transform 1 0 1564 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1710841341
transform 1 0 1564 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1710841341
transform 1 0 1260 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1710841341
transform 1 0 940 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1710841341
transform 1 0 940 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1710841341
transform 1 0 908 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3019
timestamp 1710841341
transform 1 0 1876 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1710841341
transform 1 0 1708 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1710841341
transform 1 0 1700 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1710841341
transform 1 0 1564 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1710841341
transform 1 0 2036 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3024
timestamp 1710841341
transform 1 0 1884 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1710841341
transform 1 0 2108 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1710841341
transform 1 0 2012 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1710841341
transform 1 0 1972 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1710841341
transform 1 0 1828 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1710841341
transform 1 0 1804 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1710841341
transform 1 0 1772 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3031
timestamp 1710841341
transform 1 0 932 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1710841341
transform 1 0 868 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1710841341
transform 1 0 1700 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1710841341
transform 1 0 1588 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1710841341
transform 1 0 1588 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1710841341
transform 1 0 1540 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1710841341
transform 1 0 1116 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1710841341
transform 1 0 932 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1710841341
transform 1 0 884 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3040
timestamp 1710841341
transform 1 0 876 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1710841341
transform 1 0 844 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1710841341
transform 1 0 804 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1710841341
transform 1 0 1780 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1710841341
transform 1 0 1684 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1710841341
transform 1 0 1596 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1710841341
transform 1 0 1524 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1710841341
transform 1 0 1524 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1710841341
transform 1 0 1484 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3049
timestamp 1710841341
transform 1 0 1460 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1710841341
transform 1 0 1460 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3051
timestamp 1710841341
transform 1 0 1428 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1710841341
transform 1 0 1428 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1710841341
transform 1 0 1396 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1710841341
transform 1 0 1388 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1710841341
transform 1 0 1388 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1710841341
transform 1 0 1196 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1710841341
transform 1 0 836 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1710841341
transform 1 0 1668 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1710841341
transform 1 0 1604 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1710841341
transform 1 0 1492 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1710841341
transform 1 0 1372 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1710841341
transform 1 0 1372 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1710841341
transform 1 0 1348 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1710841341
transform 1 0 972 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1710841341
transform 1 0 1748 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1710841341
transform 1 0 1668 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1710841341
transform 1 0 1612 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1710841341
transform 1 0 1596 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1710841341
transform 1 0 1540 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1710841341
transform 1 0 1532 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1710841341
transform 1 0 1508 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1710841341
transform 1 0 1356 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1710841341
transform 1 0 1356 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1710841341
transform 1 0 796 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1710841341
transform 1 0 1580 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1710841341
transform 1 0 1516 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1710841341
transform 1 0 1500 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1710841341
transform 1 0 1052 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1710841341
transform 1 0 1124 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1710841341
transform 1 0 1084 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1710841341
transform 1 0 1004 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1710841341
transform 1 0 980 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1710841341
transform 1 0 1356 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1710841341
transform 1 0 1276 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1710841341
transform 1 0 1444 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1710841341
transform 1 0 1324 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1710841341
transform 1 0 1388 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1710841341
transform 1 0 772 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1710841341
transform 1 0 1572 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1710841341
transform 1 0 1484 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1710841341
transform 1 0 1340 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1710841341
transform 1 0 1252 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1710841341
transform 1 0 1356 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1710841341
transform 1 0 1236 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1710841341
transform 1 0 1388 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1710841341
transform 1 0 1268 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1710841341
transform 1 0 1236 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1710841341
transform 1 0 1260 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1710841341
transform 1 0 1196 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1710841341
transform 1 0 1132 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1710841341
transform 1 0 1396 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1710841341
transform 1 0 1332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1710841341
transform 1 0 1348 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1710841341
transform 1 0 1028 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1710841341
transform 1 0 1476 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1710841341
transform 1 0 1412 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1710841341
transform 1 0 1492 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1710841341
transform 1 0 1436 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1710841341
transform 1 0 1228 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1710841341
transform 1 0 1092 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1710841341
transform 1 0 1236 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1710841341
transform 1 0 1132 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1710841341
transform 1 0 1004 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1710841341
transform 1 0 1372 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1710841341
transform 1 0 1300 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1710841341
transform 1 0 1332 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1710841341
transform 1 0 1284 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1710841341
transform 1 0 1212 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1710841341
transform 1 0 1052 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1710841341
transform 1 0 1412 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1710841341
transform 1 0 1340 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1710841341
transform 1 0 1316 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1710841341
transform 1 0 1140 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1710841341
transform 1 0 1172 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1710841341
transform 1 0 1124 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1710841341
transform 1 0 1100 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1710841341
transform 1 0 1068 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1710841341
transform 1 0 1044 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1710841341
transform 1 0 852 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1710841341
transform 1 0 852 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1710841341
transform 1 0 772 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1710841341
transform 1 0 772 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1710841341
transform 1 0 724 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1710841341
transform 1 0 1428 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1710841341
transform 1 0 1404 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1710841341
transform 1 0 1236 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1710841341
transform 1 0 1156 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1710841341
transform 1 0 1396 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1710841341
transform 1 0 1268 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3140
timestamp 1710841341
transform 1 0 1508 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1710841341
transform 1 0 1404 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1710841341
transform 1 0 1572 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1710841341
transform 1 0 1540 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1710841341
transform 1 0 1508 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1710841341
transform 1 0 1028 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1710841341
transform 1 0 916 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1710841341
transform 1 0 1244 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1710841341
transform 1 0 1180 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1710841341
transform 1 0 1148 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1710841341
transform 1 0 1148 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1710841341
transform 1 0 1268 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1710841341
transform 1 0 1188 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1710841341
transform 1 0 1212 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1710841341
transform 1 0 1140 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1710841341
transform 1 0 1164 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1710841341
transform 1 0 1132 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1710841341
transform 1 0 1268 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1710841341
transform 1 0 1220 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1710841341
transform 1 0 1292 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1710841341
transform 1 0 1116 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1710841341
transform 1 0 1196 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1710841341
transform 1 0 1164 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1710841341
transform 1 0 1292 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1710841341
transform 1 0 1212 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1710841341
transform 1 0 1036 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3166
timestamp 1710841341
transform 1 0 964 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1710841341
transform 1 0 1036 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1710841341
transform 1 0 972 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1710841341
transform 1 0 1460 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1710841341
transform 1 0 1132 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1710841341
transform 1 0 1164 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1710841341
transform 1 0 1036 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3173
timestamp 1710841341
transform 1 0 1036 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1710841341
transform 1 0 1012 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1710841341
transform 1 0 1020 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1710841341
transform 1 0 988 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1710841341
transform 1 0 740 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1710841341
transform 1 0 716 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1710841341
transform 1 0 644 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3180
timestamp 1710841341
transform 1 0 972 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1710841341
transform 1 0 908 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1710841341
transform 1 0 924 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1710841341
transform 1 0 884 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1710841341
transform 1 0 1556 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1710841341
transform 1 0 1500 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3186
timestamp 1710841341
transform 1 0 1068 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1710841341
transform 1 0 1012 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1710841341
transform 1 0 868 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1710841341
transform 1 0 788 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1710841341
transform 1 0 916 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1710841341
transform 1 0 852 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1710841341
transform 1 0 900 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1710841341
transform 1 0 884 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3194
timestamp 1710841341
transform 1 0 964 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1710841341
transform 1 0 892 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1710841341
transform 1 0 1428 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3197
timestamp 1710841341
transform 1 0 996 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1710841341
transform 1 0 908 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1710841341
transform 1 0 828 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1710841341
transform 1 0 884 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1710841341
transform 1 0 844 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1710841341
transform 1 0 940 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1710841341
transform 1 0 860 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1710841341
transform 1 0 748 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1710841341
transform 1 0 756 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3206
timestamp 1710841341
transform 1 0 612 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1710841341
transform 1 0 612 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1710841341
transform 1 0 532 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1710841341
transform 1 0 780 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1710841341
transform 1 0 716 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1710841341
transform 1 0 828 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1710841341
transform 1 0 708 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1710841341
transform 1 0 732 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1710841341
transform 1 0 660 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1710841341
transform 1 0 484 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1710841341
transform 1 0 444 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1710841341
transform 1 0 380 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1710841341
transform 1 0 508 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3219
timestamp 1710841341
transform 1 0 300 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3220
timestamp 1710841341
transform 1 0 268 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3221
timestamp 1710841341
transform 1 0 268 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1710841341
transform 1 0 228 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3223
timestamp 1710841341
transform 1 0 228 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1710841341
transform 1 0 188 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1710841341
transform 1 0 276 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1710841341
transform 1 0 204 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1710841341
transform 1 0 364 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3228
timestamp 1710841341
transform 1 0 204 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1710841341
transform 1 0 284 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1710841341
transform 1 0 172 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1710841341
transform 1 0 348 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1710841341
transform 1 0 188 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1710841341
transform 1 0 268 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3234
timestamp 1710841341
transform 1 0 180 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3235
timestamp 1710841341
transform 1 0 228 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1710841341
transform 1 0 204 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1710841341
transform 1 0 84 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3238
timestamp 1710841341
transform 1 0 380 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1710841341
transform 1 0 284 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3240
timestamp 1710841341
transform 1 0 220 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3241
timestamp 1710841341
transform 1 0 340 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1710841341
transform 1 0 316 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1710841341
transform 1 0 180 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_3244
timestamp 1710841341
transform 1 0 332 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1710841341
transform 1 0 244 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1710841341
transform 1 0 236 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3247
timestamp 1710841341
transform 1 0 92 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3248
timestamp 1710841341
transform 1 0 348 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1710841341
transform 1 0 116 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1710841341
transform 1 0 444 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1710841341
transform 1 0 348 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1710841341
transform 1 0 292 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1710841341
transform 1 0 212 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1710841341
transform 1 0 388 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1710841341
transform 1 0 220 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1710841341
transform 1 0 516 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1710841341
transform 1 0 420 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1710841341
transform 1 0 468 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1710841341
transform 1 0 284 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1710841341
transform 1 0 1524 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1710841341
transform 1 0 1404 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1710841341
transform 1 0 1708 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1710841341
transform 1 0 1572 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1710841341
transform 1 0 2516 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3265
timestamp 1710841341
transform 1 0 2420 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1710841341
transform 1 0 2676 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1710841341
transform 1 0 2580 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1710841341
transform 1 0 2676 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1710841341
transform 1 0 2556 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1710841341
transform 1 0 2012 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1710841341
transform 1 0 1916 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1710841341
transform 1 0 2668 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1710841341
transform 1 0 2540 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1710841341
transform 1 0 2668 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1710841341
transform 1 0 2556 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1710841341
transform 1 0 2668 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1710841341
transform 1 0 2612 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1710841341
transform 1 0 2668 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1710841341
transform 1 0 2540 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1710841341
transform 1 0 2564 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1710841341
transform 1 0 2412 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1710841341
transform 1 0 2508 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1710841341
transform 1 0 2364 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1710841341
transform 1 0 2532 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1710841341
transform 1 0 2404 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1710841341
transform 1 0 2084 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1710841341
transform 1 0 1956 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1710841341
transform 1 0 444 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1710841341
transform 1 0 348 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3290
timestamp 1710841341
transform 1 0 172 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1710841341
transform 1 0 100 0 1 2395
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1710841341
transform 1 0 224 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1710841341
transform 1 0 1256 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1710841341
transform 1 0 1248 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1710841341
transform 1 0 1192 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1710841341
transform 1 0 376 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1710841341
transform 1 0 344 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1710841341
transform 1 0 248 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1710841341
transform 1 0 248 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1710841341
transform 1 0 160 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1710841341
transform 1 0 328 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1710841341
transform 1 0 560 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1710841341
transform 1 0 1088 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1710841341
transform 1 0 928 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1710841341
transform 1 0 1136 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1710841341
transform 1 0 968 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1710841341
transform 1 0 896 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1710841341
transform 1 0 1088 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1710841341
transform 1 0 976 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1710841341
transform 1 0 848 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1710841341
transform 1 0 1032 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1710841341
transform 1 0 800 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1710841341
transform 1 0 1144 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1710841341
transform 1 0 1024 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1710841341
transform 1 0 616 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1710841341
transform 1 0 728 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1710841341
transform 1 0 640 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1710841341
transform 1 0 1264 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1710841341
transform 1 0 544 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1710841341
transform 1 0 1000 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1710841341
transform 1 0 1232 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1710841341
transform 1 0 808 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1710841341
transform 1 0 944 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1710841341
transform 1 0 1336 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1710841341
transform 1 0 1208 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1710841341
transform 1 0 1136 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1710841341
transform 1 0 1440 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1710841341
transform 1 0 1144 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1710841341
transform 1 0 1536 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1710841341
transform 1 0 1376 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1710841341
transform 1 0 1360 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1710841341
transform 1 0 1560 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1710841341
transform 1 0 1528 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1710841341
transform 1 0 1296 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1710841341
transform 1 0 1200 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1710841341
transform 1 0 1256 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1710841341
transform 1 0 1312 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1710841341
transform 1 0 1656 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1710841341
transform 1 0 1168 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1710841341
transform 1 0 1528 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1710841341
transform 1 0 1760 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1710841341
transform 1 0 1464 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1710841341
transform 1 0 2112 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1710841341
transform 1 0 1712 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1710841341
transform 1 0 2216 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1710841341
transform 1 0 2272 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1710841341
transform 1 0 1240 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1710841341
transform 1 0 1104 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1710841341
transform 1 0 2288 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1710841341
transform 1 0 2072 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1710841341
transform 1 0 2552 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1710841341
transform 1 0 1592 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1710841341
transform 1 0 2512 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1710841341
transform 1 0 2240 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1710841341
transform 1 0 1984 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1710841341
transform 1 0 2616 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1710841341
transform 1 0 1648 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1710841341
transform 1 0 2560 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1710841341
transform 1 0 2368 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1710841341
transform 1 0 1824 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1710841341
transform 1 0 1528 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1710841341
transform 1 0 2240 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1710841341
transform 1 0 2336 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1710841341
transform 1 0 2104 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1710841341
transform 1 0 2128 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1710841341
transform 1 0 2112 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1710841341
transform 1 0 1848 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1710841341
transform 1 0 1792 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1710841341
transform 1 0 1496 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1710841341
transform 1 0 1640 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1710841341
transform 1 0 760 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1710841341
transform 1 0 1664 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1710841341
transform 1 0 1952 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1710841341
transform 1 0 1712 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1710841341
transform 1 0 1768 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1710841341
transform 1 0 1720 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1710841341
transform 1 0 1744 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1710841341
transform 1 0 1640 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1710841341
transform 1 0 2376 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_88
timestamp 1710841341
transform 1 0 2464 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_89
timestamp 1710841341
transform 1 0 1584 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1710841341
transform 1 0 2552 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_91
timestamp 1710841341
transform 1 0 2120 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_92
timestamp 1710841341
transform 1 0 1632 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1710841341
transform 1 0 2264 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_94
timestamp 1710841341
transform 1 0 1936 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_95
timestamp 1710841341
transform 1 0 1816 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1710841341
transform 1 0 1672 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_97
timestamp 1710841341
transform 1 0 1920 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_98
timestamp 1710841341
transform 1 0 1616 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1710841341
transform 1 0 1448 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_100
timestamp 1710841341
transform 1 0 1320 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_101
timestamp 1710841341
transform 1 0 1592 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1710841341
transform 1 0 1584 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_103
timestamp 1710841341
transform 1 0 1776 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1710841341
transform 1 0 1536 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1710841341
transform 1 0 1416 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_106
timestamp 1710841341
transform 1 0 1544 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_107
timestamp 1710841341
transform 1 0 1216 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_108
timestamp 1710841341
transform 1 0 1416 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_109
timestamp 1710841341
transform 1 0 1264 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_110
timestamp 1710841341
transform 1 0 1536 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_111
timestamp 1710841341
transform 1 0 1376 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_112
timestamp 1710841341
transform 1 0 1256 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1710841341
transform 1 0 760 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_114
timestamp 1710841341
transform 1 0 792 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_115
timestamp 1710841341
transform 1 0 928 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_116
timestamp 1710841341
transform 1 0 1472 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_117
timestamp 1710841341
transform 1 0 1296 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1710841341
transform 1 0 872 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_119
timestamp 1710841341
transform 1 0 1280 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_120
timestamp 1710841341
transform 1 0 1312 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1710841341
transform 1 0 984 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_122
timestamp 1710841341
transform 1 0 680 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1710841341
transform 1 0 472 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1710841341
transform 1 0 528 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1710841341
transform 1 0 168 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_126
timestamp 1710841341
transform 1 0 352 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_127
timestamp 1710841341
transform 1 0 504 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_128
timestamp 1710841341
transform 1 0 376 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_129
timestamp 1710841341
transform 1 0 504 0 1 1370
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1710841341
transform 1 0 632 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1710841341
transform 1 0 600 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1710841341
transform 1 0 840 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1710841341
transform 1 0 880 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1710841341
transform 1 0 904 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1710841341
transform 1 0 808 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1710841341
transform 1 0 1064 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1710841341
transform 1 0 1136 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1710841341
transform 1 0 440 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1710841341
transform 1 0 472 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1710841341
transform 1 0 560 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1710841341
transform 1 0 392 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1710841341
transform 1 0 648 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1710841341
transform 1 0 672 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1710841341
transform 1 0 728 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1710841341
transform 1 0 584 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1710841341
transform 1 0 1112 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1710841341
transform 1 0 1056 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1710841341
transform 1 0 936 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1710841341
transform 1 0 856 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1710841341
transform 1 0 1296 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1710841341
transform 1 0 1248 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1710841341
transform 1 0 1288 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1710841341
transform 1 0 1232 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1710841341
transform 1 0 1384 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1710841341
transform 1 0 1448 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1710841341
transform 1 0 1576 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1710841341
transform 1 0 1696 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1710841341
transform 1 0 1632 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1710841341
transform 1 0 1384 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1710841341
transform 1 0 1744 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1710841341
transform 1 0 1840 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1710841341
transform 1 0 1744 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1710841341
transform 1 0 1624 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1710841341
transform 1 0 1752 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1710841341
transform 1 0 1696 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1710841341
transform 1 0 2264 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1710841341
transform 1 0 2296 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1710841341
transform 1 0 2192 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1710841341
transform 1 0 2240 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1710841341
transform 1 0 2248 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1710841341
transform 1 0 2192 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1710841341
transform 1 0 2344 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1710841341
transform 1 0 2104 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1710841341
transform 1 0 2024 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1710841341
transform 1 0 2080 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1710841341
transform 1 0 2440 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1710841341
transform 1 0 2560 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_48
timestamp 1710841341
transform 1 0 2136 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_49
timestamp 1710841341
transform 1 0 2328 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_50
timestamp 1710841341
transform 1 0 2632 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_51
timestamp 1710841341
transform 1 0 2552 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_52
timestamp 1710841341
transform 1 0 2416 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_53
timestamp 1710841341
transform 1 0 2320 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_54
timestamp 1710841341
transform 1 0 2224 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1710841341
transform 1 0 1944 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_56
timestamp 1710841341
transform 1 0 2312 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_57
timestamp 1710841341
transform 1 0 1704 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_58
timestamp 1710841341
transform 1 0 1544 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_59
timestamp 1710841341
transform 1 0 2152 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_60
timestamp 1710841341
transform 1 0 1976 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_61
timestamp 1710841341
transform 1 0 2216 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_62
timestamp 1710841341
transform 1 0 2048 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_63
timestamp 1710841341
transform 1 0 1768 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_64
timestamp 1710841341
transform 1 0 1856 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_65
timestamp 1710841341
transform 1 0 2424 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_66
timestamp 1710841341
transform 1 0 2288 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_67
timestamp 1710841341
transform 1 0 2232 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_68
timestamp 1710841341
transform 1 0 2464 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_69
timestamp 1710841341
transform 1 0 2376 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_70
timestamp 1710841341
transform 1 0 2328 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_71
timestamp 1710841341
transform 1 0 2496 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_72
timestamp 1710841341
transform 1 0 2600 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_73
timestamp 1710841341
transform 1 0 2176 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_74
timestamp 1710841341
transform 1 0 2120 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_75
timestamp 1710841341
transform 1 0 2160 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_76
timestamp 1710841341
transform 1 0 2224 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_77
timestamp 1710841341
transform 1 0 1864 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_78
timestamp 1710841341
transform 1 0 1808 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_79
timestamp 1710841341
transform 1 0 1864 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_80
timestamp 1710841341
transform 1 0 1960 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_81
timestamp 1710841341
transform 1 0 1688 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_82
timestamp 1710841341
transform 1 0 1576 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_83
timestamp 1710841341
transform 1 0 888 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_84
timestamp 1710841341
transform 1 0 728 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_85
timestamp 1710841341
transform 1 0 1336 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_86
timestamp 1710841341
transform 1 0 1384 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_87
timestamp 1710841341
transform 1 0 1384 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_88
timestamp 1710841341
transform 1 0 848 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_89
timestamp 1710841341
transform 1 0 576 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_90
timestamp 1710841341
transform 1 0 1448 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_91
timestamp 1710841341
transform 1 0 592 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_92
timestamp 1710841341
transform 1 0 1192 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_93
timestamp 1710841341
transform 1 0 1248 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_94
timestamp 1710841341
transform 1 0 704 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_95
timestamp 1710841341
transform 1 0 632 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_96
timestamp 1710841341
transform 1 0 1456 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_97
timestamp 1710841341
transform 1 0 1344 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_98
timestamp 1710841341
transform 1 0 688 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_99
timestamp 1710841341
transform 1 0 992 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_100
timestamp 1710841341
transform 1 0 936 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_101
timestamp 1710841341
transform 1 0 648 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_102
timestamp 1710841341
transform 1 0 1416 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_103
timestamp 1710841341
transform 1 0 1376 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_104
timestamp 1710841341
transform 1 0 1328 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_105
timestamp 1710841341
transform 1 0 536 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_106
timestamp 1710841341
transform 1 0 600 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_107
timestamp 1710841341
transform 1 0 1408 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_108
timestamp 1710841341
transform 1 0 648 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_109
timestamp 1710841341
transform 1 0 232 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_110
timestamp 1710841341
transform 1 0 240 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_111
timestamp 1710841341
transform 1 0 328 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_112
timestamp 1710841341
transform 1 0 408 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_113
timestamp 1710841341
transform 1 0 232 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_114
timestamp 1710841341
transform 1 0 304 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_115
timestamp 1710841341
transform 1 0 272 0 1 2370
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1710841341
transform 1 0 160 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1710841341
transform 1 0 272 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1710841341
transform 1 0 200 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1710841341
transform 1 0 168 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1710841341
transform 1 0 440 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1710841341
transform 1 0 144 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1710841341
transform 1 0 344 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1710841341
transform 1 0 840 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1710841341
transform 1 0 616 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1710841341
transform 1 0 408 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1710841341
transform 1 0 512 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1710841341
transform 1 0 456 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1710841341
transform 1 0 336 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1710841341
transform 1 0 576 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1710841341
transform 1 0 688 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1710841341
transform 1 0 736 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1710841341
transform 1 0 984 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1710841341
transform 1 0 1272 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1710841341
transform 1 0 1104 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1710841341
transform 1 0 296 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1710841341
transform 1 0 280 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1710841341
transform 1 0 592 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1710841341
transform 1 0 560 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1710841341
transform 1 0 408 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1710841341
transform 1 0 480 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1710841341
transform 1 0 664 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1710841341
transform 1 0 688 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1710841341
transform 1 0 440 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1710841341
transform 1 0 936 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1710841341
transform 1 0 392 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1710841341
transform 1 0 680 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1710841341
transform 1 0 576 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1710841341
transform 1 0 544 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1710841341
transform 1 0 1080 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1710841341
transform 1 0 1008 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1710841341
transform 1 0 968 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1710841341
transform 1 0 1296 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1710841341
transform 1 0 912 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1710841341
transform 1 0 600 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1710841341
transform 1 0 976 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1710841341
transform 1 0 1024 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1710841341
transform 1 0 936 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1710841341
transform 1 0 840 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1710841341
transform 1 0 1168 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1710841341
transform 1 0 1416 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1710841341
transform 1 0 1264 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1710841341
transform 1 0 1408 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1710841341
transform 1 0 1192 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1710841341
transform 1 0 1216 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1710841341
transform 1 0 1352 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1710841341
transform 1 0 1368 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1710841341
transform 1 0 1256 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1710841341
transform 1 0 1520 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1710841341
transform 1 0 1392 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1710841341
transform 1 0 1424 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1710841341
transform 1 0 1520 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1710841341
transform 1 0 1504 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1710841341
transform 1 0 1672 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1710841341
transform 1 0 1792 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1710841341
transform 1 0 1704 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1710841341
transform 1 0 1864 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1710841341
transform 1 0 1952 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1710841341
transform 1 0 1952 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1710841341
transform 1 0 1816 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1710841341
transform 1 0 1816 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1710841341
transform 1 0 1728 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1710841341
transform 1 0 1960 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1710841341
transform 1 0 2360 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1710841341
transform 1 0 2424 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1710841341
transform 1 0 1992 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1710841341
transform 1 0 1936 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1710841341
transform 1 0 2128 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1710841341
transform 1 0 2392 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1710841341
transform 1 0 2224 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1710841341
transform 1 0 2392 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1710841341
transform 1 0 1344 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1710841341
transform 1 0 2416 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1710841341
transform 1 0 2176 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1710841341
transform 1 0 2264 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1710841341
transform 1 0 2232 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1710841341
transform 1 0 1896 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1710841341
transform 1 0 2112 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1710841341
transform 1 0 2168 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1710841341
transform 1 0 2200 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1710841341
transform 1 0 1968 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1710841341
transform 1 0 2448 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1710841341
transform 1 0 1696 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1710841341
transform 1 0 2528 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1710841341
transform 1 0 2520 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1710841341
transform 1 0 2600 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1710841341
transform 1 0 2624 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1710841341
transform 1 0 2536 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1710841341
transform 1 0 2480 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1710841341
transform 1 0 1944 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1710841341
transform 1 0 2640 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1710841341
transform 1 0 2640 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1710841341
transform 1 0 2456 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1710841341
transform 1 0 2472 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1710841341
transform 1 0 2512 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1710841341
transform 1 0 1968 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1710841341
transform 1 0 1944 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1710841341
transform 1 0 2440 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1710841341
transform 1 0 2480 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1710841341
transform 1 0 816 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1710841341
transform 1 0 1896 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1710841341
transform 1 0 2240 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1710841341
transform 1 0 2488 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1710841341
transform 1 0 2576 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1710841341
transform 1 0 1344 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1710841341
transform 1 0 2288 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1710841341
transform 1 0 1960 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1710841341
transform 1 0 1832 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1710841341
transform 1 0 1872 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1710841341
transform 1 0 1176 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1710841341
transform 1 0 1720 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1710841341
transform 1 0 2456 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1710841341
transform 1 0 2584 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1710841341
transform 1 0 2216 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1710841341
transform 1 0 1896 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1710841341
transform 1 0 856 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1710841341
transform 1 0 2528 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1710841341
transform 1 0 2520 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1710841341
transform 1 0 2432 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1710841341
transform 1 0 2416 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1710841341
transform 1 0 2536 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1710841341
transform 1 0 1872 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_126
timestamp 1710841341
transform 1 0 1120 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_127
timestamp 1710841341
transform 1 0 2632 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_128
timestamp 1710841341
transform 1 0 2416 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_129
timestamp 1710841341
transform 1 0 2520 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_130
timestamp 1710841341
transform 1 0 2544 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_131
timestamp 1710841341
transform 1 0 2328 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_132
timestamp 1710841341
transform 1 0 2248 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_133
timestamp 1710841341
transform 1 0 2224 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_134
timestamp 1710841341
transform 1 0 2072 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_135
timestamp 1710841341
transform 1 0 2344 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_136
timestamp 1710841341
transform 1 0 1752 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_137
timestamp 1710841341
transform 1 0 2320 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_138
timestamp 1710841341
transform 1 0 2152 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_139
timestamp 1710841341
transform 1 0 2176 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_140
timestamp 1710841341
transform 1 0 2280 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_141
timestamp 1710841341
transform 1 0 2000 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_142
timestamp 1710841341
transform 1 0 1872 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_143
timestamp 1710841341
transform 1 0 2040 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_144
timestamp 1710841341
transform 1 0 2040 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_145
timestamp 1710841341
transform 1 0 2032 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_146
timestamp 1710841341
transform 1 0 1984 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_147
timestamp 1710841341
transform 1 0 1784 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_148
timestamp 1710841341
transform 1 0 1824 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_149
timestamp 1710841341
transform 1 0 1928 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_150
timestamp 1710841341
transform 1 0 1760 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_151
timestamp 1710841341
transform 1 0 1816 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_152
timestamp 1710841341
transform 1 0 1816 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_153
timestamp 1710841341
transform 1 0 840 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_154
timestamp 1710841341
transform 1 0 1728 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_155
timestamp 1710841341
transform 1 0 1600 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_156
timestamp 1710841341
transform 1 0 1536 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_157
timestamp 1710841341
transform 1 0 1664 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_158
timestamp 1710841341
transform 1 0 984 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_159
timestamp 1710841341
transform 1 0 1440 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_160
timestamp 1710841341
transform 1 0 1096 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_161
timestamp 1710841341
transform 1 0 1048 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_162
timestamp 1710841341
transform 1 0 1288 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_163
timestamp 1710841341
transform 1 0 1368 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_164
timestamp 1710841341
transform 1 0 1128 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_165
timestamp 1710841341
transform 1 0 960 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_166
timestamp 1710841341
transform 1 0 1136 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_167
timestamp 1710841341
transform 1 0 1304 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_168
timestamp 1710841341
transform 1 0 1088 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_169
timestamp 1710841341
transform 1 0 904 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_170
timestamp 1710841341
transform 1 0 992 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_171
timestamp 1710841341
transform 1 0 784 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_172
timestamp 1710841341
transform 1 0 720 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_173
timestamp 1710841341
transform 1 0 768 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_174
timestamp 1710841341
transform 1 0 816 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_175
timestamp 1710841341
transform 1 0 488 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_176
timestamp 1710841341
transform 1 0 1456 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_177
timestamp 1710841341
transform 1 0 976 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_178
timestamp 1710841341
transform 1 0 768 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_179
timestamp 1710841341
transform 1 0 832 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_180
timestamp 1710841341
transform 1 0 632 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_181
timestamp 1710841341
transform 1 0 760 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_182
timestamp 1710841341
transform 1 0 200 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_183
timestamp 1710841341
transform 1 0 224 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_184
timestamp 1710841341
transform 1 0 432 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_185
timestamp 1710841341
transform 1 0 480 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_186
timestamp 1710841341
transform 1 0 136 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_187
timestamp 1710841341
transform 1 0 88 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_0
timestamp 1710841341
transform 1 0 192 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1710841341
transform 1 0 104 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1710841341
transform 1 0 200 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1710841341
transform 1 0 88 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1710841341
transform 1 0 248 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1710841341
transform 1 0 288 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1710841341
transform 1 0 112 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1710841341
transform 1 0 192 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1710841341
transform 1 0 80 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1710841341
transform 1 0 264 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1710841341
transform 1 0 248 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1710841341
transform 1 0 232 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1710841341
transform 1 0 88 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1710841341
transform 1 0 184 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1710841341
transform 1 0 88 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1710841341
transform 1 0 240 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1710841341
transform 1 0 200 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1710841341
transform 1 0 640 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1710841341
transform 1 0 688 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1710841341
transform 1 0 696 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1710841341
transform 1 0 440 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1710841341
transform 1 0 624 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1710841341
transform 1 0 536 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1710841341
transform 1 0 472 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1710841341
transform 1 0 560 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1710841341
transform 1 0 688 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1710841341
transform 1 0 776 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1710841341
transform 1 0 680 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1710841341
transform 1 0 696 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1710841341
transform 1 0 688 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1710841341
transform 1 0 928 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1710841341
transform 1 0 1032 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1710841341
transform 1 0 1096 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1710841341
transform 1 0 952 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1710841341
transform 1 0 1008 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1710841341
transform 1 0 1152 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1710841341
transform 1 0 1024 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1710841341
transform 1 0 1088 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1710841341
transform 1 0 336 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1710841341
transform 1 0 312 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1710841341
transform 1 0 576 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1710841341
transform 1 0 744 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1710841341
transform 1 0 736 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1710841341
transform 1 0 712 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1710841341
transform 1 0 632 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1710841341
transform 1 0 528 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1710841341
transform 1 0 912 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1710841341
transform 1 0 1008 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1710841341
transform 1 0 848 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1710841341
transform 1 0 1288 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1710841341
transform 1 0 1296 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1710841341
transform 1 0 1240 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1710841341
transform 1 0 1464 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1710841341
transform 1 0 1416 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1710841341
transform 1 0 1464 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1710841341
transform 1 0 1616 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1710841341
transform 1 0 1568 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1710841341
transform 1 0 1536 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1710841341
transform 1 0 1632 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1710841341
transform 1 0 1584 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1710841341
transform 1 0 1568 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1710841341
transform 1 0 1672 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1710841341
transform 1 0 1832 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1710841341
transform 1 0 1880 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1710841341
transform 1 0 1776 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1710841341
transform 1 0 1832 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1710841341
transform 1 0 1896 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1710841341
transform 1 0 1960 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1710841341
transform 1 0 1472 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1710841341
transform 1 0 1416 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1710841341
transform 1 0 1728 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1710841341
transform 1 0 1632 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1710841341
transform 1 0 1568 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1710841341
transform 1 0 2296 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1710841341
transform 1 0 2144 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1710841341
transform 1 0 2112 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1710841341
transform 1 0 1976 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1710841341
transform 1 0 2240 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1710841341
transform 1 0 2224 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1710841341
transform 1 0 2160 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1710841341
transform 1 0 2376 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1710841341
transform 1 0 2624 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1710841341
transform 1 0 2624 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1710841341
transform 1 0 2584 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1710841341
transform 1 0 2568 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1710841341
transform 1 0 2512 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1710841341
transform 1 0 2080 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1710841341
transform 1 0 2024 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1710841341
transform 1 0 2280 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1710841341
transform 1 0 2504 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1710841341
transform 1 0 2144 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1710841341
transform 1 0 2192 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1710841341
transform 1 0 1848 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1710841341
transform 1 0 1736 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1710841341
transform 1 0 1656 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1710841341
transform 1 0 760 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1710841341
transform 1 0 1800 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1710841341
transform 1 0 2088 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1710841341
transform 1 0 2344 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1710841341
transform 1 0 2288 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1710841341
transform 1 0 1856 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1710841341
transform 1 0 1840 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1710841341
transform 1 0 1072 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1710841341
transform 1 0 1920 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1710841341
transform 1 0 2152 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1710841341
transform 1 0 2120 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1710841341
transform 1 0 2096 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1710841341
transform 1 0 1792 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1710841341
transform 1 0 1696 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1710841341
transform 1 0 928 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1710841341
transform 1 0 1688 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1710841341
transform 1 0 2384 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1710841341
transform 1 0 2344 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1710841341
transform 1 0 2168 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1710841341
transform 1 0 1904 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1710841341
transform 1 0 2152 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1710841341
transform 1 0 2472 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1710841341
transform 1 0 2496 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1710841341
transform 1 0 2552 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1710841341
transform 1 0 2168 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1710841341
transform 1 0 1648 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1710841341
transform 1 0 2176 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1710841341
transform 1 0 2248 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1710841341
transform 1 0 1928 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1710841341
transform 1 0 1856 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1710841341
transform 1 0 1944 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1710841341
transform 1 0 1632 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1710841341
transform 1 0 1760 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1710841341
transform 1 0 1640 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1710841341
transform 1 0 1576 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1710841341
transform 1 0 1512 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1710841341
transform 1 0 1528 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1710841341
transform 1 0 1264 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1710841341
transform 1 0 1328 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1710841341
transform 1 0 1312 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1710841341
transform 1 0 1416 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1710841341
transform 1 0 1304 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1710841341
transform 1 0 1320 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1710841341
transform 1 0 1256 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1710841341
transform 1 0 1352 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1710841341
transform 1 0 1096 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1710841341
transform 1 0 1144 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1710841341
transform 1 0 1208 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1710841341
transform 1 0 1256 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1710841341
transform 1 0 1376 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1710841341
transform 1 0 1192 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1710841341
transform 1 0 1128 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1710841341
transform 1 0 1136 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1710841341
transform 1 0 1248 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1710841341
transform 1 0 1144 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1710841341
transform 1 0 960 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1710841341
transform 1 0 1016 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1710841341
transform 1 0 1080 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1710841341
transform 1 0 1088 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1710841341
transform 1 0 1040 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1710841341
transform 1 0 1000 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1710841341
transform 1 0 1000 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1710841341
transform 1 0 1128 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1710841341
transform 1 0 1040 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1710841341
transform 1 0 840 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1710841341
transform 1 0 896 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1710841341
transform 1 0 880 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1710841341
transform 1 0 936 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_163
timestamp 1710841341
transform 1 0 880 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_164
timestamp 1710841341
transform 1 0 800 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_165
timestamp 1710841341
transform 1 0 752 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_166
timestamp 1710841341
transform 1 0 616 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_167
timestamp 1710841341
transform 1 0 800 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_168
timestamp 1710841341
transform 1 0 912 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_169
timestamp 1710841341
transform 1 0 400 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_170
timestamp 1710841341
transform 1 0 344 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_171
timestamp 1710841341
transform 1 0 248 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_172
timestamp 1710841341
transform 1 0 336 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_173
timestamp 1710841341
transform 1 0 256 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_174
timestamp 1710841341
transform 1 0 320 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_175
timestamp 1710841341
transform 1 0 240 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_176
timestamp 1710841341
transform 1 0 80 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_177
timestamp 1710841341
transform 1 0 360 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_178
timestamp 1710841341
transform 1 0 440 0 -1 2170
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1710841341
transform 1 0 392 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1710841341
transform 1 0 520 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1710841341
transform 1 0 512 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1710841341
transform 1 0 408 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1710841341
transform 1 0 624 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1710841341
transform 1 0 1200 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1710841341
transform 1 0 1280 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1710841341
transform 1 0 520 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1710841341
transform 1 0 336 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1710841341
transform 1 0 848 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1710841341
transform 1 0 600 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1710841341
transform 1 0 792 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1710841341
transform 1 0 368 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1710841341
transform 1 0 472 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1710841341
transform 1 0 1168 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1710841341
transform 1 0 1080 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1710841341
transform 1 0 848 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1710841341
transform 1 0 920 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1710841341
transform 1 0 880 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1710841341
transform 1 0 1360 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1710841341
transform 1 0 1200 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1710841341
transform 1 0 960 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1710841341
transform 1 0 1144 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1710841341
transform 1 0 1304 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1710841341
transform 1 0 1464 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1710841341
transform 1 0 920 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1710841341
transform 1 0 1416 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1710841341
transform 1 0 1568 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1710841341
transform 1 0 1608 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1710841341
transform 1 0 1792 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1710841341
transform 1 0 1744 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1710841341
transform 1 0 1800 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1710841341
transform 1 0 1896 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1710841341
transform 1 0 1784 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1710841341
transform 1 0 1784 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1710841341
transform 1 0 1888 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_36
timestamp 1710841341
transform 1 0 2368 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_37
timestamp 1710841341
transform 1 0 2064 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_38
timestamp 1710841341
transform 1 0 2040 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1710841341
transform 1 0 2312 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_40
timestamp 1710841341
transform 1 0 2072 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_41
timestamp 1710841341
transform 1 0 2352 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1710841341
transform 1 0 2328 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_43
timestamp 1710841341
transform 1 0 2040 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_44
timestamp 1710841341
transform 1 0 2136 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_45
timestamp 1710841341
transform 1 0 2064 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_46
timestamp 1710841341
transform 1 0 2584 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_47
timestamp 1710841341
transform 1 0 2528 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_48
timestamp 1710841341
transform 1 0 2400 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_49
timestamp 1710841341
transform 1 0 2024 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_50
timestamp 1710841341
transform 1 0 2616 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_51
timestamp 1710841341
transform 1 0 2512 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_52
timestamp 1710841341
transform 1 0 2448 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_53
timestamp 1710841341
transform 1 0 2032 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_54
timestamp 1710841341
transform 1 0 2040 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_55
timestamp 1710841341
transform 1 0 2376 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_56
timestamp 1710841341
transform 1 0 2280 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_57
timestamp 1710841341
transform 1 0 2424 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_58
timestamp 1710841341
transform 1 0 2480 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_59
timestamp 1710841341
transform 1 0 1032 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_60
timestamp 1710841341
transform 1 0 1984 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_61
timestamp 1710841341
transform 1 0 1784 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_62
timestamp 1710841341
transform 1 0 1776 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_63
timestamp 1710841341
transform 1 0 912 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_64
timestamp 1710841341
transform 1 0 2320 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_65
timestamp 1710841341
transform 1 0 2504 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_66
timestamp 1710841341
transform 1 0 1968 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_67
timestamp 1710841341
transform 1 0 2448 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_68
timestamp 1710841341
transform 1 0 2344 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_69
timestamp 1710841341
transform 1 0 2072 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_70
timestamp 1710841341
transform 1 0 2560 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_71
timestamp 1710841341
transform 1 0 2600 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_72
timestamp 1710841341
transform 1 0 2240 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_73
timestamp 1710841341
transform 1 0 2272 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_74
timestamp 1710841341
transform 1 0 2336 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_75
timestamp 1710841341
transform 1 0 2216 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_76
timestamp 1710841341
transform 1 0 1944 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_77
timestamp 1710841341
transform 1 0 2080 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_78
timestamp 1710841341
transform 1 0 2024 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_79
timestamp 1710841341
transform 1 0 2008 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_80
timestamp 1710841341
transform 1 0 1872 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_81
timestamp 1710841341
transform 1 0 1752 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_82
timestamp 1710841341
transform 1 0 1648 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_83
timestamp 1710841341
transform 1 0 1712 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_84
timestamp 1710841341
transform 1 0 1472 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_85
timestamp 1710841341
transform 1 0 1456 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_86
timestamp 1710841341
transform 1 0 1048 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_87
timestamp 1710841341
transform 1 0 1256 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_88
timestamp 1710841341
transform 1 0 1112 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_89
timestamp 1710841341
transform 1 0 888 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_90
timestamp 1710841341
transform 1 0 1184 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_91
timestamp 1710841341
transform 1 0 480 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_92
timestamp 1710841341
transform 1 0 192 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_93
timestamp 1710841341
transform 1 0 152 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_94
timestamp 1710841341
transform 1 0 272 0 -1 2170
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1710841341
transform 1 0 672 0 -1 1970
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1710841341
transform 1 0 168 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1710841341
transform 1 0 344 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1710841341
transform 1 0 160 0 -1 770
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1710841341
transform 1 0 752 0 -1 1570
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1710841341
transform 1 0 1024 0 -1 1770
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1710841341
transform 1 0 528 0 1 1970
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1710841341
transform 1 0 200 0 -1 2170
box -8 -3 40 105
use OR2X2  OR2X2_0
timestamp 1710841341
transform 1 0 496 0 1 1570
box -7 -3 35 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1710841341
transform 1 0 2720 0 1 2517
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1710841341
transform 1 0 2720 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1710841341
transform 1 0 24 0 1 2517
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1710841341
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1710841341
transform 1 0 2696 0 1 2493
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1710841341
transform 1 0 2696 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1710841341
transform 1 0 48 0 1 2493
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1710841341
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1710841341
transform 1 0 2720 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1710841341
transform 1 0 2720 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1710841341
transform 1 0 2720 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1710841341
transform 1 0 2720 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1710841341
transform 1 0 2720 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1710841341
transform 1 0 2720 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1710841341
transform 1 0 2720 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1710841341
transform 1 0 2720 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1710841341
transform 1 0 2720 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1710841341
transform 1 0 2720 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1710841341
transform 1 0 2720 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1710841341
transform 1 0 2720 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1710841341
transform 1 0 2720 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1710841341
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1710841341
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1710841341
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1710841341
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1710841341
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1710841341
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1710841341
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1710841341
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1710841341
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1710841341
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1710841341
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1710841341
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1710841341
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1710841341
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1710841341
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1710841341
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1710841341
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1710841341
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1710841341
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1710841341
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1710841341
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1710841341
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1710841341
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1710841341
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1710841341
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1710841341
transform 1 0 2696 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1710841341
transform 1 0 2696 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1710841341
transform 1 0 2696 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1710841341
transform 1 0 2696 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1710841341
transform 1 0 2696 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1710841341
transform 1 0 2696 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1710841341
transform 1 0 2696 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1710841341
transform 1 0 2696 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1710841341
transform 1 0 2696 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1710841341
transform 1 0 2696 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1710841341
transform 1 0 2696 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1710841341
transform 1 0 2696 0 1 2370
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1710841341
transform 1 0 240 0 -1 1770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1710841341
transform 1 0 224 0 1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1710841341
transform 1 0 336 0 1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1710841341
transform 1 0 128 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1710841341
transform 1 0 72 0 1 1570
box -8 -3 64 105
<< labels >>
rlabel electrodecontact s 356 2395 356 2395 4 in_clka
rlabel electrodecontact s 2636 145 2636 145 4 in_clkb
rlabel electrodecontact s 84 1345 84 1345 4 in_restart
rlabel electrodecontact s 172 2415 172 2415 4 in_move[1]
rlabel electrodecontact s 76 2405 76 2405 4 in_move[0]
rlabel metal1 220 1325 220 1325 4 board_out[31]
rlabel electrodecontact s 204 925 204 925 4 board_out[30]
rlabel metal1 180 325 180 325 4 board_out[29]
rlabel metal1 372 1015 372 1015 4 board_out[28]
rlabel metal1 420 725 420 725 4 board_out[27]
rlabel metal1 740 615 740 615 4 board_out[26]
rlabel metal1 1068 615 1068 615 4 board_out[25]
rlabel electrodecontact s 252 215 252 215 4 board_out[24]
rlabel metal1 332 125 332 125 4 board_out[23]
rlabel electrodecontact s 820 125 820 125 4 board_out[22]
rlabel electrodecontact s 1148 125 1148 125 4 board_out[21]
rlabel electrodecontact s 1716 125 1716 125 4 board_out[20]
rlabel metal1 1924 125 1924 125 4 board_out[19]
rlabel electrodecontact s 2084 125 2084 125 4 board_out[18]
rlabel metal1 1932 725 1932 725 4 board_out[17]
rlabel electrodecontact s 2532 925 2532 925 4 board_out[16]
rlabel metal1 2500 615 2500 615 4 board_out[15]
rlabel electrodecontact s 2564 125 2564 125 4 board_out[14]
rlabel electrodecontact s 2668 615 2668 615 4 board_out[13]
rlabel electrodecontact s 2668 1215 2668 1215 4 board_out[12]
rlabel electrodecontact s 2668 1415 2668 1415 4 board_out[11]
rlabel electrodecontact s 2668 1615 2668 1615 4 board_out[10]
rlabel electrodecontact s 2012 1925 2012 1925 4 board_out[9]
rlabel metal1 2668 1815 2668 1815 4 board_out[8]
rlabel metal1 2668 2015 2668 2015 4 board_out[7]
rlabel metal1 2500 2415 2500 2415 4 board_out[6]
rlabel electrodecontact s 2148 2415 2148 2415 4 board_out[5]
rlabel electrodecontact s 1708 2415 1708 2415 4 board_out[4]
rlabel electrodecontact s 1524 2415 1524 2415 4 board_out[3]
rlabel metal1 1188 2415 1188 2415 4 board_out[2]
rlabel metal1 1076 2415 1076 2415 4 board_out[1]
rlabel metal1 908 2415 908 2415 4 board_out[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 4788.000 12825.001 4788.000 14355.001 
<< end >>
