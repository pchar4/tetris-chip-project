magic
tech scmos
timestamp 1712256841
<< end >>
