magic
tech scmos
timestamp 1711307567
<< m2contact >>
rect -2 -2 2 2
<< end >>
