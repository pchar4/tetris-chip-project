magic
tech scmos
timestamp 1710841341
<< m2contact >>
rect -2 -2 2 2
<< end >>
