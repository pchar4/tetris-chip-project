magic
tech scmos
timestamp 1713638986
<< metal1 >>
rect -1366 4092 -1327 4120
rect -1057 4089 -1030 4126
rect -773 4086 -725 4121
rect -473 4089 -427 4120
rect -162 4090 -124 4120
rect 135 4094 181 4128
rect 431 4091 477 4125
rect 732 4091 773 4124
rect 1039 4095 1075 4121
rect 1333 4098 1391 4125
rect 1636 4102 1672 4118
rect 1928 4097 1969 4117
rect 2228 4094 2265 4114
rect 2844 4104 2866 4117
rect 3133 4092 3167 4108
rect -1389 3386 -1385 3402
rect -1471 3382 -1385 3386
rect -1089 3386 -1085 3402
rect -1171 3382 -1085 3386
rect -789 3386 -785 3402
rect -871 3382 -785 3386
rect -489 3386 -485 3402
rect -571 3382 -485 3386
rect -189 3386 -185 3402
rect -271 3382 -185 3386
rect 111 3386 115 3402
rect 29 3382 115 3386
rect 435 3360 458 3407
rect 711 3386 715 3402
rect 629 3382 715 3386
rect 1011 3386 1015 3402
rect 929 3382 1015 3386
rect 1311 3386 1315 3402
rect 1229 3382 1315 3386
rect 1611 3386 1615 3402
rect 1529 3382 1615 3386
rect 1911 3386 1915 3402
rect 1829 3382 1915 3386
rect 2211 3386 2215 3402
rect 2129 3382 2215 3386
rect 2811 3386 2815 3402
rect 2729 3382 2815 3386
rect 3111 3386 3115 3388
rect 3029 3382 3115 3386
rect 435 3337 903 3360
rect -2229 3227 -2200 3273
rect -1490 3211 -1482 3215
rect -1486 3129 -1482 3211
rect -2222 2934 -2193 2981
rect -1502 2911 -1482 2915
rect -1486 2829 -1482 2911
rect 880 2676 903 3337
rect -2226 2635 -2197 2671
rect -880 2652 -802 2671
rect -1502 2611 -1482 2615
rect -1486 2529 -1482 2611
rect -2219 2326 -2188 2374
rect -1502 2311 -1482 2315
rect -1486 2229 -1482 2311
rect -1486 1789 -1482 1871
rect -1488 1785 -1482 1789
rect -2226 1718 -2203 1775
rect -2228 1435 -2194 1467
rect -1490 1411 -1482 1415
rect -1486 1329 -1482 1411
rect -2227 1137 -2200 1173
rect -1489 1111 -1482 1115
rect -1486 1029 -1482 1111
rect -880 1002 -861 2652
rect -1454 983 -861 1002
rect -2224 828 -2191 864
rect -1489 811 -1482 815
rect -1486 729 -1482 811
rect -2216 527 -2189 574
rect -1491 511 -1482 515
rect -1486 429 -1482 511
rect -1454 259 -1435 983
rect -1489 240 -1435 259
rect -1486 -11 -1482 71
rect -1490 -15 -1482 -11
rect -2219 -75 -2192 -32
rect -2218 -366 -2194 -331
rect -1490 -389 -1482 -385
rect -1486 -471 -1482 -389
rect -2224 -665 -2193 -628
rect -1493 -689 -1482 -685
rect -1486 -771 -1482 -689
rect -2227 -977 -2197 -934
rect -1494 -989 -1482 -985
rect -1486 -1071 -1482 -989
rect -2220 -1267 -2201 -1235
rect -1471 -1376 -1385 -1372
rect -1389 -1392 -1385 -1376
rect -1171 -1386 -1085 -1382
rect -1089 -1391 -1085 -1386
rect -871 -1386 -785 -1382
rect -789 -1390 -785 -1386
rect 29 -1386 115 -1382
rect 111 -1390 115 -1386
rect -1363 -2120 -1337 -2097
rect -1061 -2122 -1035 -2100
rect -761 -2124 -735 -2105
rect -458 -2123 -430 -2096
rect 140 -2118 171 -2098
rect 440 -2117 464 -2100
rect 743 -2117 773 -2098
rect 1035 -2117 1070 -2090
rect 1337 -2116 1359 -2101
<< m2contact >>
rect -1477 3381 -1471 3387
rect -1177 3381 -1171 3387
rect -877 3381 -871 3387
rect -577 3381 -571 3387
rect -277 3381 -271 3387
rect 23 3381 29 3387
rect 623 3381 629 3387
rect 923 3381 929 3387
rect 1223 3381 1229 3387
rect 1523 3381 1529 3387
rect 1823 3381 1829 3387
rect 2123 3381 2129 3387
rect 2723 3381 2729 3387
rect 3023 3381 3029 3387
rect -1487 3123 -1481 3129
rect -1487 2823 -1481 2829
rect -1487 2523 -1481 2529
rect -1487 2223 -1481 2229
rect -1487 1871 -1481 1877
rect -1487 1323 -1481 1329
rect -1487 1023 -1481 1029
rect -1487 723 -1481 729
rect -1487 423 -1481 429
rect -1487 71 -1481 77
rect -1487 -477 -1481 -471
rect -1487 -777 -1481 -771
rect -1487 -1077 -1481 -1071
rect -1477 -1377 -1471 -1371
rect -1177 -1387 -1171 -1381
rect -877 -1387 -871 -1381
rect 23 -1387 29 -1381
<< metal2 >>
rect -1456 3334 -1453 3381
rect -1156 3340 -1153 3381
rect -856 3346 -853 3381
rect -556 3352 -553 3381
rect -256 3358 -253 3381
rect 44 3364 47 3381
rect 650 3370 653 3381
rect 944 3370 947 3381
rect 650 3367 891 3370
rect 44 3361 885 3364
rect -256 3355 879 3358
rect -556 3349 873 3352
rect -856 3343 867 3346
rect -1156 3337 861 3340
rect -1456 3331 855 3334
rect -1481 3150 -1431 3153
rect -1481 2850 -1437 2853
rect -1481 2550 -1443 2553
rect -1482 2250 -1449 2253
rect -1481 1853 -1455 1856
rect -1481 1350 -1461 1353
rect -1481 1050 -1467 1053
rect -1470 997 -1467 1050
rect -1464 1003 -1461 1350
rect -1458 1009 -1455 1853
rect -1452 1015 -1449 2250
rect -1446 1021 -1443 2550
rect -1440 1027 -1437 2850
rect -1434 1033 -1431 3150
rect 852 2787 855 3331
rect -887 2784 855 2787
rect -887 1595 -884 2784
rect 858 2781 861 3337
rect -881 2778 861 2781
rect -881 1625 -878 2778
rect 864 2775 867 3343
rect -875 2772 867 2775
rect -875 1695 -872 2772
rect 870 2769 873 3349
rect -869 2766 873 2769
rect -869 1775 -866 2766
rect 876 2763 879 3355
rect -863 2760 879 2763
rect -863 1835 -860 2760
rect 882 2757 885 3361
rect -857 2754 885 2757
rect -857 1895 -854 2754
rect 888 2751 891 3367
rect -851 2748 891 2751
rect 894 3367 947 3370
rect -851 2045 -848 2748
rect 894 2745 897 3367
rect 1244 3364 1247 3381
rect -845 2742 897 2745
rect 900 3361 1247 3364
rect -845 2205 -842 2742
rect 900 2739 903 3361
rect 1544 3358 1547 3381
rect -84 2736 903 2739
rect 906 3355 1547 3358
rect -84 2706 -81 2736
rect 906 2733 909 3355
rect 1844 3352 1847 3381
rect -36 2730 909 2733
rect 912 3349 1847 3352
rect -36 2705 -33 2730
rect 912 2727 915 3349
rect 2144 3346 2147 3381
rect -12 2724 915 2727
rect 918 3343 2147 3346
rect -12 2706 -9 2724
rect 918 2721 921 3343
rect 2744 3340 2747 3381
rect 4 2718 921 2721
rect 924 3337 2747 3340
rect 4 2705 7 2718
rect 924 2715 927 3337
rect 3044 3334 3047 3381
rect 20 2712 927 2715
rect 930 3331 3047 3334
rect 20 2706 23 2712
rect 930 2709 933 3331
rect 3273 3195 3288 3199
rect 3273 3129 3277 3195
rect 3273 3123 3296 3129
rect 3273 2895 3288 2899
rect 3273 2829 3277 2895
rect 3273 2823 3296 2829
rect 116 2706 933 2709
rect 3273 2595 3288 2599
rect 3273 2529 3277 2595
rect 3273 2523 3296 2529
rect 3273 2295 3288 2299
rect 3273 2229 3277 2295
rect 3273 2223 3296 2229
rect -851 2042 -845 2045
rect 3273 1995 3288 1999
rect 3273 1929 3277 1995
rect 3273 1923 3296 1929
rect -857 1892 -845 1895
rect -863 1832 -845 1835
rect -869 1772 -845 1775
rect -875 1692 -845 1695
rect -881 1622 -845 1625
rect -887 1592 -845 1595
rect -887 1552 -845 1555
rect -887 1033 -884 1552
rect -1434 1030 -884 1033
rect -881 1412 -845 1415
rect -881 1027 -878 1412
rect 3273 1395 3288 1399
rect 3273 1329 3277 1395
rect 3273 1323 3296 1329
rect -1440 1024 -878 1027
rect -875 1252 -845 1255
rect -875 1021 -872 1252
rect -1446 1018 -872 1021
rect -869 1162 -845 1165
rect -869 1015 -866 1162
rect -1452 1012 -866 1015
rect -863 1102 -845 1105
rect -863 1009 -860 1102
rect 3273 1095 3288 1099
rect -1458 1006 -860 1009
rect -857 1082 -845 1085
rect -857 1003 -854 1082
rect 3273 1029 3277 1095
rect 3273 1023 3296 1029
rect -1464 1000 -854 1003
rect -1470 994 -842 997
rect -1470 988 -848 991
rect -1470 747 -1467 988
rect -1481 744 -1467 747
rect -1464 982 -854 985
rect -1464 453 -1461 982
rect -1481 450 -1461 453
rect -1458 976 -860 979
rect -1458 56 -1455 976
rect -1481 53 -1455 56
rect -1452 970 -866 973
rect -1452 -447 -1449 970
rect -1481 -450 -1449 -447
rect -1446 964 -872 967
rect -1446 -747 -1443 964
rect -1482 -750 -1443 -747
rect -1440 958 -878 961
rect -1440 -1047 -1437 958
rect -1481 -1050 -1437 -1047
rect -1434 952 -884 955
rect -1434 -1347 -1431 952
rect -887 305 -884 952
rect -881 325 -878 958
rect -875 355 -872 964
rect -869 375 -866 970
rect -863 765 -860 976
rect -857 795 -854 982
rect -851 865 -848 988
rect -845 915 -842 994
rect -851 862 -845 865
rect 3273 795 3288 799
rect -857 792 -845 795
rect -863 762 -845 765
rect 3273 729 3277 795
rect 3273 723 3296 729
rect 3273 495 3288 499
rect 3273 429 3277 495
rect 3273 423 3296 429
rect -869 372 -845 375
rect -875 352 -845 355
rect -881 322 -845 325
rect -887 302 -845 305
rect -887 282 -845 285
rect -887 -776 -884 282
rect -881 262 -845 265
rect -881 -770 -878 262
rect -875 242 -845 245
rect -875 -764 -872 242
rect -869 222 -845 225
rect -869 -758 -866 222
rect -863 202 -845 205
rect -863 -752 -860 202
rect 3273 195 3288 199
rect 3273 129 3277 195
rect 3273 123 3296 129
rect 3273 -405 3288 -401
rect 3273 -471 3277 -405
rect 3273 -477 3296 -471
rect 3273 -705 3288 -701
rect -164 -746 -161 -731
rect 260 -740 263 -728
rect 884 -734 887 -731
rect 884 -737 897 -734
rect 260 -743 891 -740
rect -164 -749 885 -746
rect -863 -755 879 -752
rect -869 -761 873 -758
rect -875 -767 867 -764
rect -881 -773 861 -770
rect -887 -779 855 -776
rect 852 -1331 855 -779
rect -1481 -1350 -1431 -1347
rect -1428 -1334 855 -1331
rect -1428 -1353 -1425 -1334
rect 858 -1337 861 -773
rect -1450 -1356 -1425 -1353
rect -1156 -1340 861 -1337
rect -1481 -1377 -1477 -1371
rect -1477 -1381 -1471 -1377
rect -1450 -1382 -1447 -1356
rect -1156 -1381 -1153 -1340
rect 864 -1343 867 -767
rect -856 -1346 867 -1343
rect -856 -1381 -853 -1346
rect 870 -1349 873 -761
rect -343 -1352 873 -1349
rect -577 -1377 -501 -1373
rect -577 -1381 -571 -1377
rect -505 -1392 -501 -1377
rect -343 -1381 -340 -1352
rect 876 -1355 879 -755
rect 44 -1358 879 -1355
rect 44 -1381 47 -1358
rect 882 -1361 885 -749
rect 557 -1364 885 -1361
rect 323 -1377 399 -1373
rect 323 -1381 329 -1377
rect 395 -1392 399 -1377
rect 557 -1381 560 -1364
rect 888 -1367 891 -743
rect 857 -1370 891 -1367
rect 894 -1367 897 -737
rect 940 -740 943 -728
rect 900 -743 943 -740
rect 900 -1361 903 -743
rect 3273 -771 3277 -705
rect 3273 -777 3296 -771
rect 3273 -1005 3288 -1001
rect 3273 -1071 3277 -1005
rect 3273 -1077 3296 -1071
rect 3273 -1305 3288 -1301
rect 900 -1364 1466 -1361
rect 894 -1370 1166 -1367
rect 623 -1377 699 -1373
rect 623 -1381 629 -1377
rect 695 -1392 699 -1377
rect 857 -1381 860 -1370
rect 923 -1377 999 -1374
rect 923 -1381 929 -1377
rect 995 -1392 999 -1377
rect 1163 -1381 1166 -1370
rect 1223 -1377 1299 -1373
rect 1223 -1381 1229 -1377
rect 1295 -1388 1299 -1377
rect 1463 -1382 1466 -1364
rect 3273 -1371 3277 -1305
rect 1823 -1377 1899 -1373
rect 1295 -1392 1299 -1391
rect 1823 -1396 1829 -1377
rect 1895 -1388 1899 -1377
rect 2123 -1377 2199 -1373
rect 2123 -1396 2129 -1377
rect 2195 -1388 2199 -1377
rect 2423 -1377 2499 -1373
rect 2423 -1396 2429 -1377
rect 2495 -1388 2499 -1377
rect 2723 -1377 2799 -1373
rect 2723 -1396 2729 -1377
rect 2795 -1388 2799 -1377
rect 3023 -1377 3099 -1373
rect 3273 -1377 3281 -1371
rect 3023 -1396 3029 -1377
rect 3095 -1388 3099 -1377
<< m3contact >>
rect -845 2200 -840 2205
rect -845 2040 -840 2045
rect -845 1890 -840 1895
rect -845 1830 -840 1835
rect -845 1770 -840 1775
rect -845 1690 -840 1695
rect -845 1620 -840 1625
rect -845 1590 -840 1595
rect -845 1552 -840 1557
rect -845 1412 -840 1417
rect -845 1252 -840 1257
rect -845 1162 -840 1167
rect -845 1102 -840 1107
rect -845 1082 -840 1087
rect -845 910 -840 915
rect -845 860 -840 865
rect -845 790 -840 795
rect -845 760 -840 765
rect -845 370 -840 375
rect -845 350 -840 355
rect -845 320 -840 325
rect -845 300 -840 305
rect -845 280 -840 285
rect -845 260 -840 265
rect -845 240 -840 245
rect -845 220 -840 225
rect -845 200 -840 205
<< metal3 >>
rect -846 2205 -839 2206
rect -846 2200 -845 2205
rect -840 2200 -839 2205
rect -846 2199 -839 2200
rect -846 2191 -841 2199
rect -846 2045 -839 2046
rect -846 2040 -845 2045
rect -840 2040 -839 2045
rect -846 2039 -839 2040
rect -846 2031 -841 2039
rect -846 1895 -839 1896
rect -846 1890 -845 1895
rect -840 1890 -839 1895
rect -846 1889 -839 1890
rect -846 1881 -841 1889
rect -846 1835 -839 1836
rect -846 1830 -845 1835
rect -840 1830 -839 1835
rect -846 1829 -839 1830
rect -846 1821 -841 1829
rect -846 1775 -839 1776
rect -846 1770 -845 1775
rect -840 1770 -839 1775
rect -846 1769 -839 1770
rect -846 1761 -841 1769
rect -846 1695 -839 1696
rect -846 1690 -845 1695
rect -840 1690 -839 1695
rect -846 1689 -839 1690
rect -846 1681 -841 1689
rect -846 1625 -839 1626
rect -846 1620 -845 1625
rect -840 1620 -839 1625
rect -846 1619 -839 1620
rect -846 1611 -841 1619
rect -846 1595 -839 1596
rect -846 1590 -845 1595
rect -840 1590 -839 1595
rect -846 1589 -839 1590
rect -846 1581 -841 1589
rect -846 1558 -841 1566
rect -846 1557 -839 1558
rect -846 1552 -845 1557
rect -840 1552 -839 1557
rect -846 1551 -839 1552
rect -846 1418 -841 1426
rect -846 1417 -839 1418
rect -846 1412 -845 1417
rect -840 1412 -839 1417
rect -846 1411 -839 1412
rect -846 1258 -841 1266
rect -846 1257 -839 1258
rect -846 1252 -845 1257
rect -840 1252 -839 1257
rect -846 1251 -839 1252
rect -846 1168 -841 1176
rect -846 1167 -839 1168
rect -846 1162 -845 1167
rect -840 1162 -839 1167
rect -846 1161 -839 1162
rect -846 1108 -841 1116
rect -846 1107 -839 1108
rect -846 1102 -845 1107
rect -840 1102 -839 1107
rect -846 1101 -839 1102
rect -846 1088 -841 1096
rect -846 1087 -839 1088
rect -846 1082 -845 1087
rect -840 1082 -839 1087
rect -846 1081 -839 1082
rect -846 915 -839 916
rect -846 910 -845 915
rect -840 910 -839 915
rect -846 909 -839 910
rect -846 901 -841 909
rect -846 865 -839 866
rect -846 860 -845 865
rect -840 860 -839 865
rect -846 859 -839 860
rect -846 851 -841 859
rect -846 795 -839 796
rect -846 790 -845 795
rect -840 790 -839 795
rect -846 789 -839 790
rect -846 781 -841 789
rect -846 765 -839 766
rect -846 760 -845 765
rect -840 760 -839 765
rect -846 759 -839 760
rect -846 751 -841 759
rect -846 375 -839 376
rect -846 370 -845 375
rect -840 370 -839 375
rect -846 369 -839 370
rect -846 361 -841 369
rect -846 355 -839 356
rect -846 350 -845 355
rect -840 350 -839 355
rect -846 349 -839 350
rect -846 341 -841 349
rect -846 325 -839 326
rect -846 320 -845 325
rect -840 320 -839 325
rect -846 319 -839 320
rect -846 311 -841 319
rect -846 305 -839 306
rect -846 300 -845 305
rect -840 300 -839 305
rect -846 299 -839 300
rect -846 291 -841 299
rect -846 285 -839 286
rect -846 280 -845 285
rect -840 280 -839 285
rect -846 279 -839 280
rect -846 271 -841 279
rect -846 265 -839 266
rect -846 260 -845 265
rect -840 260 -839 265
rect -846 259 -839 260
rect -846 251 -841 259
rect -846 245 -839 246
rect -846 240 -845 245
rect -840 240 -839 245
rect -846 239 -839 240
rect -846 231 -841 239
rect -846 225 -839 226
rect -846 220 -845 225
rect -840 220 -839 225
rect -846 219 -839 220
rect -846 211 -841 219
rect -846 205 -839 206
rect -846 200 -845 205
rect -840 200 -839 205
rect -846 199 -839 200
rect -846 191 -841 199
use PadFC  16_0
timestamp 1681001061
transform 1 0 -2500 0 1 3400
box 327 -3 1003 673
use PadFC  16_1
timestamp 1681001061
transform 0 1 3300 -1 0 4400
box 327 -3 1003 673
use PadFC  16_2
timestamp 1681001061
transform 0 -1 -1500 1 0 -2400
box 327 -3 1003 673
use PadFC  16_3
timestamp 1681001061
transform -1 0 4300 0 -1 -1400
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1711830429
transform 1 0 -1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1711830429
transform 1 0 -1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1711830429
transform 1 0 -900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1711830429
transform 1 0 -600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1711830429
transform 1 0 -300 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_5
timestamp 1711830429
transform 1 0 0 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1711830429
transform 1 0 600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1711830429
transform 1 0 900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1711830429
transform 1 0 1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1711830429
transform 0 -1 -1500 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1711830429
transform 0 -1 -1500 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1711830429
transform 0 -1 -1500 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1711830429
transform 0 -1 -1500 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_13
timestamp 1711830429
transform 0 -1 -1500 -1 0 1900
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1711830429
transform 0 -1 -1500 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1711830429
transform 0 -1 -1500 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1711830429
transform 0 -1 -1500 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1711830429
transform 0 1 3300 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1711830429
transform 0 1 3300 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_19
timestamp 1711830429
transform 0 1 3300 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1711830429
transform 0 1 3300 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1711830429
transform 0 1 3300 1 0 1900
box -36 -19 303 1000
use PadBiDir  17_22
timestamp 1711830429
transform 0 1 3300 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1711830429
transform 0 1 3300 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1711830429
transform 0 1 3300 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1711830429
transform 0 -1 -1500 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_26
timestamp 1711830429
transform 1 0 -1500 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1711830429
transform 1 0 -1200 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1711830429
transform 1 0 -900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1711830429
transform 1 0 -600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_30
timestamp 1711830429
transform 1 0 0 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1711830429
transform 1 0 300 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1711830429
transform 1 0 600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1711830429
transform 1 0 900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1711830429
transform 0 1 3300 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1711830429
transform 1 0 1200 0 -1 -1400
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1711831643
transform 1 0 300 0 1 3400
box -3 -16 303 1000
use PadVdd  18_1
timestamp 1711831643
transform 1 0 -300 0 -1 -1400
box -3 -16 303 1000
use PadGnd  19_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 2200
box -3 -11 303 1000
use PadGnd  19_1
timestamp 1711831454
transform 0 1 3300 -1 0 1900
box -3 -11 303 1000
use PadBiDir  PadBiDir_0
timestamp 1711830429
transform 1 0 1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_1
timestamp 1711830429
transform 1 0 1800 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_2
timestamp 1711830429
transform 1 0 2100 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_3
timestamp 1711830429
transform 1 0 2700 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_4
timestamp 1711830429
transform 1 0 3000 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_5
timestamp 1711830429
transform 1 0 1800 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_6
timestamp 1711830429
transform 1 0 2100 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_7
timestamp 1711830429
transform 1 0 2400 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_8
timestamp 1711830429
transform 1 0 2700 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_9
timestamp 1711830429
transform 1 0 3000 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_10
timestamp 1711830429
transform 0 -1 -1500 -1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_11
timestamp 1711830429
transform 0 -1 -1500 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_12
timestamp 1711830429
transform 0 -1 -1500 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_13
timestamp 1711830429
transform 0 -1 -1500 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_14
timestamp 1711830429
transform 0 -1 -1500 1 0 1300
box -36 -19 303 1000
use PadBiDir  PadBiDir_15
timestamp 1711830429
transform 0 1 3300 1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_16
timestamp 1711830429
transform 0 1 3300 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_17
timestamp 1711830429
transform 0 1 3300 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_18
timestamp 1711830429
transform 0 1 3300 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_19
timestamp 1711830429
transform 0 1 3300 1 0 1300
box -36 -19 303 1000
use PadGnd  PadGnd_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 400
box -3 -11 303 1000
use PadGnd  PadGnd_1
timestamp 1711831454
transform 0 1 3300 -1 0 100
box -3 -11 303 1000
use PadVdd  PadVdd_0
timestamp 1711831643
transform 1 0 2400 0 1 3400
box -3 -16 303 1000
use PadVdd  PadVdd_1
timestamp 1711831643
transform 1 0 1500 0 -1 -1400
box -3 -16 303 1000
use top_module  top_module_0
timestamp 1713453518
transform 1 0 -846 0 1 -731
box 0 0 3506 3440
<< labels >>
rlabel metal1 3149 4102 3149 4102 1 p_board_out[29]
rlabel metal1 2855 4111 2855 4111 1 p_board_out[25]
rlabel metal1 2246 4106 2246 4106 1 p_board_out[30]
rlabel metal1 1946 4107 1946 4107 1 p_board_out[31]
rlabel metal1 1651 4111 1651 4111 1 p_board_out[26]
rlabel metal1 1360 4113 1360 4113 1 p_board_out[27]
rlabel metal1 1054 4106 1054 4106 1 p_board_out[28]
rlabel metal1 754 4108 754 4108 1 p_board_out[24]
rlabel metal1 152 4111 152 4111 1 p_board_out[23]
rlabel metal1 -146 4108 -146 4108 1 p_board_out[22]
rlabel metal1 -445 4103 -445 4103 1 p_board_out[21]
rlabel metal1 -751 4104 -751 4104 1 p_board_out[20]
rlabel metal1 -1045 4110 -1045 4110 1 p_board_out[19]
rlabel metal1 -1345 4108 -1345 4108 1 p_board_out[18]
rlabel metal1 -2213 3252 -2213 3252 1 p_board_out[16]
rlabel metal1 -2206 2956 -2206 2956 1 p_board_out[17]
rlabel metal1 -2212 2649 -2212 2649 1 p_board_out[15]
rlabel metal1 -2203 2351 -2203 2351 1 p_board_out[14]
rlabel metal1 -2213 1751 -2213 1751 1 p_board_out[13]
rlabel metal1 -2209 1454 -2209 1454 1 p_board_out[12]
rlabel metal1 -2211 1153 -2211 1153 1 p_board_out[11]
rlabel metal1 -2205 845 -2205 845 1 p_board_out[8]
rlabel metal1 -2207 548 -2207 548 1 p_board_out[10]
rlabel metal1 -2202 -49 -2202 -49 1 p_board_out[9]
rlabel metal1 -2205 -347 -2205 -347 1 p_board_out[7]
rlabel metal1 -2205 -646 -2205 -646 1 p_board_out[6]
rlabel metal1 -2209 -953 -2209 -953 1 p_board_out[5]
rlabel metal1 -2210 -1252 -2210 -1252 1 p_board_out[4]
rlabel metal1 -1350 -2110 -1350 -2110 1 p_board_out[3]
rlabel metal1 -1049 -2113 -1049 -2113 1 p_board_out[2]
rlabel metal1 -750 -2115 -750 -2115 1 p_board_out[1]
rlabel metal1 -446 -2110 -446 -2110 1 p_in_clkb
rlabel metal1 153 -2108 153 -2108 1 p_board_out[0]
rlabel metal1 453 -2108 453 -2108 1 p_in_clka
rlabel metal1 755 -2106 755 -2106 1 p_in_restart
rlabel metal1 1052 -2104 1052 -2104 1 p_in_move[0]
rlabel metal1 1349 -2107 1349 -2107 1 p_in_move[1]
<< end >>
