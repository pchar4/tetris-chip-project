magic
tech scmos
timestamp 1711653199
<< m2contact >>
rect -2 -2 2 2
<< end >>
