magic
tech scmos
timestamp 1711307567
<< end >>
