magic
tech scmos
timestamp 1712020386
<< m2contact >>
rect -2 -2 2 2
<< end >>
