magic
tech scmos
timestamp 1712622712
<< m2contact >>
rect -2 -2 2 2
<< end >>
