magic
tech scmos
timestamp 1712256841
<< metal1 >>
rect 14 3307 3490 3327
rect 38 3283 3466 3303
rect 14 3267 3490 3273
rect 954 3233 980 3236
rect 1602 3233 1652 3236
rect 1842 3233 1860 3236
rect 1922 3233 1932 3236
rect 1946 3233 1980 3236
rect 588 3223 613 3226
rect 658 3216 661 3226
rect 954 3216 957 3233
rect 988 3223 997 3226
rect 1092 3223 1101 3226
rect 1252 3223 1277 3226
rect 1340 3223 1357 3226
rect 1436 3223 1469 3226
rect 1596 3223 1645 3226
rect 1868 3223 1885 3226
rect 1940 3223 1957 3226
rect 1964 3223 1973 3226
rect 2020 3223 2053 3226
rect 1274 3216 1277 3223
rect 1466 3216 1469 3223
rect 2106 3216 2109 3225
rect 2210 3216 2213 3225
rect 2428 3223 2437 3226
rect 2556 3223 2573 3226
rect 2908 3223 2941 3226
rect 3412 3223 3421 3226
rect 196 3213 221 3216
rect 252 3213 269 3216
rect 276 3213 285 3216
rect 332 3213 357 3216
rect 444 3213 461 3216
rect 506 3213 540 3216
rect 594 3213 620 3216
rect 658 3213 668 3216
rect 700 3213 717 3216
rect 722 3213 740 3216
rect 804 3213 829 3216
rect 914 3213 957 3216
rect 994 3213 1004 3216
rect 1010 3213 1044 3216
rect 1050 3213 1076 3216
rect 1090 3213 1124 3216
rect 1138 3213 1156 3216
rect 1274 3213 1285 3216
rect 1338 3213 1396 3216
rect 1412 3213 1421 3216
rect 1466 3213 1484 3216
rect 1498 3213 1532 3216
rect 1546 3213 1581 3216
rect 1682 3213 1700 3216
rect 1788 3213 1821 3216
rect 266 3205 269 3213
rect 722 3206 725 3213
rect 826 3206 829 3213
rect 644 3203 669 3206
rect 692 3203 725 3206
rect 764 3203 789 3206
rect 802 3203 812 3206
rect 826 3203 852 3206
rect 882 3203 892 3206
rect 1010 3203 1013 3213
rect 1140 3203 1148 3206
rect 1186 3203 1196 3206
rect 1282 3205 1285 3213
rect 1316 3203 1324 3206
rect 1362 3203 1388 3206
rect 1500 3203 1517 3206
rect 1554 3203 1564 3206
rect 1748 3203 1764 3206
rect 1900 3203 1909 3206
rect 770 3193 788 3196
rect 1706 3193 1740 3196
rect 1794 3193 1820 3196
rect 1874 3193 1892 3196
rect 1922 3193 1925 3214
rect 2106 3213 2124 3216
rect 2138 3213 2164 3216
rect 2178 3213 2196 3216
rect 2210 3213 2228 3216
rect 2258 3213 2276 3216
rect 2292 3213 2325 3216
rect 2332 3213 2349 3216
rect 2452 3213 2461 3216
rect 2468 3213 2509 3216
rect 2516 3213 2525 3216
rect 2530 3213 2540 3216
rect 2612 3213 2637 3216
rect 2668 3213 2701 3216
rect 2788 3213 2797 3216
rect 2922 3213 2956 3216
rect 2970 3213 2988 3216
rect 2994 3213 3045 3216
rect 3116 3213 3133 3216
rect 3284 3213 3309 3216
rect 3346 3213 3380 3216
rect 3386 3213 3396 3216
rect 2020 3203 2045 3206
rect 2130 3203 2156 3206
rect 2346 3205 2349 3213
rect 2378 3203 2404 3206
rect 2498 3203 2508 3206
rect 2698 3205 2701 3213
rect 2740 3203 2765 3206
rect 2786 3203 2804 3206
rect 2914 3203 2948 3206
rect 2994 3203 3028 3206
rect 3042 3205 3045 3213
rect 38 3167 3466 3173
rect 802 3143 844 3146
rect 1082 3143 1101 3146
rect 3298 3143 3332 3146
rect 1098 3136 1101 3143
rect 210 3126 213 3134
rect 258 3133 284 3136
rect 532 3133 549 3136
rect 572 3133 613 3136
rect 642 3133 652 3136
rect 770 3133 780 3136
rect 858 3133 876 3136
rect 1034 3133 1052 3136
rect 1068 3133 1093 3136
rect 1098 3133 1116 3136
rect 1146 3133 1156 3136
rect 1522 3133 1532 3136
rect 1554 3133 1604 3136
rect 1634 3133 1652 3136
rect 1658 3133 1700 3136
rect 1754 3133 1764 3136
rect 1786 3133 1812 3136
rect 1826 3133 1852 3136
rect 1930 3133 1940 3136
rect 1964 3133 1989 3136
rect 2020 3133 2029 3136
rect 2082 3133 2100 3136
rect 2130 3133 2164 3136
rect 2234 3133 2260 3136
rect 2282 3133 2316 3136
rect 2354 3133 2364 3136
rect 2410 3133 2444 3136
rect 2450 3133 2460 3136
rect 2490 3133 2516 3136
rect 2554 3133 2596 3136
rect 2620 3133 2629 3136
rect 2724 3133 2741 3136
rect 2780 3133 2789 3136
rect 2884 3133 2892 3136
rect 2914 3133 2948 3136
rect 116 3123 141 3126
rect 172 3123 213 3126
rect 220 3123 236 3126
rect 340 3123 356 3126
rect 428 3123 444 3126
rect 586 3123 612 3126
rect 650 3123 660 3126
rect 858 3125 861 3133
rect 2786 3126 2789 3133
rect 2978 3126 2981 3134
rect 3018 3133 3044 3136
rect 3058 3133 3076 3136
rect 3090 3133 3124 3136
rect 3148 3133 3173 3136
rect 3178 3126 3181 3134
rect 3212 3133 3237 3136
rect 3260 3133 3268 3136
rect 3340 3133 3364 3136
rect 3404 3133 3421 3136
rect 946 3123 980 3126
rect 986 3123 996 3126
rect 1018 3123 1044 3126
rect 1076 3123 1117 3126
rect 1180 3123 1221 3126
rect 1260 3123 1269 3126
rect 1276 3123 1301 3126
rect 1370 3123 1388 3126
rect 1410 3123 1420 3126
rect 1660 3123 1677 3126
rect 1682 3123 1692 3126
rect 1730 3123 1756 3126
rect 1828 3123 1853 3126
rect 1882 3123 1924 3126
rect 1930 3123 1948 3126
rect 1962 3123 2004 3126
rect 2066 3123 2101 3126
rect 2188 3123 2197 3126
rect 2340 3123 2372 3126
rect 2458 3123 2468 3126
rect 2490 3123 2524 3126
rect 2556 3123 2597 3126
rect 2652 3123 2685 3126
rect 2738 3123 2756 3126
rect 2786 3123 2804 3126
rect 2810 3123 2860 3126
rect 2930 3123 2956 3126
rect 2970 3123 2981 3126
rect 2988 3123 3045 3126
rect 3052 3123 3077 3126
rect 3084 3123 3125 3126
rect 3154 3123 3181 3126
rect 3188 3123 3196 3126
rect 3218 3123 3244 3126
rect 3266 3123 3276 3126
rect 3292 3123 3333 3126
rect 3372 3123 3381 3126
rect 252 3113 277 3116
rect 308 3113 325 3116
rect 372 3113 413 3116
rect 460 3113 501 3116
rect 666 3113 708 3116
rect 898 3113 916 3116
rect 940 3113 949 3116
rect 1012 3113 1037 3116
rect 1436 3113 1477 3116
rect 714 3103 724 3106
rect 898 3103 932 3106
rect 1882 3103 1885 3123
rect 1930 3115 1933 3123
rect 2194 3116 2197 3123
rect 1964 3113 1981 3116
rect 2124 3113 2149 3116
rect 2194 3113 2204 3116
rect 2404 3113 2421 3116
rect 2484 3113 2493 3116
rect 2490 3083 2493 3113
rect 14 3067 3490 3073
rect 220 3023 237 3026
rect 492 3023 509 3026
rect 628 3023 645 3026
rect 1420 3023 1429 3026
rect 1548 3023 1581 3026
rect 2148 3023 2165 3026
rect 2892 3023 2925 3026
rect 2922 3016 2925 3023
rect 116 3013 141 3016
rect 172 3013 181 3016
rect 188 3013 204 3016
rect 276 3013 301 3016
rect 380 3013 405 3016
rect 436 3013 453 3016
rect 460 3013 476 3016
rect 498 3013 516 3016
rect 562 3013 580 3016
rect 634 3013 652 3016
rect 756 3013 773 3016
rect 178 3005 181 3013
rect 450 3005 453 3013
rect 786 3006 789 3014
rect 682 3003 692 3006
rect 754 3003 789 3006
rect 818 3006 821 3014
rect 940 3013 949 3016
rect 970 3013 980 3016
rect 1066 3006 1069 3014
rect 1138 3013 1172 3016
rect 1234 3013 1245 3016
rect 1290 3013 1316 3016
rect 1370 3013 1404 3016
rect 1418 3013 1436 3016
rect 1468 3013 1477 3016
rect 1682 3013 1692 3016
rect 1786 3013 1796 3016
rect 1874 3013 1900 3016
rect 1970 3013 2004 3016
rect 2066 3013 2076 3016
rect 2122 3013 2132 3016
rect 2234 3013 2244 3016
rect 2258 3013 2301 3016
rect 2364 3013 2413 3016
rect 2426 3013 2436 3016
rect 2442 3013 2452 3016
rect 2458 3013 2476 3016
rect 818 3003 829 3006
rect 852 3003 893 3006
rect 954 3003 972 3006
rect 1028 3003 1069 3006
rect 1146 3003 1180 3006
rect 1242 2996 1245 3013
rect 1282 3003 1308 3006
rect 1378 3003 1396 3006
rect 1466 3003 1492 3006
rect 1562 3003 1596 3006
rect 1618 3003 1636 3006
rect 1666 3003 1700 3006
rect 1722 3003 1732 3006
rect 1770 3003 1804 3006
rect 1866 3003 1908 3006
rect 2114 3003 2124 3006
rect 2154 3003 2180 3006
rect 2298 3005 2301 3013
rect 2538 3006 2541 3014
rect 2578 3013 2620 3016
rect 2740 3013 2765 3016
rect 2850 3013 2860 3016
rect 2922 3013 2957 3016
rect 2964 3013 3021 3016
rect 3042 3013 3060 3016
rect 3308 3013 3317 3016
rect 2356 3003 2373 3006
rect 2378 3003 2412 3006
rect 2458 3003 2468 3006
rect 2524 3003 2541 3006
rect 2564 3003 2573 3006
rect 2578 3003 2628 3006
rect 2892 3003 2933 3006
rect 3018 3005 3021 3013
rect 874 2993 892 2996
rect 1242 2993 1268 2996
rect 2194 2993 2212 2996
rect 2482 2993 2516 2996
rect 38 2967 3466 2973
rect 1490 2936 1493 2946
rect 106 2933 148 2936
rect 154 2933 172 2936
rect 204 2933 221 2936
rect 316 2933 333 2936
rect 106 2923 109 2933
rect 482 2926 485 2935
rect 530 2926 533 2935
rect 652 2933 677 2936
rect 722 2933 732 2936
rect 748 2933 789 2936
rect 794 2933 804 2936
rect 860 2933 892 2936
rect 908 2933 925 2936
rect 1002 2933 1012 2936
rect 1228 2933 1253 2936
rect 1386 2933 1396 2936
rect 1484 2933 1493 2936
rect 1676 2933 1685 2936
rect 1738 2933 1764 2936
rect 1820 2933 1845 2936
rect 1922 2933 1932 2936
rect 2242 2933 2252 2936
rect 2322 2933 2332 2936
rect 2426 2933 2460 2936
rect 3186 2933 3212 2936
rect 922 2927 925 2933
rect 156 2923 165 2926
rect 268 2923 284 2926
rect 396 2923 421 2926
rect 452 2923 485 2926
rect 492 2923 508 2926
rect 522 2923 533 2926
rect 682 2923 700 2926
rect 756 2923 789 2926
rect 922 2924 940 2927
rect 1842 2926 1845 2933
rect 1010 2923 1020 2926
rect 1084 2923 1109 2926
rect 1146 2923 1180 2926
rect 1194 2923 1204 2926
rect 1316 2923 1341 2926
rect 1378 2923 1404 2926
rect 1490 2923 1516 2926
rect 1538 2923 1548 2926
rect 1570 2923 1596 2926
rect 1634 2923 1652 2926
rect 1786 2923 1796 2926
rect 1842 2923 1860 2926
rect 1866 2923 1892 2926
rect 1924 2923 1933 2926
rect 1970 2923 1988 2926
rect 2020 2923 2037 2926
rect 2146 2923 2164 2926
rect 2196 2923 2205 2926
rect 2244 2923 2253 2926
rect 2260 2923 2277 2926
rect 2354 2923 2388 2926
rect 2474 2923 2500 2926
rect 2538 2923 2581 2926
rect 2676 2923 2685 2926
rect 2740 2923 2749 2926
rect 2844 2923 2853 2926
rect 3186 2925 3189 2933
rect 3194 2923 3220 2926
rect 3372 2923 3381 2926
rect 956 2913 965 2916
rect 1420 2913 1429 2916
rect 1564 2913 1589 2916
rect 1732 2913 1757 2916
rect 1956 2913 1965 2916
rect 3010 2913 3028 2916
rect 3140 2913 3149 2916
rect 930 2903 948 2906
rect 3018 2903 3044 2906
rect 3114 2903 3156 2906
rect 14 2867 3490 2873
rect 3186 2833 3204 2836
rect 892 2823 901 2826
rect 3108 2823 3141 2826
rect 3180 2823 3188 2826
rect 556 2813 581 2816
rect 612 2813 637 2816
rect 674 2813 684 2816
rect 698 2813 724 2816
rect 770 2813 788 2816
rect 794 2813 820 2816
rect 850 2813 876 2816
rect 946 2813 964 2816
rect 1140 2813 1165 2816
rect 1202 2813 1236 2816
rect 1258 2813 1292 2816
rect 1324 2813 1357 2816
rect 1452 2813 1469 2816
rect 1500 2813 1517 2816
rect 1556 2813 1565 2816
rect 1700 2813 1725 2816
rect 1756 2813 1765 2816
rect 1828 2813 1853 2816
rect 1972 2813 1989 2816
rect 2034 2813 2052 2816
rect 2066 2813 2084 2816
rect 2140 2813 2165 2816
rect 2234 2813 2252 2816
rect 2378 2813 2396 2816
rect 2410 2813 2428 2816
rect 2596 2813 2605 2816
rect 2668 2813 2677 2816
rect 2730 2813 2740 2816
rect 2834 2813 2844 2816
rect 2874 2813 2884 2816
rect 2972 2813 2980 2816
rect 3106 2813 3172 2816
rect 3276 2813 3293 2816
rect 770 2806 773 2813
rect 428 2803 437 2806
rect 442 2803 452 2806
rect 458 2803 476 2806
rect 618 2803 644 2806
rect 748 2803 773 2806
rect 802 2803 812 2806
rect 858 2803 868 2806
rect 970 2803 1020 2806
rect 1210 2803 1228 2806
rect 1266 2803 1284 2806
rect 1466 2805 1469 2813
rect 1618 2803 1636 2806
rect 1762 2805 1765 2813
rect 2370 2803 2388 2806
rect 2570 2803 2588 2806
rect 2602 2803 2620 2806
rect 2660 2803 2685 2806
rect 2722 2803 2732 2806
rect 2802 2803 2820 2806
rect 2826 2803 2836 2806
rect 3108 2803 3117 2806
rect 3218 2803 3268 2806
rect 402 2793 420 2796
rect 898 2793 924 2796
rect 2698 2793 2708 2796
rect 3290 2795 3293 2813
rect 3300 2803 3317 2806
rect 38 2767 3466 2773
rect 506 2743 540 2746
rect 1082 2743 1100 2746
rect 1138 2743 1165 2746
rect 1402 2743 1436 2746
rect 1450 2743 1460 2746
rect 602 2733 628 2736
rect 634 2733 660 2736
rect 834 2733 860 2736
rect 1050 2726 1053 2735
rect 1066 2733 1076 2736
rect 1108 2733 1141 2736
rect 1146 2733 1180 2736
rect 1402 2733 1444 2736
rect 1468 2733 1485 2736
rect 1532 2733 1573 2736
rect 1706 2726 1709 2735
rect 1722 2726 1725 2745
rect 1802 2743 1828 2746
rect 1836 2733 1861 2736
rect 1882 2726 1885 2745
rect 2026 2726 2029 2745
rect 2978 2743 2996 2746
rect 2036 2733 2053 2736
rect 2060 2733 2101 2736
rect 2228 2733 2253 2736
rect 2354 2733 2388 2736
rect 2978 2733 3004 2736
rect 3226 2733 3260 2736
rect 3274 2733 3284 2736
rect 164 2723 173 2726
rect 324 2723 349 2726
rect 380 2723 405 2726
rect 572 2723 613 2726
rect 642 2723 668 2726
rect 684 2723 709 2726
rect 764 2723 789 2726
rect 820 2723 853 2726
rect 964 2723 981 2726
rect 1020 2723 1053 2726
rect 1084 2723 1093 2726
rect 1194 2723 1204 2726
rect 1268 2723 1277 2726
rect 1452 2723 1461 2726
rect 1498 2723 1516 2726
rect 1612 2723 1637 2726
rect 1668 2723 1709 2726
rect 1716 2723 1725 2726
rect 1762 2723 1796 2726
rect 1876 2723 1885 2726
rect 1988 2723 2029 2726
rect 2292 2723 2317 2726
rect 2444 2723 2469 2726
rect 2564 2723 2573 2726
rect 2620 2723 2637 2726
rect 2676 2723 2685 2726
rect 2796 2723 2805 2726
rect 2916 2723 2941 2726
rect 3132 2723 3141 2726
rect 3146 2723 3172 2726
rect 3186 2723 3253 2726
rect 3268 2723 3285 2726
rect 3364 2723 3389 2726
rect 14 2667 3490 2673
rect 3058 2636 3061 2646
rect 3018 2633 3037 2636
rect 3058 2633 3092 2636
rect 116 2613 149 2616
rect 188 2613 221 2616
rect 226 2606 229 2614
rect 260 2613 277 2616
rect 282 2613 292 2616
rect 324 2613 357 2616
rect 396 2613 405 2616
rect 516 2613 533 2616
rect 538 2613 548 2616
rect 596 2613 605 2616
rect 812 2613 837 2616
rect 924 2613 941 2616
rect 1028 2613 1045 2616
rect 1196 2613 1213 2616
rect 1356 2613 1381 2616
rect 1412 2613 1429 2616
rect 1468 2613 1485 2616
rect 1524 2613 1533 2616
rect 1628 2613 1645 2616
rect 1780 2613 1805 2616
rect 1836 2613 1845 2616
rect 1940 2613 1949 2616
rect 2154 2613 2164 2616
rect 2244 2613 2253 2616
rect 2300 2613 2317 2616
rect 2436 2613 2477 2616
rect 2524 2613 2565 2616
rect 2572 2613 2597 2616
rect 2852 2613 2877 2616
rect 2924 2613 2949 2616
rect 3034 2615 3037 2633
rect 3058 2623 3076 2626
rect 3114 2613 3156 2616
rect 3172 2613 3229 2616
rect 108 2603 141 2606
rect 146 2603 164 2606
rect 202 2603 229 2606
rect 322 2603 372 2606
rect 522 2603 540 2606
rect 2380 2603 2397 2606
rect 2434 2603 2500 2606
rect 2522 2603 2564 2606
rect 2578 2603 2612 2606
rect 2778 2603 2828 2606
rect 146 2596 149 2603
rect 122 2593 149 2596
rect 3114 2593 3117 2613
rect 3138 2603 3148 2606
rect 3178 2603 3228 2606
rect 3266 2603 3316 2606
rect 3332 2603 3357 2606
rect 3362 2603 3396 2606
rect 3362 2593 3365 2603
rect 38 2567 3466 2573
rect 554 2543 573 2546
rect 554 2536 557 2543
rect 1842 2536 1845 2546
rect 3034 2543 3068 2546
rect 410 2533 436 2536
rect 458 2533 524 2536
rect 540 2533 557 2536
rect 562 2533 620 2536
rect 706 2533 716 2536
rect 826 2533 861 2536
rect 884 2533 917 2536
rect 1026 2533 1044 2536
rect 1202 2533 1212 2536
rect 1250 2533 1260 2536
rect 1276 2533 1293 2536
rect 1554 2533 1572 2536
rect 1610 2533 1620 2536
rect 1666 2533 1700 2536
rect 1746 2533 1796 2536
rect 1818 2533 1845 2536
rect 1914 2533 1949 2536
rect 164 2523 189 2526
rect 324 2523 349 2526
rect 460 2523 493 2526
rect 740 2523 749 2526
rect 826 2525 829 2533
rect 892 2523 925 2526
rect 964 2523 981 2526
rect 1020 2523 1036 2526
rect 1068 2523 1085 2526
rect 1124 2523 1141 2526
rect 1180 2523 1197 2526
rect 1242 2523 1252 2526
rect 1284 2523 1301 2526
rect 1340 2523 1365 2526
rect 1396 2523 1404 2526
rect 1548 2523 1564 2526
rect 1602 2523 1612 2526
rect 1818 2525 1821 2533
rect 1914 2525 1917 2533
rect 1922 2523 1956 2526
rect 2002 2523 2012 2526
rect 2042 2525 2045 2536
rect 2050 2533 2100 2536
rect 2122 2533 2149 2536
rect 2186 2533 2196 2536
rect 2322 2533 2356 2536
rect 2554 2533 2588 2536
rect 2644 2533 2700 2536
rect 2730 2533 2788 2536
rect 2810 2533 2868 2536
rect 3226 2533 3244 2536
rect 2082 2523 2092 2526
rect 2122 2525 2125 2533
rect 3274 2526 3277 2545
rect 3284 2533 3309 2536
rect 2178 2523 2188 2526
rect 2220 2523 2269 2526
rect 2386 2523 2412 2526
rect 2474 2523 2484 2526
rect 2554 2523 2604 2526
rect 2724 2523 2765 2526
rect 2812 2523 2853 2526
rect 2892 2523 2933 2526
rect 2972 2523 2989 2526
rect 3028 2523 3061 2526
rect 3154 2523 3180 2526
rect 3218 2523 3252 2526
rect 3266 2523 3277 2526
rect 3114 2513 3124 2516
rect 3148 2513 3165 2516
rect 3196 2513 3237 2516
rect 3266 2515 3269 2523
rect 3098 2503 3140 2506
rect 14 2467 3490 2473
rect 1028 2423 1037 2426
rect 1092 2423 1117 2426
rect 1340 2423 1357 2426
rect 124 2413 133 2416
rect 180 2413 205 2416
rect 244 2413 269 2416
rect 356 2413 381 2416
rect 412 2413 429 2416
rect 468 2413 493 2416
rect 580 2413 605 2416
rect 692 2413 709 2416
rect 916 2413 941 2416
rect 1042 2413 1076 2416
rect 1228 2413 1253 2416
rect 1290 2413 1324 2416
rect 1564 2413 1581 2416
rect 1620 2413 1645 2416
rect 1676 2413 1693 2416
rect 1732 2413 1757 2416
rect 1836 2413 1861 2416
rect 1932 2413 1957 2416
rect 2028 2413 2053 2416
rect 2220 2413 2245 2416
rect 2316 2413 2325 2416
rect 2412 2413 2437 2416
rect 2604 2413 2629 2416
rect 2700 2413 2717 2416
rect 2796 2413 2821 2416
rect 2988 2413 2997 2416
rect 3084 2413 3093 2416
rect 3236 2413 3245 2416
rect 3292 2413 3317 2416
rect 3362 2415 3365 2426
rect 3388 2423 3397 2426
rect 3412 2423 3429 2426
rect 978 2403 1004 2406
rect 1042 2403 1068 2406
rect 1098 2403 1124 2406
rect 1394 2403 1420 2406
rect 1444 2403 1469 2406
rect 3242 2405 3245 2413
rect 38 2367 3466 2373
rect 202 2333 220 2336
rect 244 2333 253 2336
rect 298 2333 340 2336
rect 378 2333 396 2336
rect 426 2333 468 2336
rect 556 2333 565 2336
rect 570 2333 596 2336
rect 620 2333 653 2336
rect 658 2326 661 2335
rect 674 2333 700 2336
rect 738 2333 772 2336
rect 852 2333 893 2336
rect 986 2333 996 2336
rect 1018 2326 1021 2335
rect 1026 2333 1036 2336
rect 1106 2326 1109 2335
rect 1114 2333 1132 2336
rect 1162 2333 1204 2336
rect 1226 2326 1229 2335
rect 1268 2333 1277 2336
rect 1378 2333 1436 2336
rect 1492 2333 1509 2336
rect 1564 2333 1573 2336
rect 1786 2333 1804 2336
rect 1842 2333 1868 2336
rect 1898 2333 1932 2336
rect 1956 2333 1981 2336
rect 2018 2333 2060 2336
rect 2084 2333 2109 2336
rect 2114 2326 2117 2335
rect 2204 2333 2237 2336
rect 2388 2333 2413 2336
rect 2458 2333 2484 2336
rect 2564 2333 2589 2336
rect 2802 2333 2820 2336
rect 2850 2333 2868 2336
rect 2898 2333 2948 2336
rect 2962 2333 2972 2336
rect 3026 2333 3044 2336
rect 3140 2333 3156 2336
rect 3170 2333 3236 2336
rect 3250 2333 3316 2336
rect 3346 2333 3364 2336
rect 3388 2333 3396 2336
rect 116 2323 125 2326
rect 172 2323 181 2326
rect 242 2323 268 2326
rect 562 2323 604 2326
rect 634 2323 661 2326
rect 668 2323 693 2326
rect 698 2323 708 2326
rect 730 2323 780 2326
rect 810 2323 836 2326
rect 850 2323 908 2326
rect 1018 2323 1029 2326
rect 1044 2323 1085 2326
rect 1106 2323 1125 2326
rect 1154 2323 1212 2326
rect 1226 2323 1252 2326
rect 1338 2323 1356 2326
rect 1370 2323 1444 2326
rect 1490 2323 1548 2326
rect 1578 2323 1596 2326
rect 1634 2323 1652 2326
rect 1674 2323 1684 2326
rect 1794 2323 1812 2326
rect 1842 2323 1876 2326
rect 2058 2323 2068 2326
rect 2082 2323 2117 2326
rect 492 2313 525 2316
rect 620 2313 645 2316
rect 724 2313 765 2316
rect 796 2313 821 2316
rect 1026 2283 1029 2323
rect 1372 2313 1429 2316
rect 1492 2313 1525 2316
rect 1612 2313 1621 2316
rect 1892 2313 1925 2316
rect 2140 2313 2157 2316
rect 2204 2313 2229 2316
rect 2234 2313 2237 2333
rect 2282 2323 2308 2326
rect 2362 2323 2372 2326
rect 2394 2323 2428 2326
rect 2450 2323 2492 2326
rect 2530 2323 2548 2326
rect 2730 2323 2756 2326
rect 2794 2323 2828 2326
rect 2842 2323 2876 2326
rect 2956 2323 2973 2326
rect 3148 2323 3157 2326
rect 3210 2323 3244 2326
rect 2324 2313 2357 2316
rect 2724 2313 2741 2316
rect 2772 2313 2781 2316
rect 2844 2313 2861 2316
rect 2996 2313 3037 2316
rect 3172 2313 3221 2316
rect 3250 2315 3253 2333
rect 3276 2323 3285 2326
rect 3362 2323 3372 2326
rect 3386 2323 3397 2326
rect 3404 2323 3429 2326
rect 3340 2313 3357 2316
rect 3386 2315 3389 2323
rect 1426 2303 1429 2313
rect 1618 2303 1621 2313
rect 14 2267 3490 2273
rect 2058 2253 2077 2256
rect 116 2223 149 2226
rect 324 2223 357 2226
rect 532 2223 573 2226
rect 1180 2223 1189 2226
rect 1804 2223 1821 2226
rect 354 2216 357 2223
rect 1938 2216 1941 2236
rect 2268 2223 2277 2226
rect 2676 2223 2693 2226
rect 2884 2223 2893 2226
rect 2996 2223 3005 2226
rect 3036 2223 3045 2226
rect 2890 2216 2893 2223
rect 66 2213 100 2216
rect 114 2213 164 2216
rect 178 2213 197 2216
rect 210 2213 236 2216
rect 194 2206 197 2213
rect 274 2206 277 2216
rect 316 2213 349 2216
rect 354 2213 365 2216
rect 386 2213 428 2216
rect 474 2213 492 2216
rect 524 2213 533 2216
rect 538 2213 580 2216
rect 626 2213 660 2216
rect 684 2213 701 2216
rect 714 2213 724 2216
rect 762 2213 796 2216
rect 802 2213 845 2216
rect 900 2213 932 2216
rect 964 2213 1013 2216
rect 1052 2213 1069 2216
rect 1074 2213 1100 2216
rect 1250 2213 1292 2216
rect 1340 2213 1357 2216
rect 1450 2213 1468 2216
rect 1556 2213 1565 2216
rect 1578 2213 1596 2216
rect 1634 2213 1644 2216
rect 1700 2213 1717 2216
rect 346 2206 349 2213
rect 1762 2206 1765 2216
rect 1778 2213 1796 2216
rect 1818 2213 1836 2216
rect 1858 2213 1900 2216
rect 1938 2213 1964 2216
rect 2092 2213 2109 2216
rect 2156 2213 2165 2216
rect 2170 2213 2204 2216
rect 2242 2213 2260 2216
rect 2274 2213 2316 2216
rect 2378 2213 2428 2216
rect 2442 2213 2451 2216
rect 2538 2213 2556 2216
rect 2562 2213 2596 2216
rect 2634 2213 2660 2216
rect 2682 2213 2716 2216
rect 2746 2213 2772 2216
rect 116 2203 125 2206
rect 130 2203 156 2206
rect 180 2203 189 2206
rect 194 2203 244 2206
rect 274 2203 308 2206
rect 346 2203 364 2206
rect 388 2203 413 2206
rect 604 2203 652 2206
rect 722 2203 732 2206
rect 748 2203 781 2206
rect 810 2203 828 2206
rect 858 2203 876 2206
rect 1058 2203 1085 2206
rect 1130 2203 1156 2206
rect 1180 2203 1189 2206
rect 1194 2203 1219 2206
rect 1266 2203 1284 2206
rect 1362 2203 1372 2206
rect 1442 2203 1460 2206
rect 1524 2203 1533 2206
rect 1548 2203 1597 2206
rect 1626 2203 1636 2206
rect 1650 2203 1692 2206
rect 1762 2203 1788 2206
rect 1802 2203 1828 2206
rect 1852 2203 1893 2206
rect 1970 2203 2020 2206
rect 2148 2203 2197 2206
rect 2202 2203 2212 2206
rect 2306 2203 2324 2206
rect 2634 2203 2652 2206
rect 2690 2203 2708 2206
rect 2732 2203 2741 2206
rect 2754 2203 2764 2206
rect 2786 2205 2789 2216
rect 2890 2213 2901 2216
rect 2994 2213 3020 2216
rect 3034 2213 3084 2216
rect 3098 2213 3108 2216
rect 3138 2213 3172 2216
rect 3322 2213 3340 2216
rect 3420 2213 3429 2216
rect 2812 2203 2821 2206
rect 2884 2203 2893 2206
rect 2924 2203 2933 2206
rect 2938 2203 2972 2206
rect 3058 2203 3076 2206
rect 3124 2203 3133 2206
rect 3362 2203 3412 2206
rect 1338 2193 1364 2196
rect 1506 2193 1516 2196
rect 2690 2193 2693 2203
rect 3178 2193 3196 2196
rect 3370 2193 3404 2196
rect 38 2167 3466 2173
rect 826 2143 852 2146
rect 914 2143 924 2146
rect 970 2143 997 2146
rect 970 2136 973 2143
rect 204 2133 237 2136
rect 274 2133 285 2136
rect 306 2133 316 2136
rect 372 2133 389 2136
rect 410 2133 428 2136
rect 676 2133 685 2136
rect 690 2133 708 2136
rect 746 2133 764 2136
rect 778 2133 788 2136
rect 850 2133 860 2136
rect 866 2133 876 2136
rect 956 2133 973 2136
rect 978 2133 1012 2136
rect 282 2126 285 2133
rect 1042 2126 1045 2146
rect 124 2123 165 2126
rect 218 2123 244 2126
rect 282 2123 324 2126
rect 338 2123 348 2126
rect 452 2123 469 2126
rect 522 2123 540 2126
rect 546 2123 580 2126
rect 626 2123 652 2126
rect 684 2123 693 2126
rect 716 2123 725 2126
rect 738 2123 772 2126
rect 796 2123 821 2126
rect 868 2123 884 2126
rect 964 2123 973 2126
rect 1036 2123 1045 2126
rect 1050 2123 1053 2156
rect 1634 2143 1644 2146
rect 1740 2143 1749 2146
rect 2994 2143 3005 2146
rect 2994 2136 2997 2143
rect 1100 2133 1109 2136
rect 1154 2133 1164 2136
rect 1188 2133 1197 2136
rect 1218 2133 1236 2136
rect 1284 2133 1301 2136
rect 1306 2133 1324 2136
rect 1386 2133 1436 2136
rect 1474 2133 1508 2136
rect 1524 2133 1541 2136
rect 1652 2133 1661 2136
rect 1738 2133 1772 2136
rect 1810 2133 1821 2136
rect 1850 2133 1900 2136
rect 1810 2126 1813 2133
rect 1058 2123 1084 2126
rect 1162 2123 1172 2126
rect 1252 2123 1261 2126
rect 1388 2123 1405 2126
rect 1426 2123 1444 2126
rect 1490 2123 1500 2126
rect 1546 2123 1580 2126
rect 1660 2123 1676 2126
rect 1740 2123 1749 2126
rect 1780 2123 1813 2126
rect 1874 2123 1908 2126
rect 332 2113 341 2116
rect 466 2113 492 2116
rect 724 2113 765 2116
rect 780 2113 789 2116
rect 458 2103 508 2106
rect 1930 2103 1933 2134
rect 2012 2133 2061 2136
rect 2130 2133 2140 2136
rect 2156 2133 2165 2136
rect 2218 2133 2252 2136
rect 2268 2133 2317 2136
rect 2338 2133 2356 2136
rect 2372 2133 2413 2136
rect 2474 2133 2500 2136
rect 2538 2133 2556 2136
rect 2692 2133 2741 2136
rect 2794 2133 2820 2136
rect 2850 2133 2860 2136
rect 2964 2133 2997 2136
rect 3002 2133 3012 2136
rect 3162 2133 3180 2136
rect 1962 2123 1988 2126
rect 2164 2123 2189 2126
rect 2194 2123 2212 2126
rect 2218 2123 2221 2133
rect 3226 2126 3229 2156
rect 3266 2133 3292 2136
rect 3298 2133 3316 2136
rect 3370 2133 3380 2136
rect 2234 2116 2237 2126
rect 2298 2123 2332 2126
rect 2338 2123 2348 2126
rect 2394 2123 2428 2126
rect 2458 2123 2468 2126
rect 2498 2123 2508 2126
rect 2594 2123 2636 2126
rect 2706 2123 2740 2126
rect 2778 2123 2788 2126
rect 2828 2123 2861 2126
rect 3010 2123 3020 2126
rect 3034 2123 3051 2126
rect 3114 2123 3124 2126
rect 3226 2123 3244 2126
rect 3260 2123 3285 2126
rect 3338 2123 3364 2126
rect 1948 2113 1981 2116
rect 2092 2113 2117 2116
rect 2220 2113 2237 2116
rect 2524 2113 2549 2116
rect 2836 2113 2845 2116
rect 14 2067 3490 2073
rect 66 2043 85 2046
rect 338 2033 356 2036
rect 442 2026 445 2036
rect 458 2033 476 2036
rect 164 2023 189 2026
rect 260 2023 301 2026
rect 316 2023 333 2026
rect 340 2023 349 2026
rect 364 2023 389 2026
rect 442 2023 460 2026
rect 532 2023 549 2026
rect 836 2023 845 2026
rect 1108 2023 1117 2026
rect 1706 2016 1709 2036
rect 1962 2033 1996 2036
rect 2410 2033 2420 2036
rect 2442 2033 2476 2036
rect 1900 2023 1917 2026
rect 1954 2023 1980 2026
rect 2004 2023 2021 2026
rect 2186 2023 2221 2026
rect 2450 2023 2460 2026
rect 2524 2023 2557 2026
rect 156 2013 197 2016
rect 234 2013 244 2016
rect 266 2013 308 2016
rect 378 2013 404 2016
rect 490 2013 524 2016
rect 580 2013 605 2016
rect 676 2013 692 2016
rect 748 2013 773 2016
rect 812 2013 821 2016
rect 1010 2013 1028 2016
rect 218 2003 236 2006
rect 260 2003 293 2006
rect 498 2003 516 2006
rect 538 2003 556 2006
rect 586 2003 620 2006
rect 804 2003 821 2006
rect 922 2003 932 2006
rect 948 2003 973 2006
rect 1018 2003 1036 2006
rect 1052 2003 1085 2006
rect 1090 2005 1093 2016
rect 1100 2013 1125 2016
rect 1234 2013 1243 2016
rect 1276 2013 1309 2016
rect 1370 2013 1380 2016
rect 1386 2013 1436 2016
rect 1482 2013 1516 2016
rect 1564 2013 1573 2016
rect 1580 2013 1605 2016
rect 1610 2006 1613 2015
rect 1644 2013 1653 2016
rect 1698 2013 1709 2016
rect 1754 2006 1757 2015
rect 1762 2013 1804 2016
rect 1850 2013 1860 2016
rect 1892 2013 1909 2016
rect 1914 2006 1917 2023
rect 2060 2013 2093 2016
rect 2242 2013 2260 2016
rect 2292 2013 2324 2016
rect 2348 2013 2357 2016
rect 2498 2013 2516 2016
rect 2546 2013 2564 2016
rect 2570 2006 2573 2025
rect 2596 2023 2605 2026
rect 2668 2023 2677 2026
rect 2828 2023 2845 2026
rect 3020 2023 3037 2026
rect 3156 2023 3181 2026
rect 2594 2013 2660 2016
rect 2738 2013 2756 2016
rect 2826 2013 2868 2016
rect 2906 2013 2925 2016
rect 2970 2013 3004 2016
rect 3058 2013 3076 2016
rect 3106 2013 3140 2016
rect 3234 2013 3244 2016
rect 3250 2013 3293 2016
rect 1106 2003 1140 2006
rect 1186 2003 1204 2006
rect 1234 2003 1245 2006
rect 1314 2003 1324 2006
rect 1356 2003 1372 2006
rect 1386 2003 1428 2006
rect 1452 2003 1461 2006
rect 1474 2003 1508 2006
rect 1530 2003 1540 2006
rect 1602 2003 1613 2006
rect 1650 2003 1676 2006
rect 1700 2003 1725 2006
rect 1754 2003 1773 2006
rect 1802 2003 1812 2006
rect 1828 2003 1845 2006
rect 1906 2003 1917 2006
rect 2018 2003 2028 2006
rect 2042 2003 2052 2006
rect 2138 2003 2148 2006
rect 2164 2003 2205 2006
rect 2242 2003 2268 2006
rect 2284 2003 2309 2006
rect 2522 2003 2556 2006
rect 2570 2003 2580 2006
rect 2618 2003 2652 2006
rect 2714 2003 2748 2006
rect 2842 2003 2860 2006
rect 2884 2003 2909 2006
rect 2922 2005 2925 2013
rect 3290 2006 3293 2013
rect 3042 2003 3068 2006
rect 3100 2003 3109 2006
rect 3114 2003 3132 2006
rect 3156 2003 3173 2006
rect 3282 2005 3293 2006
rect 3282 2003 3292 2005
rect 3306 2003 3324 2006
rect 1234 1996 1237 2003
rect 1220 1993 1237 1996
rect 1282 1993 1316 1996
rect 1338 1993 1348 1996
rect 1386 1993 1389 2003
rect 1458 1995 1461 2003
rect 3106 1983 3109 2003
rect 3186 1993 3204 1996
rect 38 1967 3466 1973
rect 82 1933 92 1936
rect 196 1933 229 1936
rect 106 1923 116 1926
rect 138 1923 172 1926
rect 204 1923 229 1926
rect 242 1925 245 1956
rect 978 1953 1005 1956
rect 386 1943 397 1946
rect 394 1936 397 1943
rect 338 1933 356 1936
rect 372 1933 389 1936
rect 394 1933 420 1936
rect 442 1933 484 1936
rect 538 1933 564 1936
rect 580 1933 605 1936
rect 658 1933 676 1936
rect 746 1933 780 1936
rect 866 1933 884 1936
rect 930 1933 948 1936
rect 964 1933 997 1936
rect 124 1913 149 1916
rect 226 1913 229 1923
rect 266 1906 269 1926
rect 338 1916 341 1933
rect 1002 1926 1005 1953
rect 1506 1943 1533 1946
rect 3178 1943 3188 1946
rect 3242 1943 3268 1946
rect 1506 1936 1509 1943
rect 1036 1933 1061 1936
rect 1082 1933 1124 1936
rect 1138 1933 1156 1936
rect 1228 1933 1236 1936
rect 1324 1933 1341 1936
rect 1450 1933 1460 1936
rect 1476 1933 1509 1936
rect 1514 1933 1540 1936
rect 1666 1933 1676 1936
rect 1692 1933 1725 1936
rect 1770 1933 1780 1936
rect 1842 1933 1876 1936
rect 1898 1933 1925 1936
rect 2026 1933 2036 1936
rect 2066 1933 2076 1936
rect 2162 1933 2180 1936
rect 2196 1933 2237 1936
rect 2298 1933 2316 1936
rect 2362 1933 2372 1936
rect 2420 1933 2429 1936
rect 2500 1933 2525 1936
rect 444 1923 461 1926
rect 492 1923 501 1926
rect 588 1923 613 1926
rect 706 1923 724 1926
rect 754 1923 772 1926
rect 796 1923 821 1926
rect 866 1923 892 1926
rect 914 1923 940 1926
rect 986 1923 1012 1926
rect 1122 1923 1132 1926
rect 1194 1923 1212 1926
rect 1226 1923 1244 1926
rect 1258 1923 1300 1926
rect 1442 1923 1452 1926
rect 1484 1923 1548 1926
rect 1554 1923 1564 1926
rect 1634 1923 1660 1926
rect 1714 1923 1748 1926
rect 1754 1923 1773 1926
rect 1820 1923 1829 1926
rect 316 1913 341 1916
rect 740 1913 765 1916
rect 210 1903 252 1906
rect 266 1903 308 1906
rect 858 1883 861 1906
rect 986 1883 989 1923
rect 1842 1916 1845 1933
rect 1898 1925 1901 1933
rect 2562 1926 2565 1936
rect 2578 1933 2588 1936
rect 2636 1933 2661 1936
rect 2714 1933 2724 1936
rect 2746 1933 2756 1936
rect 2786 1933 2796 1936
rect 2810 1933 2820 1936
rect 2866 1933 2876 1936
rect 2996 1933 3005 1936
rect 1906 1923 1940 1926
rect 2138 1923 2156 1926
rect 2210 1923 2252 1926
rect 2306 1923 2324 1926
rect 2380 1923 2389 1926
rect 2466 1923 2476 1926
rect 2562 1923 2596 1926
rect 1084 1913 1125 1916
rect 1364 1913 1373 1916
rect 1412 1913 1421 1916
rect 1842 1913 1861 1916
rect 1370 1893 1373 1913
rect 1378 1903 1428 1906
rect 1498 1903 1509 1906
rect 1970 1903 1973 1915
rect 2268 1913 2277 1916
rect 2292 1913 2301 1916
rect 2532 1913 2541 1916
rect 2658 1906 2661 1933
rect 2746 1926 2749 1933
rect 3010 1926 3013 1934
rect 3042 1933 3084 1936
rect 3108 1933 3117 1936
rect 3130 1933 3148 1936
rect 3154 1933 3196 1936
rect 3226 1933 3276 1936
rect 3300 1933 3317 1936
rect 2698 1923 2749 1926
rect 2786 1923 2804 1926
rect 2818 1923 2828 1926
rect 2850 1923 2884 1926
rect 2924 1923 2957 1926
rect 2962 1923 2980 1926
rect 2994 1923 3013 1926
rect 3066 1923 3092 1926
rect 3156 1923 3197 1926
rect 3372 1923 3397 1926
rect 3228 1913 3261 1916
rect 1978 1903 1988 1906
rect 2522 1903 2548 1906
rect 2658 1903 2684 1906
rect 1498 1893 1501 1903
rect 2522 1893 2525 1903
rect 14 1867 3490 1873
rect 1498 1833 1509 1836
rect 1770 1833 1780 1836
rect 124 1823 149 1826
rect 244 1823 253 1826
rect 300 1823 325 1826
rect 362 1823 381 1826
rect 802 1823 821 1826
rect 916 1823 925 1826
rect 362 1816 365 1823
rect 818 1816 821 1823
rect 266 1813 292 1816
rect 332 1813 365 1816
rect 378 1813 388 1816
rect 420 1813 429 1816
rect 500 1813 541 1816
rect 580 1813 613 1816
rect 634 1813 676 1816
rect 764 1813 781 1816
rect 796 1813 813 1816
rect 818 1813 844 1816
rect 890 1813 900 1816
rect 978 1813 1012 1816
rect 1044 1813 1053 1816
rect 1154 1813 1164 1816
rect 1234 1813 1245 1816
rect 1252 1813 1285 1816
rect 1316 1813 1341 1816
rect 1348 1813 1356 1816
rect 362 1806 365 1813
rect 124 1803 149 1806
rect 164 1803 205 1806
rect 210 1803 220 1806
rect 244 1803 277 1806
rect 298 1803 324 1806
rect 362 1803 396 1806
rect 412 1803 453 1806
rect 458 1803 476 1806
rect 498 1803 556 1806
rect 572 1803 605 1806
rect 636 1803 684 1806
rect 700 1803 733 1806
rect 146 1796 149 1803
rect 146 1793 156 1796
rect 778 1795 781 1813
rect 866 1803 876 1806
rect 986 1803 1020 1806
rect 1036 1803 1045 1806
rect 1140 1803 1149 1806
rect 1234 1805 1237 1813
rect 1266 1803 1300 1806
rect 1330 1803 1340 1806
rect 1410 1803 1428 1806
rect 1490 1803 1493 1815
rect 1506 1806 1509 1833
rect 1618 1823 1637 1826
rect 1514 1813 1540 1816
rect 1612 1813 1629 1816
rect 1634 1806 1637 1823
rect 1810 1816 1813 1836
rect 1858 1816 1861 1836
rect 1722 1813 1732 1816
rect 1810 1813 1820 1816
rect 1852 1813 1861 1816
rect 1866 1833 1900 1836
rect 2434 1833 2468 1836
rect 1866 1806 1869 1833
rect 1874 1823 1884 1826
rect 1964 1823 1973 1826
rect 2274 1823 2285 1826
rect 2282 1816 2285 1823
rect 1930 1813 1956 1816
rect 1994 1813 2036 1816
rect 2122 1813 2148 1816
rect 2186 1813 2228 1816
rect 2260 1813 2277 1816
rect 2282 1813 2292 1816
rect 2330 1813 2372 1816
rect 2402 1813 2420 1816
rect 2434 1813 2437 1833
rect 2594 1816 2597 1826
rect 3060 1823 3069 1826
rect 2482 1813 2532 1816
rect 2546 1813 2564 1816
rect 2594 1813 2612 1816
rect 2666 1813 2692 1816
rect 2916 1813 2949 1816
rect 2994 1813 3037 1816
rect 3074 1813 3092 1816
rect 2330 1806 2333 1813
rect 1506 1803 1517 1806
rect 1570 1803 1588 1806
rect 1634 1803 1660 1806
rect 1818 1803 1828 1806
rect 1858 1803 1869 1806
rect 1938 1803 1948 1806
rect 2146 1803 2156 1806
rect 2194 1803 2236 1806
rect 2252 1803 2285 1806
rect 2316 1803 2333 1806
rect 2570 1803 2604 1806
rect 2636 1803 2677 1806
rect 2708 1803 2725 1806
rect 2780 1803 2821 1806
rect 2882 1803 2908 1806
rect 2922 1803 2964 1806
rect 2980 1803 3005 1806
rect 3026 1803 3036 1806
rect 3060 1803 3069 1806
rect 1282 1793 1292 1796
rect 2570 1793 2573 1803
rect 3074 1786 3077 1813
rect 3194 1806 3197 1815
rect 3170 1803 3188 1806
rect 3194 1803 3252 1806
rect 3258 1796 3261 1815
rect 3306 1806 3309 1815
rect 3314 1813 3324 1816
rect 3282 1803 3300 1806
rect 3306 1803 3316 1806
rect 3258 1793 3292 1796
rect 434 1783 453 1786
rect 3066 1783 3077 1786
rect 38 1767 3466 1773
rect 74 1743 85 1746
rect 130 1743 141 1746
rect 866 1743 876 1746
rect 970 1743 1020 1746
rect 1156 1743 1181 1746
rect 74 1726 77 1743
rect 138 1736 141 1743
rect 1178 1736 1181 1743
rect 82 1733 100 1736
rect 116 1733 133 1736
rect 138 1733 180 1736
rect 194 1733 204 1736
rect 266 1733 284 1736
rect 298 1733 308 1736
rect 386 1733 396 1736
rect 410 1733 445 1736
rect 74 1723 92 1726
rect 124 1723 141 1726
rect 162 1723 188 1726
rect 218 1723 245 1726
rect 346 1723 380 1726
rect 404 1723 429 1726
rect 442 1716 445 1733
rect 634 1733 668 1736
rect 682 1733 715 1736
rect 786 1733 820 1736
rect 898 1733 940 1736
rect 956 1733 981 1736
rect 1058 1733 1092 1736
rect 1178 1733 1188 1736
rect 1218 1733 1252 1736
rect 1314 1733 1323 1736
rect 1348 1733 1357 1736
rect 1604 1733 1613 1736
rect 1636 1733 1653 1736
rect 490 1723 516 1726
rect 634 1723 637 1733
rect 1690 1726 1693 1734
rect 1698 1733 1716 1736
rect 1746 1733 1764 1736
rect 1836 1733 1877 1736
rect 2170 1733 2220 1736
rect 2236 1733 2245 1736
rect 2426 1733 2444 1736
rect 2458 1733 2468 1736
rect 2594 1733 2636 1736
rect 2754 1733 2772 1736
rect 2794 1733 2804 1736
rect 2860 1733 2885 1736
rect 2930 1733 2956 1736
rect 3036 1733 3076 1736
rect 3194 1733 3220 1736
rect 3300 1733 3325 1736
rect 1874 1726 1877 1733
rect 2594 1726 2597 1733
rect 706 1723 724 1726
rect 746 1723 780 1726
rect 892 1723 932 1726
rect 964 1723 1021 1726
rect 1100 1723 1117 1726
rect 1156 1723 1173 1726
rect 1186 1723 1196 1726
rect 412 1713 437 1716
rect 442 1713 452 1716
rect 476 1713 501 1716
rect 594 1713 604 1716
rect 706 1713 709 1723
rect 1348 1713 1357 1716
rect 434 1703 437 1713
rect 1394 1706 1397 1725
rect 1412 1713 1437 1716
rect 1458 1706 1461 1725
rect 1482 1723 1516 1726
rect 1570 1723 1588 1726
rect 1602 1723 1620 1726
rect 1650 1723 1676 1726
rect 1690 1723 1701 1726
rect 1740 1723 1765 1726
rect 1772 1723 1781 1726
rect 1794 1723 1812 1726
rect 1874 1723 1892 1726
rect 1994 1723 2012 1726
rect 2044 1723 2053 1726
rect 2092 1723 2109 1726
rect 2114 1723 2132 1726
rect 2146 1723 2212 1726
rect 2244 1723 2301 1726
rect 2306 1723 2316 1726
rect 2348 1723 2357 1726
rect 2370 1723 2388 1726
rect 2420 1723 2437 1726
rect 2452 1723 2461 1726
rect 2586 1723 2597 1726
rect 2626 1723 2644 1726
rect 2738 1723 2748 1726
rect 2786 1723 2812 1726
rect 2874 1723 2900 1726
rect 2922 1723 2948 1726
rect 3042 1723 3068 1726
rect 3114 1723 3148 1726
rect 3258 1723 3276 1726
rect 1476 1713 1501 1716
rect 1532 1713 1541 1716
rect 1604 1713 1613 1716
rect 1692 1713 1709 1716
rect 1780 1713 1789 1716
rect 1794 1706 1797 1723
rect 2306 1716 2309 1723
rect 1964 1713 1973 1716
rect 2100 1713 2117 1716
rect 2140 1713 2149 1716
rect 2298 1713 2309 1716
rect 2506 1713 2532 1716
rect 2676 1713 2685 1716
rect 2916 1713 2933 1716
rect 442 1703 468 1706
rect 570 1703 620 1706
rect 1370 1703 1397 1706
rect 1442 1703 1461 1706
rect 1786 1703 1797 1706
rect 1930 1703 1973 1706
rect 2514 1703 2548 1706
rect 2650 1703 2668 1706
rect 14 1667 3490 1673
rect 2202 1653 2221 1656
rect 74 1643 85 1646
rect 74 1606 77 1643
rect 82 1616 85 1636
rect 338 1633 388 1636
rect 1098 1626 1101 1636
rect 1514 1633 1556 1636
rect 1634 1633 1684 1636
rect 1930 1633 1949 1636
rect 2154 1633 2172 1636
rect 180 1623 189 1626
rect 332 1623 349 1626
rect 396 1623 405 1626
rect 706 1616 709 1625
rect 804 1623 813 1626
rect 996 1623 1005 1626
rect 1092 1623 1101 1626
rect 1298 1623 1309 1626
rect 1356 1623 1365 1626
rect 1444 1623 1469 1626
rect 1514 1623 1540 1626
rect 1564 1623 1573 1626
rect 1658 1623 1668 1626
rect 1716 1623 1725 1626
rect 82 1613 92 1616
rect 130 1613 172 1616
rect 234 1613 276 1616
rect 482 1613 492 1616
rect 572 1613 589 1616
rect 604 1613 613 1616
rect 626 1613 660 1616
rect 706 1613 757 1616
rect 764 1613 773 1616
rect 778 1613 788 1616
rect 130 1606 133 1613
rect 74 1603 85 1606
rect 116 1603 133 1606
rect 220 1603 277 1606
rect 402 1603 426 1606
rect 530 1603 564 1606
rect 596 1603 645 1606
rect 708 1603 717 1606
rect 754 1605 757 1613
rect 810 1606 813 1623
rect 924 1613 980 1616
rect 1090 1613 1108 1616
rect 1164 1613 1173 1616
rect 1218 1613 1252 1616
rect 1276 1613 1301 1616
rect 1306 1606 1309 1623
rect 1402 1613 1428 1616
rect 810 1603 828 1606
rect 850 1603 876 1606
rect 900 1603 909 1606
rect 916 1603 957 1606
rect 1034 1603 1076 1606
rect 1156 1603 1189 1606
rect 1220 1603 1229 1606
rect 1306 1603 1324 1606
rect 1386 1603 1420 1606
rect 1444 1603 1453 1606
rect 1500 1603 1533 1606
rect 1594 1603 1604 1606
rect 1658 1603 1661 1623
rect 1826 1616 1829 1626
rect 1754 1613 1780 1616
rect 1812 1613 1829 1616
rect 1834 1613 1844 1616
rect 1850 1613 1884 1616
rect 1946 1615 1949 1633
rect 2156 1623 2165 1626
rect 1970 1613 2004 1616
rect 2068 1613 2077 1616
rect 2098 1613 2148 1616
rect 1804 1603 1821 1606
rect 1826 1603 1836 1606
rect 1882 1603 1892 1606
rect 1908 1603 1933 1606
rect 1994 1603 2012 1606
rect 2028 1603 2037 1606
rect 2042 1603 2060 1606
rect 810 1593 820 1596
rect 2074 1595 2077 1613
rect 2186 1596 2189 1646
rect 2202 1616 2205 1653
rect 2210 1633 2244 1636
rect 2346 1633 2365 1636
rect 2410 1633 2421 1636
rect 2346 1626 2349 1633
rect 2228 1623 2237 1626
rect 2332 1623 2349 1626
rect 2202 1613 2213 1616
rect 2258 1613 2268 1616
rect 2298 1613 2316 1616
rect 2418 1615 2421 1633
rect 2436 1623 2453 1626
rect 2474 1616 2477 1636
rect 2658 1626 2661 1646
rect 2786 1633 2821 1636
rect 2882 1633 2901 1636
rect 2540 1623 2557 1626
rect 2604 1623 2629 1626
rect 2644 1623 2653 1626
rect 2658 1623 2668 1626
rect 2778 1623 2812 1626
rect 2442 1613 2468 1616
rect 2474 1613 2508 1616
rect 2522 1613 2532 1616
rect 2602 1613 2636 1616
rect 2740 1613 2757 1616
rect 2818 1615 2821 1633
rect 2836 1623 2845 1626
rect 2874 1623 2892 1626
rect 2868 1613 2877 1616
rect 2898 1615 2901 1633
rect 3274 1616 3277 1636
rect 2922 1613 2964 1616
rect 3010 1606 3013 1614
rect 3018 1613 3060 1616
rect 3204 1613 3229 1616
rect 3274 1613 3285 1616
rect 2274 1603 2308 1606
rect 2332 1603 2341 1606
rect 2474 1603 2500 1606
rect 2562 1603 2580 1606
rect 2698 1603 2732 1606
rect 2842 1603 2860 1606
rect 2930 1603 2956 1606
rect 2970 1603 2988 1606
rect 3010 1603 3052 1606
rect 3066 1603 3092 1606
rect 3282 1605 3285 1613
rect 2186 1593 2213 1596
rect 2842 1593 2852 1596
rect 38 1567 3466 1573
rect 124 1543 133 1546
rect 82 1533 108 1536
rect 236 1533 245 1536
rect 90 1523 100 1526
rect 124 1523 133 1526
rect 130 1506 133 1523
rect 146 1506 149 1525
rect 164 1513 205 1516
rect 130 1503 149 1506
rect 282 1483 309 1486
rect 314 1483 317 1556
rect 442 1543 450 1546
rect 834 1543 852 1546
rect 866 1543 876 1546
rect 1330 1543 1356 1546
rect 362 1533 397 1536
rect 450 1533 460 1536
rect 482 1533 493 1536
rect 332 1523 341 1526
rect 348 1523 389 1526
rect 394 1525 397 1533
rect 430 1523 437 1526
rect 476 1523 485 1526
rect 434 1513 437 1523
rect 490 1516 493 1533
rect 538 1533 564 1536
rect 580 1533 636 1536
rect 812 1533 853 1536
rect 884 1533 901 1536
rect 994 1533 1004 1536
rect 1138 1533 1164 1536
rect 1202 1533 1205 1543
rect 1290 1536 1293 1543
rect 1370 1536 1373 1546
rect 1546 1543 1556 1546
rect 2106 1543 2124 1546
rect 2282 1536 2285 1546
rect 1258 1533 1276 1536
rect 1290 1533 1301 1536
rect 1308 1533 1341 1536
rect 1364 1533 1373 1536
rect 1378 1533 1388 1536
rect 1426 1533 1452 1536
rect 1564 1533 1589 1536
rect 1626 1533 1668 1536
rect 1794 1533 1804 1536
rect 538 1516 541 1533
rect 546 1523 555 1526
rect 594 1523 628 1526
rect 652 1523 669 1526
rect 482 1513 493 1516
rect 498 1513 508 1516
rect 532 1513 541 1516
rect 706 1513 740 1516
rect 482 1486 485 1513
rect 746 1506 749 1525
rect 770 1523 796 1526
rect 892 1523 917 1526
rect 932 1523 949 1526
rect 764 1513 773 1516
rect 940 1513 964 1516
rect 970 1506 973 1525
rect 1012 1523 1061 1526
rect 1130 1523 1172 1526
rect 1220 1523 1237 1526
rect 1317 1523 1333 1526
rect 1386 1523 1396 1526
rect 1426 1523 1460 1526
rect 1572 1523 1581 1526
rect 1124 1513 1157 1516
rect 1476 1513 1485 1516
rect 1500 1513 1509 1516
rect 1524 1513 1533 1516
rect 1586 1506 1589 1533
rect 1794 1523 1797 1533
rect 1818 1526 1821 1536
rect 1834 1533 1868 1536
rect 1890 1533 1900 1536
rect 1922 1533 1933 1536
rect 2034 1533 2068 1536
rect 2114 1533 2132 1536
rect 2170 1533 2180 1536
rect 2204 1533 2213 1536
rect 2218 1533 2244 1536
rect 2260 1533 2277 1536
rect 2282 1533 2316 1536
rect 2338 1533 2348 1536
rect 2378 1533 2412 1536
rect 1922 1526 1925 1533
rect 2426 1526 2429 1546
rect 2994 1543 3036 1546
rect 2474 1533 2508 1536
rect 2522 1533 2540 1536
rect 2562 1533 2573 1536
rect 2628 1533 2637 1536
rect 2676 1533 2709 1536
rect 2714 1533 2732 1536
rect 2738 1533 2756 1536
rect 2762 1533 2812 1536
rect 2836 1533 2845 1536
rect 1812 1523 1821 1526
rect 1876 1523 1885 1526
rect 1908 1523 1925 1526
rect 2050 1523 2076 1526
rect 2140 1523 2181 1526
rect 2226 1523 2236 1526
rect 2268 1523 2285 1526
rect 2298 1523 2356 1526
rect 2420 1523 2429 1526
rect 2498 1523 2516 1526
rect 2538 1523 2548 1526
rect 1716 1513 1757 1516
rect 1764 1513 1773 1516
rect 1788 1513 1797 1516
rect 1820 1513 1853 1516
rect 2204 1513 2229 1516
rect 2372 1513 2405 1516
rect 2468 1513 2477 1516
rect 2562 1506 2565 1533
rect 2850 1526 2853 1534
rect 2876 1533 2917 1536
rect 2946 1526 2949 1534
rect 3002 1533 3044 1536
rect 3274 1526 3277 1534
rect 2570 1523 2612 1526
rect 2626 1523 2653 1526
rect 2740 1523 2749 1526
rect 2770 1523 2820 1526
rect 2834 1523 2853 1526
rect 2922 1523 2932 1526
rect 2946 1523 2957 1526
rect 3156 1523 3181 1526
rect 3268 1523 3277 1526
rect 3370 1523 3380 1526
rect 2836 1513 2845 1516
rect 2954 1506 2957 1523
rect 2964 1513 2973 1516
rect 3060 1513 3069 1516
rect 3084 1513 3093 1516
rect 490 1503 524 1506
rect 714 1503 749 1506
rect 954 1503 973 1506
rect 1490 1503 1516 1506
rect 1586 1503 1612 1506
rect 1754 1503 1780 1506
rect 2562 1503 2573 1506
rect 2954 1503 2980 1506
rect 3058 1503 3076 1506
rect 482 1483 501 1486
rect 14 1467 3490 1473
rect 314 1433 340 1436
rect 172 1423 189 1426
rect 228 1423 253 1426
rect 138 1413 164 1416
rect 170 1413 196 1416
rect 210 1413 220 1416
rect 258 1413 276 1416
rect 354 1413 404 1416
rect 138 1406 141 1413
rect 116 1403 141 1406
rect 178 1403 188 1406
rect 202 1403 212 1406
rect 258 1396 261 1413
rect 410 1406 413 1425
rect 546 1416 549 1456
rect 1410 1443 1421 1446
rect 642 1433 660 1436
rect 746 1433 764 1436
rect 748 1423 757 1426
rect 454 1413 485 1416
rect 538 1413 555 1416
rect 588 1413 597 1416
rect 706 1413 724 1416
rect 538 1406 541 1413
rect 300 1403 309 1406
rect 386 1403 396 1406
rect 410 1403 421 1406
rect 450 1403 508 1406
rect 530 1403 541 1406
rect 586 1403 628 1406
rect 690 1403 715 1406
rect 234 1393 261 1396
rect 786 1386 789 1436
rect 868 1423 909 1426
rect 1260 1423 1269 1426
rect 794 1413 828 1416
rect 882 1413 916 1416
rect 1010 1413 1061 1416
rect 1058 1406 1061 1413
rect 1098 1406 1101 1415
rect 1106 1413 1140 1416
rect 1242 1413 1252 1416
rect 1338 1413 1364 1416
rect 810 1403 820 1406
rect 914 1403 924 1406
rect 938 1403 972 1406
rect 1058 1403 1076 1406
rect 1098 1403 1109 1406
rect 1114 1403 1132 1406
rect 1156 1403 1173 1406
rect 1186 1403 1196 1406
rect 1298 1403 1308 1406
rect 1314 1403 1323 1406
rect 1346 1403 1356 1406
rect 940 1393 965 1396
rect 1282 1393 1299 1396
rect 1410 1386 1413 1443
rect 1890 1433 1924 1436
rect 2090 1433 2109 1436
rect 1794 1423 1821 1426
rect 1860 1423 1908 1426
rect 1794 1416 1797 1423
rect 2066 1416 2069 1424
rect 2074 1423 2100 1426
rect 2130 1423 2133 1446
rect 2298 1433 2308 1436
rect 2522 1433 2533 1436
rect 2914 1433 2973 1436
rect 3058 1433 3085 1436
rect 2228 1423 2237 1426
rect 2316 1423 2341 1426
rect 1418 1413 1436 1416
rect 1466 1413 1476 1416
rect 1562 1413 1572 1416
rect 1644 1413 1653 1416
rect 1746 1413 1764 1416
rect 1778 1413 1797 1416
rect 1802 1413 1828 1416
rect 1842 1413 1852 1416
rect 1986 1413 2028 1416
rect 2066 1413 2093 1416
rect 2188 1413 2205 1416
rect 2330 1413 2364 1416
rect 2378 1413 2396 1416
rect 2434 1413 2460 1416
rect 2484 1413 2525 1416
rect 1778 1406 1781 1413
rect 1482 1403 1532 1406
rect 1578 1403 1636 1406
rect 1660 1403 1717 1406
rect 1724 1403 1756 1406
rect 1986 1396 1989 1413
rect 2010 1403 2020 1406
rect 2130 1403 2172 1406
rect 2202 1405 2205 1413
rect 2242 1403 2276 1406
rect 2394 1403 2404 1406
rect 2426 1403 2452 1406
rect 2530 1396 2533 1433
rect 2698 1423 2717 1426
rect 2868 1423 2877 1426
rect 2914 1423 2964 1426
rect 2698 1416 2701 1423
rect 2612 1413 2629 1416
rect 2634 1413 2652 1416
rect 2684 1413 2701 1416
rect 2706 1413 2732 1416
rect 2970 1415 2973 1433
rect 3106 1426 3109 1436
rect 3066 1423 3076 1426
rect 3100 1423 3109 1426
rect 3396 1423 3405 1426
rect 2706 1406 2709 1413
rect 2994 1406 2997 1416
rect 3132 1413 3157 1416
rect 3170 1413 3180 1416
rect 3268 1413 3277 1416
rect 3292 1413 3317 1416
rect 3370 1413 3380 1416
rect 2570 1403 2596 1406
rect 2618 1403 2660 1406
rect 2676 1403 2709 1406
rect 2714 1403 2724 1406
rect 2746 1403 2780 1406
rect 2810 1403 2844 1406
rect 2994 1403 3004 1406
rect 3106 1403 3124 1406
rect 3242 1403 3269 1406
rect 3284 1403 3301 1406
rect 2714 1396 2717 1403
rect 1980 1393 1989 1396
rect 2188 1393 2197 1396
rect 2498 1393 2533 1396
rect 2612 1393 2621 1396
rect 2690 1393 2717 1396
rect 3106 1393 3116 1396
rect 3234 1393 3252 1396
rect 786 1383 805 1386
rect 1410 1383 1421 1386
rect 3298 1383 3301 1403
rect 3314 1396 3317 1413
rect 3338 1403 3356 1406
rect 3362 1403 3372 1406
rect 3396 1403 3413 1406
rect 3314 1393 3348 1396
rect 38 1367 3466 1373
rect 106 1343 133 1346
rect 106 1326 109 1343
rect 164 1333 213 1336
rect 218 1333 228 1336
rect 92 1323 109 1326
rect 114 1323 140 1326
rect 236 1323 261 1326
rect 306 1316 309 1346
rect 866 1343 876 1346
rect 1034 1336 1037 1346
rect 314 1323 332 1326
rect 378 1323 381 1335
rect 466 1333 484 1336
rect 508 1333 573 1336
rect 676 1333 693 1336
rect 754 1333 764 1336
rect 850 1333 884 1336
rect 906 1333 932 1336
rect 962 1333 972 1336
rect 1004 1333 1037 1336
rect 1050 1333 1076 1336
rect 1146 1333 1156 1336
rect 1188 1333 1221 1336
rect 906 1326 909 1333
rect 1218 1326 1221 1333
rect 1250 1326 1253 1345
rect 1260 1333 1277 1336
rect 1290 1333 1323 1336
rect 1386 1326 1389 1345
rect 1652 1343 1685 1346
rect 1890 1336 1893 1356
rect 2546 1353 2581 1356
rect 1906 1343 1924 1346
rect 2082 1343 2109 1346
rect 2370 1343 2381 1346
rect 2434 1343 2460 1346
rect 2634 1343 2644 1346
rect 1396 1333 1445 1336
rect 1514 1333 1548 1336
rect 1580 1333 1589 1336
rect 1610 1333 1636 1336
rect 1698 1333 1708 1336
rect 1732 1333 1749 1336
rect 1802 1333 1852 1336
rect 1890 1333 1932 1336
rect 2050 1333 2060 1336
rect 2114 1333 2124 1336
rect 2156 1333 2189 1336
rect 2242 1333 2260 1336
rect 2284 1333 2293 1336
rect 2298 1333 2324 1336
rect 2348 1333 2365 1336
rect 2370 1326 2373 1343
rect 2378 1333 2388 1336
rect 2442 1333 2468 1336
rect 2562 1333 2588 1336
rect 2618 1333 2652 1336
rect 2684 1333 2749 1336
rect 2754 1333 2764 1336
rect 2788 1333 2813 1336
rect 2818 1333 2836 1336
rect 2874 1333 2916 1336
rect 2948 1333 2965 1336
rect 2970 1333 2980 1336
rect 3002 1333 3036 1336
rect 3290 1333 3340 1336
rect 2754 1326 2757 1333
rect 420 1323 437 1326
rect 458 1323 492 1326
rect 516 1323 525 1326
rect 562 1323 572 1326
rect 604 1323 613 1326
rect 642 1323 660 1326
rect 754 1323 772 1326
rect 300 1313 309 1316
rect 676 1313 709 1316
rect 794 1313 820 1316
rect 826 1306 829 1325
rect 892 1323 909 1326
rect 914 1323 940 1326
rect 1084 1323 1093 1326
rect 1100 1323 1109 1326
rect 1122 1323 1164 1326
rect 1218 1323 1253 1326
rect 1274 1323 1332 1326
rect 1338 1323 1389 1326
rect 1426 1323 1460 1326
rect 1498 1323 1556 1326
rect 1602 1323 1628 1326
rect 1652 1323 1693 1326
rect 1988 1323 2021 1326
rect 2036 1323 2045 1326
rect 2068 1323 2085 1326
rect 2258 1323 2268 1326
rect 2370 1323 2381 1326
rect 2476 1323 2493 1326
rect 2578 1323 2596 1326
rect 2612 1323 2637 1326
rect 2668 1323 2677 1326
rect 2706 1323 2757 1326
rect 2802 1323 2844 1326
rect 2874 1323 2924 1326
rect 2996 1323 3044 1326
rect 3066 1323 3085 1326
rect 3156 1323 3181 1326
rect 3212 1323 3229 1326
rect 3242 1323 3252 1326
rect 3284 1323 3301 1326
rect 3314 1323 3348 1326
rect 3362 1323 3389 1326
rect 3404 1323 3413 1326
rect 844 1313 861 1316
rect 1732 1313 1741 1316
rect 1772 1313 1781 1316
rect 2220 1313 2237 1316
rect 2348 1313 2373 1316
rect 2378 1313 2381 1323
rect 3268 1313 3277 1316
rect 3362 1315 3365 1323
rect 250 1303 292 1306
rect 810 1303 829 1306
rect 1018 1303 1053 1306
rect 2178 1303 2212 1306
rect 14 1267 3490 1273
rect 1434 1253 1461 1256
rect 258 1243 285 1246
rect 186 1233 244 1236
rect 258 1233 316 1236
rect 650 1233 660 1236
rect 882 1233 893 1236
rect 1738 1233 1788 1236
rect 1802 1233 1852 1236
rect 1986 1233 2013 1236
rect 124 1223 157 1226
rect 186 1223 228 1226
rect 252 1223 269 1226
rect 324 1223 357 1226
rect 604 1223 613 1226
rect 186 1216 189 1223
rect 754 1216 757 1225
rect 818 1216 821 1226
rect 178 1213 189 1216
rect 362 1213 372 1216
rect 418 1213 460 1216
rect 684 1213 693 1216
rect 722 1213 748 1216
rect 754 1213 772 1216
rect 810 1213 828 1216
rect 852 1213 861 1216
rect 890 1215 893 1233
rect 908 1223 949 1226
rect 1364 1223 1389 1226
rect 1572 1223 1589 1226
rect 1732 1223 1765 1226
rect 1802 1223 1845 1226
rect 2010 1216 2013 1233
rect 2028 1223 2053 1226
rect 2178 1216 2181 1246
rect 3186 1233 3197 1236
rect 3242 1233 3268 1236
rect 3386 1233 3404 1236
rect 2220 1223 2237 1226
rect 3090 1216 3093 1226
rect 3156 1223 3181 1226
rect 946 1213 964 1216
rect 1188 1213 1197 1216
rect 1212 1213 1268 1216
rect 1362 1213 1396 1216
rect 1420 1213 1429 1216
rect 1458 1213 1469 1216
rect 1506 1213 1556 1216
rect 1586 1213 1604 1216
rect 1642 1213 1669 1216
rect 1692 1213 1716 1216
rect 1930 1213 1941 1216
rect 1954 1213 1964 1216
rect 2010 1213 2020 1216
rect 2026 1213 2068 1216
rect 2090 1213 2132 1216
rect 2164 1213 2189 1216
rect 2212 1213 2245 1216
rect 82 1203 100 1206
rect 124 1203 133 1206
rect 346 1203 380 1206
rect 396 1203 405 1206
rect 442 1203 452 1206
rect 524 1203 565 1206
rect 698 1203 740 1206
rect 810 1183 813 1213
rect 818 1203 836 1206
rect 938 1203 956 1206
rect 988 1203 1021 1206
rect 1058 1203 1084 1206
rect 1122 1203 1132 1206
rect 1146 1203 1180 1206
rect 852 1193 869 1196
rect 1090 1193 1124 1196
rect 1194 1195 1197 1213
rect 1298 1203 1340 1206
rect 1386 1203 1404 1206
rect 1458 1196 1461 1213
rect 1506 1206 1509 1213
rect 1642 1206 1645 1213
rect 1938 1206 1941 1213
rect 2250 1206 2253 1215
rect 2378 1213 2396 1216
rect 2428 1213 2445 1216
rect 2618 1213 2660 1216
rect 2716 1213 2749 1216
rect 2820 1213 2829 1216
rect 2874 1213 2908 1216
rect 3050 1213 3060 1216
rect 3084 1213 3093 1216
rect 3194 1215 3197 1233
rect 3242 1223 3261 1226
rect 3282 1213 3324 1216
rect 1498 1203 1509 1206
rect 1530 1203 1548 1206
rect 1602 1203 1612 1206
rect 1628 1203 1645 1206
rect 1650 1203 1684 1206
rect 1698 1203 1708 1206
rect 1866 1203 1892 1206
rect 1916 1203 1933 1206
rect 1938 1203 1956 1206
rect 1986 1203 2012 1206
rect 2106 1203 2140 1206
rect 2170 1203 2204 1206
rect 2226 1203 2253 1206
rect 2276 1203 2285 1206
rect 2298 1203 2332 1206
rect 2410 1203 2420 1206
rect 2434 1203 2484 1206
rect 2522 1203 2564 1206
rect 2666 1203 2684 1206
rect 2764 1203 2805 1206
rect 2812 1203 2821 1206
rect 2836 1203 2869 1206
rect 2874 1203 2900 1206
rect 2932 1203 2941 1206
rect 2978 1203 3012 1206
rect 3036 1203 3045 1206
rect 3106 1203 3132 1206
rect 3330 1205 3333 1226
rect 3354 1223 3388 1226
rect 1298 1193 1325 1196
rect 1420 1193 1461 1196
rect 2746 1193 2756 1196
rect 2818 1193 2828 1196
rect 3084 1193 3093 1196
rect 38 1167 3466 1173
rect 564 1143 581 1146
rect 626 1136 629 1156
rect 898 1143 908 1146
rect 946 1143 956 1146
rect 978 1143 996 1146
rect 1026 1143 1061 1146
rect 1274 1143 1300 1146
rect 1834 1143 1868 1146
rect 82 1133 100 1136
rect 162 1133 196 1136
rect 236 1133 293 1136
rect 378 1133 404 1136
rect 514 1133 548 1136
rect 626 1133 652 1136
rect 882 1133 916 1136
rect 946 1133 964 1136
rect 1010 1133 1068 1136
rect 1100 1133 1125 1136
rect 1154 1133 1188 1136
rect 1266 1133 1308 1136
rect 1322 1133 1349 1136
rect 1402 1133 1420 1136
rect 82 1093 85 1133
rect 946 1126 949 1133
rect 130 1123 140 1126
rect 186 1123 197 1126
rect 282 1123 308 1126
rect 378 1123 396 1126
rect 450 1123 460 1126
rect 506 1123 540 1126
rect 564 1123 589 1126
rect 594 1123 604 1126
rect 618 1123 660 1126
rect 722 1123 764 1126
rect 786 1123 797 1126
rect 804 1123 821 1126
rect 924 1123 949 1126
rect 1012 1123 1045 1126
rect 1050 1123 1076 1126
rect 1154 1123 1157 1133
rect 1322 1126 1325 1133
rect 1554 1126 1557 1136
rect 1570 1133 1580 1136
rect 1610 1126 1613 1134
rect 1690 1133 1724 1136
rect 1738 1133 1780 1136
rect 1796 1133 1869 1136
rect 1908 1133 1941 1136
rect 1186 1123 1196 1126
rect 1252 1123 1301 1126
rect 1317 1123 1325 1126
rect 186 1116 189 1123
rect 282 1116 285 1123
rect 378 1116 381 1123
rect 786 1116 789 1123
rect 148 1113 189 1116
rect 250 1113 285 1116
rect 348 1113 381 1116
rect 620 1113 645 1116
rect 684 1113 693 1116
rect 780 1113 789 1116
rect 1156 1113 1189 1116
rect 1204 1113 1221 1116
rect 1260 1113 1269 1116
rect 1322 1106 1325 1123
rect 1330 1113 1356 1116
rect 1362 1106 1365 1125
rect 1476 1123 1485 1126
rect 1522 1106 1525 1125
rect 1554 1123 1588 1126
rect 1594 1123 1613 1126
rect 1620 1123 1629 1126
rect 1698 1123 1732 1126
rect 1738 1123 1772 1126
rect 1916 1123 1933 1126
rect 1938 1123 1941 1133
rect 1540 1113 1557 1116
rect 1594 1113 1597 1123
rect 1930 1116 1933 1123
rect 1930 1113 1965 1116
rect 674 1103 700 1106
rect 1322 1103 1365 1106
rect 1498 1103 1525 1106
rect 2002 1103 2005 1126
rect 2010 1103 2013 1146
rect 2738 1143 2772 1146
rect 2842 1143 2868 1146
rect 2914 1143 2924 1146
rect 2162 1133 2188 1136
rect 2202 1133 2236 1136
rect 2242 1133 2276 1136
rect 2298 1133 2332 1136
rect 2356 1133 2397 1136
rect 2402 1133 2412 1136
rect 2506 1133 2524 1136
rect 2586 1133 2604 1136
rect 2042 1123 2109 1126
rect 2178 1123 2196 1126
rect 2244 1123 2261 1126
rect 2266 1123 2284 1126
rect 2362 1123 2404 1126
rect 2442 1123 2500 1126
rect 2506 1123 2532 1126
rect 2586 1123 2589 1133
rect 2738 1126 2741 1143
rect 2938 1136 2941 1146
rect 2746 1133 2780 1136
rect 2826 1126 2829 1134
rect 2858 1133 2876 1136
rect 2932 1133 2941 1136
rect 3308 1133 3325 1136
rect 2706 1123 2741 1126
rect 2788 1123 2829 1126
rect 2892 1123 2925 1126
rect 2940 1123 2949 1126
rect 2978 1123 2996 1126
rect 3156 1123 3181 1126
rect 3226 1123 3284 1126
rect 3314 1123 3381 1126
rect 2978 1116 2981 1123
rect 2092 1113 2117 1116
rect 2124 1113 2133 1116
rect 2148 1113 2181 1116
rect 2292 1113 2317 1116
rect 2508 1113 2525 1116
rect 2540 1113 2549 1116
rect 2954 1113 2981 1116
rect 3378 1116 3381 1123
rect 3378 1113 3388 1116
rect 2114 1106 2117 1113
rect 3394 1106 3397 1125
rect 3412 1113 3429 1116
rect 2114 1103 2140 1106
rect 3314 1103 3341 1106
rect 3362 1103 3397 1106
rect 162 1093 181 1096
rect 3226 1083 3269 1086
rect 14 1067 3490 1073
rect 1978 1053 1997 1056
rect 324 1023 349 1026
rect 578 1016 581 1046
rect 3378 1043 3389 1046
rect 666 1033 692 1036
rect 1058 1033 1101 1036
rect 1882 1033 1909 1036
rect 2074 1033 2092 1036
rect 2170 1033 2204 1036
rect 2578 1033 2613 1036
rect 2738 1033 2780 1036
rect 2794 1033 2837 1036
rect 2874 1033 2900 1036
rect 2946 1033 2972 1036
rect 666 1016 669 1033
rect 996 1023 1021 1026
rect 1082 1023 1092 1026
rect 148 1013 181 1016
rect 194 1013 204 1016
rect 236 1013 261 1016
rect 282 1013 308 1016
rect 372 1013 381 1016
rect 442 1013 460 1016
rect 532 1013 541 1016
rect 548 1013 581 1016
rect 612 1013 637 1016
rect 644 1013 669 1016
rect 730 1013 756 1016
rect 810 1013 820 1016
rect 906 1013 924 1016
rect 994 1013 1028 1016
rect 1052 1013 1061 1016
rect 1098 1015 1101 1033
rect 1116 1023 1157 1026
rect 1796 1023 1829 1026
rect 2050 1023 2076 1026
rect 2100 1023 2141 1026
rect 2156 1023 2173 1026
rect 2212 1023 2229 1026
rect 2276 1023 2301 1026
rect 2332 1023 2349 1026
rect 2418 1023 2437 1026
rect 2532 1023 2549 1026
rect 2570 1023 2604 1026
rect 1154 1016 1157 1023
rect 2418 1016 2421 1023
rect 1154 1013 1165 1016
rect 1186 1013 1205 1016
rect 1308 1013 1317 1016
rect 1364 1013 1389 1016
rect 1474 1013 1509 1016
rect 1524 1013 1533 1016
rect 1554 1013 1596 1016
rect 1746 1013 1780 1016
rect 1866 1013 1876 1016
rect 1890 1013 1925 1016
rect 1962 1013 1972 1016
rect 2002 1013 2028 1016
rect 2058 1013 2069 1016
rect 2148 1013 2181 1016
rect 634 1006 637 1013
rect 114 1003 140 1006
rect 178 1003 212 1006
rect 228 1003 253 1006
rect 324 1003 349 1006
rect 490 1003 516 1006
rect 562 1003 604 1006
rect 626 1005 637 1006
rect 626 1003 636 1005
rect 738 1003 748 1006
rect 778 1003 828 1006
rect 892 1003 909 1006
rect 930 1003 972 1006
rect 1026 1003 1036 1006
rect 1186 1005 1189 1013
rect 1194 1003 1220 1006
rect 1290 1003 1300 1006
rect 1314 996 1317 1013
rect 1322 1003 1356 1006
rect 1404 1003 1437 1006
rect 330 993 356 996
rect 466 993 508 996
rect 1052 993 1077 996
rect 1234 993 1276 996
rect 1314 993 1348 996
rect 1362 993 1396 996
rect 1506 995 1509 1013
rect 1530 1003 1588 1006
rect 1650 1003 1660 1006
rect 1684 1003 1725 1006
rect 1732 1003 1772 1006
rect 1796 1003 1805 1006
rect 1844 1003 1853 1006
rect 1858 1003 1868 1006
rect 1882 1003 1924 1006
rect 2044 1003 2061 1006
rect 2066 996 2069 1013
rect 2106 1003 2140 1006
rect 2194 1003 2197 1014
rect 2218 1013 2245 1016
rect 2362 1013 2372 1016
rect 2404 1013 2421 1016
rect 2426 1013 2444 1016
rect 2498 1013 2524 1016
rect 2538 1013 2573 1016
rect 2610 1015 2613 1033
rect 2802 1023 2828 1026
rect 2634 1013 2644 1016
rect 2650 1013 2708 1016
rect 2834 1015 2837 1033
rect 3378 1026 3381 1043
rect 3386 1033 3412 1036
rect 2858 1023 2884 1026
rect 2914 1023 2956 1026
rect 3188 1023 3229 1026
rect 3378 1023 3396 1026
rect 3420 1023 3429 1026
rect 2986 1013 2996 1016
rect 3060 1013 3085 1016
rect 3116 1013 3133 1016
rect 3226 1013 3236 1016
rect 3268 1013 3277 1016
rect 2218 1003 2252 1006
rect 2332 1003 2341 1006
rect 2354 1003 2380 1006
rect 2442 1003 2452 1006
rect 2468 1003 2501 1006
rect 2538 1003 2556 1006
rect 2724 1003 2749 1006
rect 3188 1003 3237 1006
rect 3260 1003 3292 1006
rect 3346 1003 3364 1006
rect 1690 993 1724 996
rect 2050 993 2069 996
rect 3338 993 3356 996
rect 38 967 3466 973
rect 74 943 85 946
rect 130 943 164 946
rect 74 926 77 943
rect 82 933 92 936
rect 138 933 172 936
rect 202 933 212 936
rect 226 933 252 936
rect 202 926 205 933
rect 74 923 100 926
rect 180 923 205 926
rect 116 913 157 916
rect 226 913 229 933
rect 282 926 285 945
rect 562 936 565 956
rect 1762 953 1797 956
rect 1234 943 1260 946
rect 1290 943 1300 946
rect 1314 943 1356 946
rect 292 933 301 936
rect 426 933 460 936
rect 524 933 565 936
rect 660 933 669 936
rect 754 933 764 936
rect 788 933 797 936
rect 866 933 892 936
rect 978 933 996 936
rect 1026 933 1052 936
rect 1156 933 1181 936
rect 1212 933 1229 936
rect 1274 933 1308 936
rect 1364 933 1389 936
rect 1500 933 1533 936
rect 1572 933 1605 936
rect 1178 926 1181 933
rect 260 923 285 926
rect 300 923 309 926
rect 378 923 412 926
rect 490 923 500 926
rect 532 923 549 926
rect 626 923 644 926
rect 420 913 445 916
rect 562 913 572 916
rect 660 913 693 916
rect 706 906 709 925
rect 730 923 772 926
rect 970 923 1004 926
rect 1018 923 1044 926
rect 1082 923 1140 926
rect 1178 923 1196 926
rect 1210 923 1221 926
rect 1316 923 1349 926
rect 1386 923 1389 933
rect 1530 926 1533 933
rect 1450 923 1484 926
rect 1530 923 1556 926
rect 1602 923 1613 926
rect 1626 925 1629 946
rect 1666 943 1700 946
rect 1722 943 1740 946
rect 1762 936 1765 953
rect 1842 943 1860 946
rect 2362 943 2381 946
rect 1666 933 1708 936
rect 1748 933 1765 936
rect 1778 933 1804 936
rect 1828 933 1853 936
rect 1868 933 1885 936
rect 1946 933 1979 936
rect 2004 933 2029 936
rect 2074 933 2092 936
rect 2162 933 2172 936
rect 2188 933 2229 936
rect 2274 933 2284 936
rect 2306 933 2332 936
rect 2362 933 2396 936
rect 2418 933 2468 936
rect 2484 933 2501 936
rect 2514 933 2532 936
rect 2578 933 2604 936
rect 2650 933 2660 936
rect 2690 933 2700 936
rect 1634 923 1685 926
rect 1756 923 1765 926
rect 1970 923 1987 926
rect 2044 923 2053 926
rect 2116 923 2149 926
rect 2266 923 2292 926
rect 2340 923 2357 926
rect 2420 923 2445 926
rect 2450 923 2460 926
rect 2506 923 2524 926
rect 2556 923 2573 926
rect 2586 923 2596 926
rect 2658 923 2668 926
rect 1218 916 1221 923
rect 1602 916 1605 923
rect 2450 916 2453 923
rect 2882 916 2885 946
rect 2946 933 2972 936
rect 3242 933 3252 936
rect 788 913 821 916
rect 826 906 829 915
rect 852 913 861 916
rect 1018 913 1037 916
rect 1218 913 1237 916
rect 1402 913 1412 916
rect 1436 913 1469 916
rect 1572 913 1605 916
rect 1906 913 1916 916
rect 1940 913 1949 916
rect 2202 913 2236 916
rect 2300 913 2309 916
rect 2442 913 2453 916
rect 2738 913 2748 916
rect 2804 913 2813 916
rect 2842 913 2852 916
rect 2876 913 2885 916
rect 2914 906 2917 925
rect 2938 923 2980 926
rect 2986 923 2996 926
rect 3076 923 3101 926
rect 3132 923 3141 926
rect 3146 923 3164 926
rect 3284 923 3309 926
rect 3330 925 3333 946
rect 3354 933 3372 936
rect 3380 924 3396 927
rect 3306 916 3309 923
rect 2932 913 2957 916
rect 3306 913 3324 916
rect 338 903 364 906
rect 562 903 588 906
rect 674 903 709 906
rect 794 903 829 906
rect 834 903 844 906
rect 1410 903 1428 906
rect 1898 903 1932 906
rect 2226 903 2252 906
rect 2778 903 2820 906
rect 2834 903 2868 906
rect 2882 903 2917 906
rect 14 867 3490 873
rect 3410 853 3429 856
rect 218 833 244 836
rect 266 833 308 836
rect 498 833 509 836
rect 642 833 684 836
rect 906 833 924 836
rect 1882 833 1908 836
rect 2194 833 2252 836
rect 108 823 141 826
rect 82 813 100 816
rect 218 813 221 833
rect 274 823 292 826
rect 316 823 341 826
rect 338 813 356 816
rect 388 813 429 816
rect 468 813 493 816
rect 426 806 429 813
rect 82 803 92 806
rect 172 803 213 806
rect 380 803 405 806
rect 426 803 444 806
rect 490 796 493 813
rect 498 806 501 833
rect 668 823 677 826
rect 890 823 908 826
rect 1004 823 1013 826
rect 1660 823 1669 826
rect 1850 823 1892 826
rect 1916 823 1957 826
rect 506 813 516 816
rect 578 813 604 816
rect 764 813 773 816
rect 802 813 868 816
rect 890 806 893 823
rect 2074 816 2077 826
rect 2210 823 2236 826
rect 2260 823 2269 826
rect 2428 823 2453 826
rect 2620 823 2629 826
rect 2898 823 2909 826
rect 2964 823 2989 826
rect 3140 823 3149 826
rect 1018 813 1044 816
rect 1074 813 1108 816
rect 1122 813 1148 816
rect 1178 813 1221 816
rect 1228 813 1277 816
rect 1330 813 1364 816
rect 1402 813 1444 816
rect 1490 813 1556 816
rect 1772 813 1781 816
rect 1786 813 1820 816
rect 1844 813 1885 816
rect 1930 813 1972 816
rect 2002 813 2044 816
rect 2074 813 2149 816
rect 2354 813 2388 816
rect 2394 813 2420 816
rect 2458 813 2468 816
rect 2474 813 2516 816
rect 2532 813 2549 816
rect 2618 813 2652 816
rect 2756 813 2781 816
rect 2868 813 2893 816
rect 1786 806 1789 813
rect 498 803 524 806
rect 540 803 612 806
rect 762 803 772 806
rect 796 803 813 806
rect 884 803 893 806
rect 946 803 980 806
rect 1004 803 1021 806
rect 1066 803 1100 806
rect 1122 803 1140 806
rect 1266 803 1276 806
rect 1314 803 1356 806
rect 1410 803 1436 806
rect 1450 803 1468 806
rect 1492 803 1501 806
rect 1514 803 1548 806
rect 1580 803 1589 806
rect 1618 803 1636 806
rect 1660 803 1709 806
rect 1716 803 1733 806
rect 1770 803 1797 806
rect 1922 803 1964 806
rect 1988 803 2013 806
rect 2018 803 2036 806
rect 2106 803 2124 806
rect 2138 803 2172 806
rect 2266 803 2316 806
rect 2018 796 2021 803
rect 2354 796 2357 813
rect 490 793 509 796
rect 738 793 748 796
rect 1738 793 1756 796
rect 2002 793 2021 796
rect 2332 793 2357 796
rect 2394 793 2397 813
rect 2898 807 2901 823
rect 3028 813 3053 816
rect 3084 813 3093 816
rect 3106 813 3124 816
rect 3284 813 3293 816
rect 3300 813 3333 816
rect 2658 803 2676 806
rect 3090 803 3116 806
rect 3186 803 3229 806
rect 3266 803 3276 806
rect 3330 795 3333 813
rect 3346 803 3372 806
rect 2266 783 2301 786
rect 38 767 3466 773
rect 2258 753 2269 756
rect 1002 743 1060 746
rect 1122 736 1125 746
rect 1482 743 1500 746
rect 2258 736 2261 753
rect 3226 746 3229 756
rect 2322 743 2341 746
rect 66 733 100 736
rect 154 733 204 736
rect 252 733 285 736
rect 314 733 324 736
rect 338 733 404 736
rect 420 733 437 736
rect 458 733 477 736
rect 434 726 437 733
rect 130 723 140 726
rect 162 723 212 726
rect 266 723 308 726
rect 332 723 341 726
rect 434 723 469 726
rect 474 716 477 733
rect 586 733 621 736
rect 642 733 652 736
rect 708 733 717 736
rect 738 733 748 736
rect 866 733 876 736
rect 900 733 909 736
rect 986 733 996 736
rect 1122 733 1164 736
rect 1250 733 1261 736
rect 538 723 556 726
rect 586 725 589 733
rect 986 726 989 733
rect 594 723 636 726
rect 660 723 693 726
rect 716 723 725 726
rect 730 723 756 726
rect 786 723 812 726
rect 914 723 964 726
rect 978 723 989 726
rect 1004 723 1061 726
rect 1122 723 1172 726
rect 1228 723 1253 726
rect 340 713 381 716
rect 474 713 500 716
rect 978 715 981 723
rect 1258 716 1261 733
rect 1322 726 1325 734
rect 1348 733 1365 736
rect 1418 733 1444 736
rect 1498 733 1508 736
rect 1514 733 1532 736
rect 1554 733 1564 736
rect 1594 733 1620 736
rect 1644 733 1661 736
rect 1666 733 1684 736
rect 1778 733 1788 736
rect 1810 733 1836 736
rect 2186 733 2220 736
rect 2236 733 2261 736
rect 2266 733 2292 736
rect 1300 723 1325 726
rect 1514 725 1517 733
rect 1554 726 1557 733
rect 1530 723 1557 726
rect 1588 723 1621 726
rect 1658 723 1676 726
rect 1084 713 1093 716
rect 1236 713 1261 716
rect 1348 713 1381 716
rect 1378 706 1381 713
rect 146 703 205 706
rect 1082 703 1100 706
rect 1378 703 1397 706
rect 1658 693 1661 723
rect 1754 706 1757 725
rect 1778 723 1796 726
rect 1844 723 1853 726
rect 1906 723 1932 726
rect 1858 713 1876 716
rect 1900 713 1909 716
rect 1938 713 1964 716
rect 1988 713 2013 716
rect 2044 713 2077 716
rect 1714 703 1757 706
rect 1906 693 1909 713
rect 2010 706 2013 713
rect 2090 706 2093 725
rect 2114 723 2140 726
rect 2172 723 2212 726
rect 2244 723 2269 726
rect 2274 723 2284 726
rect 2274 716 2277 723
rect 2108 713 2133 716
rect 2250 713 2277 716
rect 2010 703 2029 706
rect 2050 703 2093 706
rect 2338 686 2341 743
rect 2946 743 2965 746
rect 3220 743 3229 746
rect 2946 736 2949 743
rect 2386 733 2428 736
rect 2444 733 2477 736
rect 2516 733 2533 736
rect 2562 733 2580 736
rect 2602 733 2612 736
rect 2778 733 2788 736
rect 2836 733 2852 736
rect 2932 733 2949 736
rect 2954 733 2980 736
rect 3114 733 3132 736
rect 3218 733 3236 736
rect 3306 733 3332 736
rect 3354 733 3364 736
rect 3066 726 3069 733
rect 2380 723 2389 726
rect 2402 723 2420 726
rect 2490 723 2500 726
rect 2538 723 2548 726
rect 2652 723 2661 726
rect 2716 723 2741 726
rect 2812 723 2845 726
rect 2866 723 2908 726
rect 3066 723 3108 726
rect 3122 723 3140 726
rect 3220 723 3229 726
rect 3234 723 3244 726
rect 3362 723 3372 726
rect 3410 723 3420 726
rect 3122 716 3125 723
rect 3234 716 3237 723
rect 3116 713 3125 716
rect 3156 713 3165 716
rect 3226 713 3237 716
rect 3260 713 3269 716
rect 3300 713 3317 716
rect 2322 683 2341 686
rect 14 667 3490 673
rect 250 633 300 636
rect 930 633 964 636
rect 1034 633 1052 636
rect 1282 633 1309 636
rect 116 623 141 626
rect 156 623 181 626
rect 308 623 333 626
rect 636 623 645 626
rect 692 623 725 626
rect 788 623 805 626
rect 852 623 877 626
rect 948 623 957 626
rect 972 623 989 626
rect 1036 623 1045 626
rect 1252 623 1269 626
rect 1274 623 1300 626
rect 330 616 333 623
rect 722 616 725 623
rect 874 616 877 623
rect 1266 616 1269 623
rect 108 613 133 616
rect 148 613 165 616
rect 228 603 277 606
rect 290 593 293 615
rect 330 613 348 616
rect 474 613 500 616
rect 506 613 548 616
rect 564 613 613 616
rect 634 613 669 616
rect 722 613 733 616
rect 740 613 765 616
rect 786 613 836 616
rect 874 613 885 616
rect 1074 613 1108 616
rect 1122 613 1132 616
rect 1162 613 1188 616
rect 1218 613 1236 616
rect 1266 613 1293 616
rect 1306 615 1309 633
rect 1482 633 1508 636
rect 1618 633 1629 636
rect 1324 623 1341 626
rect 1482 616 1485 633
rect 1330 613 1356 616
rect 1452 613 1485 616
rect 1596 613 1613 616
rect 1626 615 1629 633
rect 1754 633 1780 636
rect 1708 623 1717 626
rect 1754 616 1757 633
rect 2108 623 2133 626
rect 2148 623 2173 626
rect 2188 623 2205 626
rect 2330 616 2333 636
rect 2338 633 2356 636
rect 2386 633 2420 636
rect 2364 623 2397 626
rect 2428 623 2453 626
rect 2468 623 2501 626
rect 2594 623 2613 626
rect 3276 623 3301 626
rect 2610 616 2613 623
rect 1650 613 1692 616
rect 1706 613 1725 616
rect 1732 613 1757 616
rect 1794 613 1804 616
rect 1922 613 1940 616
rect 1954 613 1980 616
rect 2002 613 2028 616
rect 2140 613 2165 616
rect 2180 613 2205 616
rect 2314 613 2333 616
rect 2434 613 2460 616
rect 2490 613 2508 616
rect 2540 613 2549 616
rect 2554 613 2605 616
rect 2610 613 2620 616
rect 2748 613 2757 616
rect 2874 613 2948 616
rect 2962 613 2973 616
rect 3002 613 3028 616
rect 3042 613 3060 616
rect 3106 613 3124 616
rect 3146 613 3156 616
rect 3202 613 3260 616
rect 372 603 444 606
rect 530 603 540 606
rect 594 603 612 606
rect 666 605 669 613
rect 730 605 733 613
rect 858 603 884 606
rect 908 603 917 606
rect 1066 603 1100 606
rect 1170 603 1180 606
rect 1338 603 1348 606
rect 1386 603 1412 606
rect 1722 605 1725 613
rect 1810 603 1868 606
rect 1946 603 1972 606
rect 1986 603 2020 606
rect 2044 603 2069 606
rect 2114 603 2132 606
rect 2146 603 2172 606
rect 2194 603 2228 606
rect 2314 605 2317 613
rect 2554 606 2557 613
rect 2602 606 2605 613
rect 2970 606 2973 613
rect 2442 603 2452 606
rect 2474 603 2516 606
rect 2532 603 2557 606
rect 2562 603 2572 606
rect 2602 603 2628 606
rect 2644 603 2661 606
rect 2666 603 2692 606
rect 2722 603 2740 606
rect 2762 603 2788 606
rect 2890 603 2916 606
rect 2970 603 3020 606
rect 3090 603 3116 606
rect 3138 603 3164 606
rect 3194 603 3252 606
rect 3346 603 3380 606
rect 3396 603 3413 606
rect 2722 593 2732 596
rect 2746 593 2780 596
rect 242 583 269 586
rect 38 567 3466 573
rect 578 543 612 546
rect 1642 543 1652 546
rect 1970 543 2004 546
rect 2330 543 2348 546
rect 2554 543 2573 546
rect 90 533 100 536
rect 116 533 133 536
rect 130 526 133 533
rect 178 533 212 536
rect 284 533 317 536
rect 410 533 428 536
rect 466 533 492 536
rect 562 533 572 536
rect 620 533 637 536
rect 660 533 685 536
rect 794 533 820 536
rect 866 533 876 536
rect 914 533 925 536
rect 954 533 996 536
rect 1012 533 1053 536
rect 1074 533 1108 536
rect 1154 533 1164 536
rect 1202 533 1220 536
rect 1266 533 1300 536
rect 1378 533 1396 536
rect 1442 533 1460 536
rect 1476 533 1485 536
rect 178 526 181 533
rect 914 526 917 533
rect 130 523 181 526
rect 194 523 204 526
rect 250 523 268 526
rect 346 523 357 526
rect 364 523 373 526
rect 388 523 397 526
rect 436 523 445 526
rect 452 523 477 526
rect 514 523 556 526
rect 844 523 861 526
rect 900 523 917 526
rect 1042 523 1068 526
rect 1138 523 1172 526
rect 1218 523 1228 526
rect 1252 523 1269 526
rect 1290 523 1308 526
rect 1356 523 1381 526
rect 1420 523 1437 526
rect 156 513 181 516
rect 346 515 349 523
rect 1514 516 1517 536
rect 1554 533 1564 536
rect 1594 533 1604 536
rect 1628 533 1653 536
rect 1690 533 1700 536
rect 1802 533 1820 536
rect 1836 533 1845 536
rect 1930 533 1940 536
rect 2042 533 2076 536
rect 1554 516 1557 533
rect 1572 523 1605 526
rect 1682 523 1708 526
rect 1802 516 1805 533
rect 2098 526 2101 534
rect 2114 533 2148 536
rect 2202 533 2212 536
rect 2242 533 2276 536
rect 2386 533 2396 536
rect 2490 533 2500 536
rect 2554 526 2557 543
rect 2570 533 2580 536
rect 2602 533 2620 536
rect 2714 533 2732 536
rect 2746 533 2788 536
rect 2794 533 2804 536
rect 2826 533 2860 536
rect 3124 533 3141 536
rect 3154 533 3172 536
rect 3258 533 3284 536
rect 3306 526 3309 534
rect 3322 533 3332 536
rect 3356 533 3365 536
rect 3370 533 3396 536
rect 3420 533 3437 536
rect 1914 523 1932 526
rect 2026 523 2036 526
rect 2084 523 2101 526
rect 2108 523 2149 526
rect 2186 523 2204 526
rect 2236 523 2261 526
rect 2274 523 2284 526
rect 2370 523 2388 526
rect 2426 523 2468 526
rect 2490 523 2508 526
rect 2548 523 2557 526
rect 2562 523 2588 526
rect 2610 523 2628 526
rect 2740 523 2781 526
rect 2802 523 2812 526
rect 2818 523 2868 526
rect 2900 523 2909 526
rect 2956 523 2973 526
rect 3084 523 3093 526
rect 3130 523 3180 526
rect 3202 523 3228 526
rect 3274 523 3292 526
rect 3306 523 3333 526
rect 3354 523 3404 526
rect 690 513 700 516
rect 724 513 733 516
rect 1034 513 1053 516
rect 1076 513 1085 516
rect 1180 513 1189 516
rect 1236 513 1245 516
rect 1316 513 1325 516
rect 1514 513 1524 516
rect 1548 513 1557 516
rect 1628 513 1637 516
rect 1724 513 1749 516
rect 1756 513 1765 516
rect 1780 513 1805 516
rect 1900 513 1925 516
rect 2172 513 2197 516
rect 2308 513 2341 516
rect 2476 513 2501 516
rect 2516 513 2533 516
rect 2636 513 2645 516
rect 2684 513 2693 516
rect 3124 513 3149 516
rect 3196 513 3213 516
rect 3244 513 3253 516
rect 3420 513 3429 516
rect 674 503 716 506
rect 746 503 772 506
rect 1498 503 1540 506
rect 1730 503 1772 506
rect 1850 503 1892 506
rect 14 467 3490 473
rect 1802 453 1821 456
rect 282 433 324 436
rect 506 433 524 436
rect 132 423 157 426
rect 276 423 301 426
rect 332 423 365 426
rect 388 423 397 426
rect 466 423 508 426
rect 532 423 541 426
rect 916 423 949 426
rect 1052 423 1077 426
rect 1132 423 1141 426
rect 1460 423 1469 426
rect 146 413 180 416
rect 210 406 213 415
rect 218 413 268 416
rect 380 413 421 416
rect 650 406 653 415
rect 658 413 708 416
rect 740 413 757 416
rect 866 413 876 416
rect 898 413 908 416
rect 1010 413 1044 416
rect 1084 413 1101 416
rect 1124 413 1180 416
rect 1242 413 1260 416
rect 1266 413 1308 416
rect 1332 413 1365 416
rect 1428 413 1437 416
rect 178 403 188 406
rect 210 403 229 406
rect 338 403 372 406
rect 410 403 436 406
rect 538 403 572 406
rect 650 403 685 406
rect 738 403 780 406
rect 1002 403 1036 406
rect 1050 403 1076 406
rect 1202 403 1220 406
rect 1324 403 1357 406
rect 1442 405 1445 416
rect 1452 413 1508 416
rect 1522 413 1549 416
rect 1626 413 1644 416
rect 1482 403 1500 406
rect 1522 405 1525 413
rect 1538 403 1556 406
rect 1570 403 1588 406
rect 1660 403 1669 406
rect 1714 405 1717 436
rect 2674 433 2724 436
rect 1844 423 1869 426
rect 1900 423 1917 426
rect 2300 423 2309 426
rect 2468 423 2501 426
rect 2682 423 2708 426
rect 1794 413 1836 416
rect 1922 413 1940 416
rect 1986 413 2020 416
rect 2034 413 2044 416
rect 2076 413 2085 416
rect 2132 413 2149 416
rect 2170 413 2204 416
rect 2250 413 2292 416
rect 2388 413 2421 416
rect 2460 413 2477 416
rect 2538 413 2548 416
rect 2554 413 2612 416
rect 2618 413 2628 416
rect 2634 413 2652 416
rect 2738 413 2748 416
rect 2836 413 2853 416
rect 2956 413 2981 416
rect 3148 413 3173 416
rect 3420 413 3429 416
rect 1796 403 1821 406
rect 1850 403 1876 406
rect 1964 403 2005 406
rect 2026 403 2052 406
rect 2068 403 2077 406
rect 2106 403 2124 406
rect 2138 403 2148 406
rect 2162 403 2212 406
rect 2258 403 2284 406
rect 2362 403 2380 406
rect 2394 403 2420 406
rect 2442 403 2452 406
rect 2466 403 2516 406
rect 3026 403 3044 406
rect 3076 403 3085 406
rect 546 393 564 396
rect 1330 393 1364 396
rect 1530 393 1548 396
rect 38 367 3466 373
rect 850 343 860 346
rect 1370 336 1373 356
rect 82 333 92 336
rect 122 333 156 336
rect 202 333 228 336
rect 274 333 340 336
rect 386 333 404 336
rect 434 333 484 336
rect 500 333 517 336
rect 658 333 708 336
rect 858 333 868 336
rect 874 333 916 336
rect 938 333 972 336
rect 1082 333 1108 336
rect 180 323 229 326
rect 250 323 268 326
rect 274 323 277 333
rect 386 326 389 333
rect 514 326 517 333
rect 364 323 389 326
rect 442 323 476 326
rect 514 323 532 326
rect 604 323 628 326
rect 650 323 725 326
rect 924 323 957 326
rect 1082 316 1085 333
rect 1130 325 1133 336
rect 1282 333 1308 336
rect 1324 333 1365 336
rect 1370 333 1380 336
rect 1394 333 1404 336
rect 1482 333 1493 336
rect 1602 333 1612 336
rect 1628 333 1645 336
rect 1706 333 1732 336
rect 1754 333 1788 336
rect 1802 333 1836 336
rect 1962 333 1972 336
rect 2066 333 2084 336
rect 2098 333 2156 336
rect 2178 333 2204 336
rect 2218 333 2276 336
rect 1282 316 1285 333
rect 1362 326 1365 333
rect 1482 326 1485 333
rect 1706 326 1709 333
rect 2298 326 2301 335
rect 2324 333 2381 336
rect 2402 333 2412 336
rect 2474 333 2492 336
rect 2514 333 2549 336
rect 1362 323 1388 326
rect 1402 323 1412 326
rect 1436 323 1485 326
rect 1586 323 1604 326
rect 1668 323 1709 326
rect 1714 323 1724 326
rect 1770 323 1796 326
rect 1946 323 2021 326
rect 2058 323 2092 326
rect 2186 323 2212 326
rect 2284 323 2301 326
rect 2330 323 2396 326
rect 2402 323 2420 326
rect 2442 323 2484 326
rect 2514 325 2517 333
rect 116 313 141 316
rect 276 313 325 316
rect 1002 313 1044 316
rect 1068 313 1085 316
rect 1162 313 1180 316
rect 1204 313 1221 316
rect 1226 313 1236 316
rect 1260 313 1285 316
rect 1676 313 1709 316
rect 1226 306 1229 313
rect 1714 306 1717 323
rect 1860 313 1901 316
rect 2060 313 2077 316
rect 2100 313 2141 316
rect 2220 313 2277 316
rect 2330 313 2333 323
rect 2404 313 2413 316
rect 2428 313 2437 316
rect 2554 313 2564 316
rect 2602 313 2628 316
rect 1050 303 1060 306
rect 1138 303 1196 306
rect 1210 303 1229 306
rect 1690 303 1717 306
rect 2138 303 2141 313
rect 2554 293 2557 313
rect 2634 306 2637 325
rect 2658 313 2692 316
rect 2722 313 2756 316
rect 2762 306 2765 325
rect 2884 323 2909 326
rect 3012 323 3037 326
rect 3124 323 3149 326
rect 3252 323 3269 326
rect 3364 323 3389 326
rect 2602 303 2637 306
rect 2674 303 2708 306
rect 2730 303 2765 306
rect 14 267 3490 273
rect 386 233 428 236
rect 906 233 925 236
rect 946 233 996 236
rect 2338 233 2388 236
rect 2402 233 2452 236
rect 2626 233 2669 236
rect 906 226 909 233
rect 244 223 261 226
rect 322 223 356 226
rect 394 223 412 226
rect 484 223 517 226
rect 668 223 685 226
rect 812 223 829 226
rect 900 223 909 226
rect 954 223 980 226
rect 1354 223 1388 226
rect 2330 223 2372 226
rect 2426 223 2436 226
rect 2460 223 2477 226
rect 2562 223 2596 226
rect 2626 223 2660 226
rect 108 213 117 216
rect 130 213 140 216
rect 442 213 476 216
rect 538 213 589 216
rect 596 213 629 216
rect 724 213 757 216
rect 762 213 772 216
rect 810 213 836 216
rect 1010 213 1044 216
rect 1050 213 1084 216
rect 1098 213 1124 216
rect 1156 213 1165 216
rect 1170 213 1196 216
rect 1306 213 1316 216
rect 100 203 109 206
rect 122 203 148 206
rect 164 203 197 206
rect 274 203 292 206
rect 308 203 349 206
rect 442 203 468 206
rect 586 205 589 213
rect 626 206 629 213
rect 746 206 749 213
rect 1474 206 1477 215
rect 1482 213 1524 216
rect 1546 213 1564 216
rect 1586 213 1596 216
rect 1628 213 1637 216
rect 1676 213 1685 216
rect 1692 213 1709 216
rect 1954 213 1964 216
rect 1996 213 2028 216
rect 2090 213 2124 216
rect 2194 213 2212 216
rect 2266 213 2292 216
rect 2324 213 2349 216
rect 2466 213 2500 216
rect 2506 213 2540 216
rect 2556 213 2589 216
rect 2666 215 2669 233
rect 3170 233 3189 236
rect 2772 223 2781 226
rect 2924 223 2933 226
rect 3170 216 3173 233
rect 2690 213 2700 216
rect 2778 213 2796 216
rect 2860 213 2893 216
rect 2922 213 2972 216
rect 3012 213 3061 216
rect 3132 213 3173 216
rect 3186 215 3189 233
rect 3220 213 3229 216
rect 3300 213 3325 216
rect 3412 213 3437 216
rect 626 203 644 206
rect 716 203 725 206
rect 746 203 764 206
rect 778 203 796 206
rect 850 203 884 206
rect 1018 203 1036 206
rect 1058 203 1076 206
rect 1090 203 1132 206
rect 1154 203 1188 206
rect 1282 203 1324 206
rect 1418 203 1452 206
rect 1474 203 1509 206
rect 1658 203 1668 206
rect 1682 205 1685 213
rect 1698 203 1764 206
rect 1802 203 1860 206
rect 2002 203 2020 206
rect 2042 203 2125 206
rect 2210 203 2220 206
rect 2316 203 2365 206
rect 2924 203 2941 206
rect 2034 193 2068 196
rect 3058 195 3061 213
rect 3068 203 3093 206
rect 3148 203 3165 206
rect 3362 203 3380 206
rect 38 167 3466 173
rect 154 136 157 146
rect 1370 143 1404 146
rect 1826 143 1836 146
rect 154 133 180 136
rect 226 133 237 136
rect 260 133 317 136
rect 426 133 436 136
rect 562 133 572 136
rect 602 133 612 136
rect 642 133 660 136
rect 714 133 725 136
rect 748 133 820 136
rect 842 133 876 136
rect 890 133 932 136
rect 948 133 1005 136
rect 1042 133 1084 136
rect 1108 133 1117 136
rect 1138 133 1180 136
rect 1196 133 1221 136
rect 1268 133 1293 136
rect 1314 133 1340 136
rect 1364 133 1397 136
rect 1402 133 1412 136
rect 1474 133 1492 136
rect 1498 133 1509 136
rect 1738 133 1772 136
rect 1834 133 1844 136
rect 1850 133 1884 136
rect 1978 133 2004 136
rect 188 123 205 126
rect 226 116 229 133
rect 602 126 605 133
rect 642 126 645 133
rect 274 123 324 126
rect 444 123 493 126
rect 538 123 605 126
rect 620 123 645 126
rect 714 116 717 133
rect 1506 126 1509 133
rect 2090 126 2093 135
rect 2106 133 2140 136
rect 2282 133 2324 136
rect 2426 133 2484 136
rect 2804 133 2837 136
rect 2890 133 2940 136
rect 3002 126 3005 134
rect 3058 126 3061 134
rect 762 123 812 126
rect 844 123 861 126
rect 866 123 884 126
rect 898 123 924 126
rect 962 123 1004 126
rect 1058 123 1092 126
rect 1132 123 1165 126
rect 1210 123 1252 126
rect 1308 123 1348 126
rect 1506 123 1524 126
rect 1612 123 1629 126
rect 1738 123 1764 126
rect 1852 123 1861 126
rect 1892 123 1901 126
rect 1914 123 1956 126
rect 1986 123 2012 126
rect 2076 123 2093 126
rect 2148 123 2181 126
rect 2282 123 2316 126
rect 2362 123 2396 126
rect 2428 123 2437 126
rect 196 113 229 116
rect 684 113 717 116
rect 892 113 917 116
rect 1532 113 1565 116
rect 1618 113 1652 116
rect 1676 113 1701 116
rect 1708 113 1717 116
rect 1732 113 1757 116
rect 1972 113 1989 116
rect 2028 113 2061 116
rect 2170 113 2188 116
rect 2226 113 2252 116
rect 2276 113 2309 116
rect 2578 113 2588 116
rect 2594 106 2597 125
rect 2618 123 2660 126
rect 2732 123 2741 126
rect 2884 123 2933 126
rect 2970 123 3005 126
rect 3012 123 3061 126
rect 3074 133 3084 136
rect 3146 133 3172 136
rect 3242 133 3252 136
rect 2740 113 2749 116
rect 2892 113 2901 116
rect 3074 115 3077 133
rect 3314 126 3317 136
rect 3370 133 3412 136
rect 3426 126 3429 136
rect 3218 123 3236 126
rect 3242 123 3317 126
rect 3346 123 3364 126
rect 3370 123 3429 126
rect 3218 116 3221 123
rect 3196 113 3221 116
rect 3346 115 3349 123
rect 3372 113 3381 116
rect 1682 103 1724 106
rect 2162 103 2204 106
rect 2218 103 2268 106
rect 2562 103 2597 106
rect 14 67 3490 73
rect 38 37 3466 57
rect 14 13 3490 33
<< metal2 >>
rect 14 13 34 3327
rect 38 37 58 3303
rect 66 2976 69 3146
rect 90 3003 93 3156
rect 170 3153 173 3206
rect 218 3173 221 3216
rect 282 3186 285 3216
rect 306 3186 309 3206
rect 282 3183 293 3186
rect 194 3163 229 3166
rect 138 3123 141 3136
rect 138 3003 141 3016
rect 162 3013 189 3016
rect 66 2973 77 2976
rect 74 2866 77 2973
rect 138 2943 141 2996
rect 162 2943 165 3013
rect 194 3003 197 3163
rect 226 3146 229 3163
rect 226 3143 261 3146
rect 226 3133 229 3143
rect 242 3133 253 3136
rect 258 3133 261 3143
rect 210 3003 221 3006
rect 226 2993 229 3126
rect 266 3076 269 3156
rect 274 3083 277 3116
rect 250 3073 269 3076
rect 234 3023 237 3046
rect 250 2993 253 3073
rect 282 3066 285 3136
rect 290 3106 293 3183
rect 298 3183 309 3186
rect 298 3153 301 3183
rect 306 3133 309 3176
rect 330 3133 333 3206
rect 322 3113 333 3116
rect 290 3103 297 3106
rect 278 3063 285 3066
rect 278 2976 281 3063
rect 294 3056 297 3103
rect 194 2943 197 2976
rect 274 2973 281 2976
rect 290 3053 297 3056
rect 290 2973 293 3053
rect 66 2863 77 2866
rect 66 2756 69 2863
rect 106 2813 109 2926
rect 154 2896 157 2936
rect 162 2923 213 2926
rect 210 2913 213 2923
rect 154 2893 173 2896
rect 170 2826 173 2893
rect 170 2823 177 2826
rect 82 2776 85 2806
rect 82 2773 141 2776
rect 66 2753 85 2756
rect 82 2646 85 2753
rect 138 2733 141 2773
rect 66 2643 85 2646
rect 66 2626 69 2643
rect 162 2626 165 2816
rect 174 2746 177 2823
rect 218 2813 221 2936
rect 258 2933 261 2946
rect 266 2923 269 2936
rect 274 2933 277 2973
rect 298 2933 301 3016
rect 306 2933 309 2946
rect 330 2943 333 3016
rect 338 2956 341 3156
rect 354 3136 357 3216
rect 386 3203 389 3216
rect 418 3193 421 3206
rect 346 3123 349 3136
rect 354 3133 373 3136
rect 354 3013 357 3126
rect 410 3113 413 3136
rect 418 3133 421 3186
rect 434 3123 437 3136
rect 458 3133 461 3216
rect 498 3183 501 3216
rect 506 3143 509 3216
rect 554 3213 557 3226
rect 610 3223 613 3246
rect 618 3216 621 3236
rect 530 3193 533 3206
rect 554 3156 557 3206
rect 562 3193 565 3206
rect 514 3153 557 3156
rect 570 3153 573 3216
rect 514 3133 517 3153
rect 586 3146 589 3206
rect 402 3013 405 3026
rect 354 2976 357 3006
rect 354 2973 373 2976
rect 338 2953 349 2956
rect 298 2903 301 2916
rect 322 2863 325 2926
rect 194 2773 197 2806
rect 274 2756 277 2816
rect 330 2813 333 2936
rect 346 2846 349 2953
rect 370 2893 373 2973
rect 338 2843 349 2846
rect 306 2776 309 2806
rect 338 2786 341 2843
rect 170 2743 177 2746
rect 266 2753 277 2756
rect 298 2773 309 2776
rect 330 2783 341 2786
rect 170 2723 173 2743
rect 66 2623 101 2626
rect 66 2576 69 2623
rect 82 2593 85 2616
rect 98 2613 101 2623
rect 146 2623 165 2626
rect 90 2596 93 2606
rect 138 2603 141 2616
rect 146 2613 149 2623
rect 90 2593 125 2596
rect 122 2583 125 2593
rect 66 2573 77 2576
rect 74 2476 77 2573
rect 154 2543 157 2616
rect 170 2596 173 2626
rect 178 2603 181 2616
rect 218 2613 221 2726
rect 266 2706 269 2753
rect 298 2733 301 2773
rect 330 2716 333 2783
rect 346 2723 349 2826
rect 386 2736 389 2816
rect 402 2793 405 3006
rect 442 2996 445 3126
rect 466 3026 469 3126
rect 498 3103 501 3116
rect 506 3066 509 3126
rect 522 3123 525 3136
rect 546 3133 549 3146
rect 554 3143 589 3146
rect 554 3133 557 3143
rect 498 3063 509 3066
rect 538 3086 541 3126
rect 546 3093 549 3126
rect 562 3103 565 3126
rect 578 3086 581 3126
rect 586 3093 589 3126
rect 538 3083 581 3086
rect 466 3023 485 3026
rect 466 3003 469 3023
rect 442 2993 453 2996
rect 418 2923 421 2946
rect 450 2856 453 2993
rect 450 2853 469 2856
rect 434 2833 453 2836
rect 434 2813 437 2833
rect 434 2786 437 2806
rect 442 2803 445 2826
rect 450 2816 453 2833
rect 458 2816 461 2826
rect 450 2813 461 2816
rect 442 2793 453 2796
rect 434 2783 445 2786
rect 450 2783 453 2793
rect 378 2733 389 2736
rect 330 2713 341 2716
rect 266 2703 277 2706
rect 166 2593 173 2596
rect 66 2473 77 2476
rect 66 2043 69 2473
rect 74 2436 77 2456
rect 74 2433 81 2436
rect 78 2366 81 2433
rect 98 2376 101 2406
rect 74 2363 81 2366
rect 90 2373 101 2376
rect 74 2296 77 2363
rect 90 2333 93 2373
rect 130 2353 133 2416
rect 138 2393 141 2536
rect 166 2366 169 2593
rect 162 2363 169 2366
rect 74 2293 85 2296
rect 82 2236 85 2293
rect 78 2233 85 2236
rect 78 2156 81 2233
rect 90 2203 93 2216
rect 74 2153 81 2156
rect 66 1523 69 2036
rect 66 983 69 1446
rect 74 1316 77 2153
rect 114 2146 117 2216
rect 122 2203 125 2326
rect 162 2316 165 2363
rect 178 2323 181 2596
rect 202 2566 205 2606
rect 202 2563 209 2566
rect 186 2476 189 2526
rect 206 2486 209 2563
rect 218 2523 221 2546
rect 234 2503 237 2606
rect 242 2576 245 2646
rect 250 2603 253 2616
rect 274 2613 277 2703
rect 298 2643 325 2646
rect 338 2643 341 2713
rect 378 2686 381 2733
rect 354 2683 381 2686
rect 242 2573 261 2576
rect 242 2546 245 2566
rect 242 2543 249 2546
rect 246 2496 249 2543
rect 202 2483 209 2486
rect 242 2493 249 2496
rect 186 2473 193 2476
rect 190 2316 193 2473
rect 202 2413 205 2483
rect 218 2393 221 2406
rect 162 2313 173 2316
rect 170 2286 173 2313
rect 162 2283 173 2286
rect 186 2313 193 2316
rect 130 2203 133 2216
rect 146 2156 149 2226
rect 162 2213 165 2283
rect 170 2223 181 2226
rect 146 2153 153 2156
rect 114 2143 125 2146
rect 82 2123 85 2136
rect 90 2123 101 2126
rect 98 2113 101 2123
rect 82 1946 85 2046
rect 90 1956 93 2096
rect 106 2033 109 2126
rect 114 2103 117 2136
rect 122 2026 125 2143
rect 130 2073 133 2126
rect 138 2093 141 2146
rect 106 2013 109 2026
rect 122 2023 133 2026
rect 98 2003 109 2006
rect 90 1953 101 1956
rect 82 1943 93 1946
rect 82 1913 85 1936
rect 82 1743 85 1906
rect 90 1736 93 1943
rect 98 1933 101 1953
rect 106 1933 109 1946
rect 98 1803 101 1926
rect 106 1913 109 1926
rect 114 1923 117 2006
rect 122 1963 125 2016
rect 130 1956 133 2023
rect 122 1953 133 1956
rect 122 1906 125 1953
rect 118 1903 125 1906
rect 82 1643 85 1736
rect 90 1733 101 1736
rect 106 1733 109 1816
rect 118 1746 121 1903
rect 118 1743 125 1746
rect 130 1743 133 1946
rect 138 1773 141 2086
rect 150 2036 153 2153
rect 150 2033 157 2036
rect 146 2003 149 2026
rect 146 1913 149 1926
rect 90 1643 93 1726
rect 98 1706 101 1733
rect 106 1723 117 1726
rect 122 1706 125 1743
rect 98 1703 105 1706
rect 102 1636 105 1703
rect 82 1633 93 1636
rect 98 1633 105 1636
rect 114 1703 125 1706
rect 98 1616 101 1633
rect 114 1623 117 1703
rect 90 1613 101 1616
rect 106 1613 117 1616
rect 82 1533 85 1606
rect 90 1563 93 1613
rect 90 1523 93 1546
rect 98 1533 101 1606
rect 106 1516 109 1606
rect 114 1546 117 1596
rect 122 1566 125 1616
rect 130 1613 133 1736
rect 138 1593 141 1766
rect 146 1613 149 1826
rect 122 1563 133 1566
rect 130 1553 133 1563
rect 114 1543 121 1546
rect 94 1513 109 1516
rect 82 1383 85 1466
rect 94 1436 97 1513
rect 90 1433 97 1436
rect 82 1333 85 1346
rect 74 1313 81 1316
rect 78 1226 81 1313
rect 74 1223 81 1226
rect 74 1066 77 1223
rect 90 1216 93 1433
rect 106 1423 109 1506
rect 118 1436 121 1543
rect 114 1433 121 1436
rect 114 1416 117 1433
rect 98 1413 109 1416
rect 114 1413 125 1416
rect 114 1406 117 1413
rect 98 1393 101 1406
rect 106 1403 117 1406
rect 98 1313 101 1386
rect 106 1316 109 1403
rect 114 1323 117 1396
rect 122 1336 125 1406
rect 130 1343 133 1546
rect 138 1513 141 1526
rect 122 1333 133 1336
rect 106 1313 117 1316
rect 114 1236 117 1313
rect 114 1233 125 1236
rect 90 1213 97 1216
rect 82 1103 85 1206
rect 94 1146 97 1213
rect 106 1203 109 1216
rect 90 1143 97 1146
rect 82 1083 85 1096
rect 74 1063 81 1066
rect 78 986 81 1063
rect 74 983 81 986
rect 74 966 77 983
rect 70 963 77 966
rect 70 756 73 963
rect 82 943 85 956
rect 82 813 85 936
rect 70 753 77 756
rect 82 753 85 806
rect 66 713 69 736
rect 66 303 69 706
rect 74 343 77 753
rect 82 333 85 736
rect 90 696 93 1143
rect 106 1123 109 1146
rect 114 1106 117 1136
rect 106 1103 117 1106
rect 106 1013 109 1103
rect 98 1003 117 1006
rect 98 906 101 996
rect 106 923 109 1003
rect 114 933 117 986
rect 98 903 105 906
rect 102 776 105 903
rect 114 803 117 916
rect 98 773 105 776
rect 98 716 101 773
rect 106 723 109 756
rect 114 733 117 746
rect 98 713 113 716
rect 90 693 101 696
rect 98 626 101 693
rect 90 623 101 626
rect 110 626 113 713
rect 110 623 117 626
rect 90 556 93 623
rect 98 603 109 606
rect 90 553 101 556
rect 90 533 93 546
rect 98 526 101 553
rect 90 523 101 526
rect 106 523 109 603
rect 90 506 93 523
rect 114 516 117 623
rect 106 513 117 516
rect 90 503 97 506
rect 94 346 97 503
rect 90 343 97 346
rect 90 293 93 343
rect 98 233 101 326
rect 106 203 109 513
rect 122 506 125 1233
rect 130 1203 133 1333
rect 130 1133 133 1146
rect 130 1103 133 1126
rect 130 943 133 1076
rect 138 993 141 1456
rect 146 1413 149 1536
rect 154 1523 157 2033
rect 162 1816 165 2126
rect 170 2106 173 2223
rect 178 2123 181 2216
rect 186 2203 189 2313
rect 202 2216 205 2336
rect 226 2323 229 2366
rect 242 2323 245 2493
rect 258 2466 261 2573
rect 282 2556 285 2616
rect 298 2603 301 2643
rect 306 2563 309 2636
rect 314 2593 317 2606
rect 322 2603 325 2643
rect 354 2613 357 2683
rect 274 2553 285 2556
rect 274 2506 277 2553
rect 298 2523 301 2536
rect 362 2526 365 2616
rect 378 2536 381 2646
rect 402 2613 405 2726
rect 418 2666 421 2776
rect 442 2723 445 2783
rect 418 2663 437 2666
rect 386 2553 389 2606
rect 410 2576 413 2616
rect 434 2603 437 2663
rect 458 2613 461 2806
rect 466 2793 469 2853
rect 474 2783 477 3016
rect 482 2986 485 3023
rect 490 3003 493 3026
rect 498 2996 501 3063
rect 506 3016 509 3026
rect 538 3016 541 3083
rect 594 3046 597 3216
rect 610 3213 621 3216
rect 626 3213 637 3216
rect 650 3213 653 3276
rect 658 3223 661 3236
rect 658 3213 677 3216
rect 682 3213 685 3246
rect 802 3216 805 3236
rect 714 3213 725 3216
rect 746 3213 805 3216
rect 586 3043 597 3046
rect 506 3013 533 3016
rect 538 3013 549 3016
rect 498 2993 509 2996
rect 522 2993 525 3006
rect 482 2983 501 2986
rect 498 2916 501 2983
rect 506 2933 509 2993
rect 522 2933 525 2946
rect 490 2913 501 2916
rect 490 2846 493 2913
rect 490 2843 501 2846
rect 482 2813 485 2826
rect 498 2813 501 2843
rect 506 2743 509 2926
rect 514 2923 525 2926
rect 538 2923 541 3006
rect 546 2963 549 3013
rect 554 2976 557 3026
rect 586 3023 589 3043
rect 594 3023 597 3036
rect 602 3016 605 3196
rect 610 3133 613 3213
rect 658 3206 661 3213
rect 626 3203 661 3206
rect 634 3173 653 3176
rect 618 3123 621 3136
rect 634 3133 637 3173
rect 642 3133 645 3166
rect 626 3083 629 3126
rect 642 3106 645 3126
rect 634 3103 645 3106
rect 650 3103 653 3173
rect 650 3066 653 3086
rect 562 2986 565 3016
rect 586 3013 605 3016
rect 610 3063 653 3066
rect 610 3013 613 3063
rect 642 3023 653 3026
rect 586 3006 589 3013
rect 570 3003 589 3006
rect 594 2993 597 3006
rect 602 3003 605 3013
rect 626 2986 629 3006
rect 562 2983 573 2986
rect 554 2973 565 2976
rect 498 2626 501 2726
rect 514 2643 517 2923
rect 522 2913 533 2916
rect 530 2753 533 2896
rect 554 2776 557 2973
rect 538 2773 557 2776
rect 498 2623 509 2626
rect 410 2573 461 2576
rect 378 2533 389 2536
rect 410 2533 413 2573
rect 274 2503 301 2506
rect 254 2463 261 2466
rect 254 2386 257 2463
rect 250 2383 257 2386
rect 250 2363 253 2383
rect 250 2333 253 2356
rect 266 2336 269 2416
rect 298 2413 301 2503
rect 346 2486 349 2526
rect 362 2523 381 2526
rect 346 2483 365 2486
rect 330 2403 333 2416
rect 354 2376 357 2476
rect 338 2373 357 2376
rect 258 2323 261 2336
rect 266 2333 285 2336
rect 298 2323 301 2336
rect 242 2256 245 2316
rect 226 2253 245 2256
rect 194 2213 205 2216
rect 210 2143 213 2246
rect 186 2133 221 2136
rect 194 2113 197 2126
rect 170 2103 177 2106
rect 174 1956 177 2103
rect 170 1953 177 1956
rect 170 1896 173 1953
rect 178 1913 181 1936
rect 186 1923 189 2026
rect 194 1996 197 2016
rect 202 2003 205 2126
rect 210 2003 213 2126
rect 218 2093 221 2133
rect 218 2013 221 2026
rect 218 1996 221 2006
rect 194 1993 221 1996
rect 170 1893 181 1896
rect 162 1813 173 1816
rect 178 1746 181 1893
rect 194 1763 197 1966
rect 202 1923 205 1986
rect 226 1946 229 2253
rect 258 2223 277 2226
rect 258 2216 261 2223
rect 250 2213 261 2216
rect 266 2206 269 2216
rect 274 2213 277 2223
rect 234 2043 237 2136
rect 242 2116 245 2156
rect 258 2146 261 2206
rect 266 2203 277 2206
rect 266 2153 269 2203
rect 258 2143 277 2146
rect 258 2136 261 2143
rect 250 2133 261 2136
rect 242 2113 249 2116
rect 246 2036 249 2113
rect 258 2103 261 2126
rect 266 2113 269 2136
rect 274 2133 277 2143
rect 274 2053 277 2126
rect 282 2036 285 2316
rect 242 2033 249 2036
rect 274 2033 285 2036
rect 234 2013 237 2026
rect 242 1963 245 2033
rect 218 1943 229 1946
rect 234 1953 245 1956
rect 210 1903 213 1926
rect 202 1793 205 1806
rect 170 1743 181 1746
rect 162 1713 165 1726
rect 154 1453 157 1506
rect 154 1356 157 1436
rect 162 1386 165 1706
rect 170 1443 173 1743
rect 178 1693 181 1736
rect 194 1723 197 1736
rect 178 1416 181 1656
rect 194 1646 197 1716
rect 186 1643 197 1646
rect 186 1493 189 1643
rect 202 1636 205 1776
rect 210 1723 213 1806
rect 218 1723 221 1943
rect 226 1923 229 1936
rect 234 1933 237 1953
rect 226 1826 229 1916
rect 234 1903 237 1916
rect 242 1876 245 1946
rect 250 1936 253 2016
rect 258 1943 261 2026
rect 266 2013 269 2026
rect 250 1933 269 1936
rect 250 1903 253 1933
rect 258 1913 261 1926
rect 266 1923 269 1933
rect 242 1873 253 1876
rect 226 1823 237 1826
rect 226 1783 229 1816
rect 234 1716 237 1823
rect 194 1633 205 1636
rect 210 1713 221 1716
rect 226 1713 237 1716
rect 194 1453 197 1633
rect 210 1613 213 1713
rect 202 1603 213 1606
rect 226 1586 229 1713
rect 234 1603 237 1616
rect 226 1583 237 1586
rect 202 1513 205 1526
rect 186 1423 205 1426
rect 170 1393 173 1416
rect 178 1413 189 1416
rect 178 1386 181 1406
rect 162 1383 181 1386
rect 154 1353 165 1356
rect 146 1183 149 1336
rect 154 1323 157 1346
rect 146 1046 149 1146
rect 154 1066 157 1316
rect 162 1203 165 1353
rect 162 1093 165 1136
rect 170 1086 173 1326
rect 186 1233 189 1413
rect 194 1403 197 1423
rect 202 1403 205 1416
rect 210 1413 213 1536
rect 226 1526 229 1576
rect 234 1533 237 1583
rect 242 1533 245 1726
rect 250 1706 253 1873
rect 266 1733 269 1916
rect 274 1803 277 2033
rect 282 1996 285 2026
rect 290 2003 293 2256
rect 298 2023 301 2236
rect 306 2123 309 2156
rect 298 2003 309 2006
rect 282 1993 293 1996
rect 290 1926 293 1993
rect 306 1973 309 2003
rect 314 1946 317 2046
rect 306 1943 317 1946
rect 282 1923 301 1926
rect 282 1803 285 1923
rect 290 1846 293 1916
rect 298 1893 301 1906
rect 290 1843 301 1846
rect 298 1756 301 1843
rect 274 1723 277 1756
rect 282 1753 301 1756
rect 306 1753 309 1943
rect 314 1816 317 1936
rect 322 1913 325 2336
rect 338 2123 341 2373
rect 362 2333 365 2483
rect 386 2456 389 2533
rect 370 2453 389 2456
rect 370 2326 373 2453
rect 378 2343 381 2416
rect 346 2323 373 2326
rect 378 2323 381 2336
rect 354 2293 357 2323
rect 362 2253 365 2316
rect 394 2286 397 2366
rect 402 2303 405 2446
rect 426 2413 429 2526
rect 442 2443 445 2566
rect 450 2533 453 2556
rect 458 2533 461 2573
rect 506 2566 509 2623
rect 490 2563 509 2566
rect 522 2563 525 2606
rect 490 2523 493 2563
rect 530 2546 533 2616
rect 538 2613 541 2773
rect 562 2766 565 2826
rect 554 2763 565 2766
rect 570 2766 573 2983
rect 594 2983 629 2986
rect 634 2983 637 3016
rect 658 3003 661 3203
rect 666 3196 669 3206
rect 674 3203 677 3213
rect 690 3196 693 3206
rect 730 3203 741 3206
rect 746 3196 749 3213
rect 666 3193 693 3196
rect 730 3193 749 3196
rect 754 3193 773 3196
rect 674 3176 677 3193
rect 674 3173 685 3176
rect 666 3113 669 3146
rect 682 3036 685 3173
rect 714 3123 717 3136
rect 666 3013 669 3036
rect 674 3033 685 3036
rect 674 2993 677 3033
rect 682 3013 693 3016
rect 682 3003 693 3006
rect 586 2923 589 2936
rect 594 2933 597 2983
rect 602 2903 605 2926
rect 578 2803 581 2816
rect 570 2763 581 2766
rect 546 2703 549 2736
rect 554 2723 557 2763
rect 562 2633 565 2736
rect 578 2666 581 2763
rect 570 2663 581 2666
rect 570 2623 573 2663
rect 570 2603 573 2616
rect 602 2613 605 2736
rect 610 2723 613 2946
rect 618 2906 621 2966
rect 682 2946 685 3003
rect 698 2983 701 3016
rect 674 2943 685 2946
rect 626 2923 629 2936
rect 634 2923 637 2936
rect 642 2913 645 2926
rect 658 2906 661 2926
rect 674 2916 677 2936
rect 690 2933 693 2946
rect 618 2903 661 2906
rect 670 2913 677 2916
rect 670 2846 673 2913
rect 670 2843 677 2846
rect 618 2803 621 2816
rect 618 2716 621 2746
rect 626 2726 629 2826
rect 634 2733 637 2816
rect 650 2736 653 2816
rect 666 2813 669 2826
rect 674 2813 677 2843
rect 682 2806 685 2926
rect 698 2813 701 2936
rect 706 2896 709 3116
rect 730 3113 733 3193
rect 786 3183 789 3206
rect 746 3133 749 3146
rect 754 3133 765 3136
rect 770 3133 773 3156
rect 714 3013 717 3106
rect 738 3093 741 3126
rect 754 3113 757 3126
rect 770 3076 773 3126
rect 786 3123 789 3136
rect 794 3116 797 3206
rect 802 3203 805 3213
rect 762 3073 773 3076
rect 786 3113 797 3116
rect 722 3003 725 3016
rect 730 3003 733 3056
rect 738 3013 741 3026
rect 746 2993 749 3006
rect 754 2986 757 3006
rect 714 2923 717 2936
rect 722 2933 725 2986
rect 730 2983 757 2986
rect 730 2926 733 2983
rect 762 2976 765 3073
rect 770 3013 773 3066
rect 786 3046 789 3113
rect 802 3053 805 3146
rect 818 3126 821 3186
rect 842 3143 845 3226
rect 882 3223 917 3226
rect 858 3193 861 3216
rect 874 3206 877 3216
rect 882 3213 885 3223
rect 906 3206 909 3216
rect 914 3213 917 3223
rect 874 3203 885 3206
rect 906 3203 917 3206
rect 818 3123 829 3126
rect 778 3043 789 3046
rect 778 2986 781 3043
rect 754 2973 765 2976
rect 774 2983 781 2986
rect 722 2923 733 2926
rect 738 2916 741 2926
rect 714 2913 741 2916
rect 706 2893 717 2896
rect 714 2806 717 2893
rect 730 2813 741 2816
rect 754 2813 757 2973
rect 774 2926 777 2983
rect 786 2933 789 3006
rect 794 2973 797 3006
rect 802 2993 805 3016
rect 810 3003 813 3106
rect 826 3056 829 3123
rect 818 3053 829 3056
rect 850 3056 853 3136
rect 874 3133 877 3203
rect 906 3183 909 3196
rect 882 3136 885 3176
rect 914 3173 917 3203
rect 890 3143 893 3156
rect 882 3133 893 3136
rect 866 3103 869 3126
rect 890 3123 893 3133
rect 898 3116 901 3136
rect 890 3113 901 3116
rect 922 3113 925 3156
rect 890 3096 893 3113
rect 886 3093 893 3096
rect 850 3053 869 3056
rect 818 3006 821 3053
rect 826 3013 829 3026
rect 818 3003 829 3006
rect 834 3003 837 3036
rect 842 3013 845 3026
rect 858 3006 861 3016
rect 842 3003 861 3006
rect 826 2996 829 3003
rect 842 2996 845 3003
rect 826 2993 845 2996
rect 850 2993 861 2996
rect 794 2933 797 2966
rect 774 2923 781 2926
rect 778 2906 781 2923
rect 786 2913 789 2926
rect 794 2906 797 2926
rect 778 2903 797 2906
rect 794 2806 797 2816
rect 658 2803 669 2806
rect 674 2803 693 2806
rect 642 2733 653 2736
rect 626 2723 637 2726
rect 642 2716 645 2733
rect 618 2713 645 2716
rect 674 2636 677 2736
rect 690 2716 693 2803
rect 706 2803 717 2806
rect 706 2723 709 2803
rect 730 2793 733 2806
rect 778 2803 797 2806
rect 802 2803 805 2946
rect 818 2933 821 2986
rect 810 2906 813 2926
rect 826 2913 829 2993
rect 834 2933 837 2946
rect 810 2903 817 2906
rect 814 2846 817 2903
rect 810 2843 817 2846
rect 810 2826 813 2843
rect 810 2823 837 2826
rect 738 2733 741 2756
rect 690 2713 725 2716
rect 658 2633 677 2636
rect 650 2556 653 2616
rect 530 2543 549 2546
rect 514 2523 525 2526
rect 442 2403 445 2416
rect 418 2333 421 2346
rect 426 2323 429 2336
rect 490 2333 493 2416
rect 522 2413 525 2523
rect 530 2506 533 2536
rect 546 2523 549 2543
rect 562 2533 565 2546
rect 570 2543 573 2556
rect 634 2533 637 2556
rect 642 2553 653 2556
rect 530 2503 541 2506
rect 538 2446 541 2503
rect 530 2443 541 2446
rect 530 2356 533 2443
rect 594 2426 597 2496
rect 610 2456 613 2526
rect 626 2463 629 2526
rect 642 2523 645 2553
rect 658 2533 661 2633
rect 674 2603 677 2616
rect 698 2613 701 2706
rect 722 2656 725 2713
rect 718 2653 725 2656
rect 706 2533 709 2646
rect 718 2546 721 2653
rect 778 2636 781 2803
rect 794 2783 797 2803
rect 786 2723 789 2746
rect 810 2646 813 2816
rect 842 2813 845 2926
rect 858 2913 861 2993
rect 866 2943 869 3053
rect 834 2793 837 2806
rect 850 2746 853 2816
rect 858 2803 861 2826
rect 874 2816 877 3086
rect 886 3026 889 3093
rect 886 3023 893 3026
rect 890 3003 893 3023
rect 898 3003 901 3106
rect 930 3103 933 3206
rect 946 3123 949 3216
rect 946 3103 949 3116
rect 906 2976 909 3016
rect 914 3003 917 3086
rect 922 2983 925 3016
rect 930 2976 933 3006
rect 946 3003 949 3016
rect 906 2973 933 2976
rect 906 2953 909 2973
rect 882 2923 893 2926
rect 898 2823 901 2926
rect 914 2883 917 2926
rect 930 2913 933 2946
rect 954 2933 957 3006
rect 938 2906 941 2926
rect 962 2913 965 3226
rect 970 3213 973 3236
rect 986 3216 989 3226
rect 994 3223 1053 3226
rect 986 3213 997 3216
rect 1050 3213 1053 3223
rect 994 3203 1013 3206
rect 970 3126 973 3136
rect 986 3133 989 3186
rect 1010 3133 1013 3146
rect 970 3123 989 3126
rect 1018 3123 1021 3136
rect 1034 3133 1037 3206
rect 1066 3203 1069 3236
rect 1074 3213 1093 3216
rect 1082 3143 1085 3186
rect 1050 3133 1077 3136
rect 986 3073 989 3123
rect 1058 3116 1061 3126
rect 1034 3113 1061 3116
rect 1074 3096 1077 3133
rect 986 3023 997 3026
rect 970 2963 973 3016
rect 1002 3013 1005 3096
rect 1066 3093 1077 3096
rect 1018 3013 1021 3046
rect 1042 3026 1045 3076
rect 1066 3046 1069 3093
rect 1066 3043 1077 3046
rect 1042 3023 1049 3026
rect 978 3003 997 3006
rect 978 2933 981 3003
rect 1010 2993 1013 3006
rect 1018 3003 1029 3006
rect 994 2933 997 2946
rect 1002 2933 1005 2966
rect 874 2813 909 2816
rect 850 2743 885 2746
rect 890 2743 893 2806
rect 898 2783 901 2796
rect 810 2643 821 2646
rect 770 2633 781 2636
rect 754 2556 757 2616
rect 718 2543 725 2546
rect 610 2453 637 2456
rect 586 2423 597 2426
rect 554 2403 557 2416
rect 514 2353 533 2356
rect 514 2326 517 2353
rect 474 2323 517 2326
rect 410 2313 421 2316
rect 410 2296 413 2313
rect 410 2293 421 2296
rect 394 2283 405 2286
rect 386 2223 389 2266
rect 354 2133 357 2146
rect 362 2123 365 2216
rect 370 2213 389 2216
rect 338 2033 341 2116
rect 330 1933 333 2026
rect 346 2023 349 2066
rect 338 2013 349 2016
rect 338 1993 341 2013
rect 354 2006 357 2056
rect 346 2003 357 2006
rect 346 1986 349 2003
rect 338 1983 349 1986
rect 338 1846 341 1983
rect 346 1926 349 1956
rect 354 1933 357 1996
rect 362 1953 365 2106
rect 346 1923 357 1926
rect 362 1923 365 1936
rect 354 1856 357 1923
rect 354 1853 361 1856
rect 338 1843 349 1846
rect 322 1823 341 1826
rect 314 1813 325 1816
rect 250 1703 261 1706
rect 258 1626 261 1703
rect 282 1683 285 1753
rect 298 1743 317 1746
rect 290 1733 301 1736
rect 250 1623 261 1626
rect 250 1583 253 1623
rect 290 1613 293 1733
rect 298 1653 301 1726
rect 314 1723 317 1743
rect 322 1716 325 1813
rect 338 1793 341 1823
rect 346 1723 349 1843
rect 358 1766 361 1853
rect 354 1763 361 1766
rect 314 1713 325 1716
rect 298 1606 301 1636
rect 218 1423 221 1526
rect 226 1523 237 1526
rect 226 1416 229 1506
rect 234 1463 237 1523
rect 250 1513 253 1556
rect 258 1533 269 1536
rect 258 1523 261 1533
rect 266 1493 269 1506
rect 274 1503 277 1606
rect 282 1543 285 1606
rect 290 1603 301 1606
rect 282 1496 285 1526
rect 274 1493 285 1496
rect 218 1413 229 1416
rect 178 1223 205 1226
rect 178 1103 181 1216
rect 186 1096 189 1176
rect 194 1116 197 1126
rect 202 1123 205 1223
rect 210 1213 213 1336
rect 218 1333 221 1413
rect 234 1376 237 1456
rect 230 1373 237 1376
rect 230 1316 233 1373
rect 226 1313 233 1316
rect 226 1226 229 1313
rect 218 1223 229 1226
rect 218 1206 221 1223
rect 210 1203 221 1206
rect 210 1123 213 1203
rect 234 1173 237 1216
rect 218 1123 221 1136
rect 226 1116 229 1126
rect 194 1113 229 1116
rect 162 1083 173 1086
rect 154 1063 165 1066
rect 146 1043 153 1046
rect 150 986 153 1043
rect 146 983 153 986
rect 138 896 141 936
rect 130 893 141 896
rect 130 736 133 893
rect 138 823 141 836
rect 130 733 141 736
rect 130 713 133 726
rect 146 703 149 983
rect 162 936 165 1063
rect 178 1013 181 1096
rect 186 1093 197 1096
rect 194 1036 197 1093
rect 186 1033 197 1036
rect 154 933 165 936
rect 154 913 157 933
rect 178 916 181 1006
rect 170 913 181 916
rect 170 856 173 913
rect 170 853 181 856
rect 162 813 165 836
rect 178 826 181 853
rect 170 823 181 826
rect 170 806 173 823
rect 154 803 173 806
rect 154 696 157 796
rect 146 693 157 696
rect 130 613 133 646
rect 138 623 141 636
rect 146 616 149 693
rect 162 623 165 746
rect 138 613 149 616
rect 138 603 141 613
rect 114 403 117 506
rect 122 503 129 506
rect 138 503 141 596
rect 126 446 129 503
rect 162 446 165 616
rect 170 573 173 776
rect 178 653 181 816
rect 178 513 181 626
rect 186 486 189 1033
rect 194 603 197 1016
rect 218 1013 221 1106
rect 234 1096 237 1166
rect 242 1153 245 1436
rect 250 1413 253 1426
rect 250 1303 253 1406
rect 258 1333 261 1456
rect 250 1146 253 1296
rect 258 1243 261 1326
rect 258 1223 261 1236
rect 266 1223 269 1486
rect 274 1463 277 1493
rect 274 1396 277 1416
rect 282 1403 285 1486
rect 290 1453 293 1603
rect 290 1396 293 1416
rect 274 1393 293 1396
rect 258 1196 261 1216
rect 258 1193 265 1196
rect 230 1093 237 1096
rect 242 1143 253 1146
rect 202 916 205 946
rect 210 933 213 966
rect 230 936 233 1093
rect 242 946 245 1143
rect 250 1003 253 1126
rect 262 1036 265 1193
rect 258 1033 265 1036
rect 242 943 249 946
rect 230 933 237 936
rect 202 913 209 916
rect 206 836 209 913
rect 202 833 209 836
rect 202 786 205 833
rect 210 803 213 816
rect 202 783 209 786
rect 206 716 209 783
rect 206 713 213 716
rect 218 713 221 926
rect 226 823 229 916
rect 234 743 237 933
rect 246 896 249 943
rect 258 936 261 1033
rect 274 943 277 1386
rect 282 1313 285 1326
rect 282 1106 285 1246
rect 290 1183 293 1336
rect 298 1273 301 1596
rect 306 1483 309 1626
rect 314 1603 317 1713
rect 330 1626 333 1656
rect 338 1633 341 1646
rect 330 1623 341 1626
rect 322 1603 325 1616
rect 322 1556 325 1596
rect 314 1553 325 1556
rect 314 1473 317 1486
rect 306 1413 309 1456
rect 306 1283 309 1406
rect 314 1323 317 1436
rect 322 1393 325 1536
rect 330 1413 333 1616
rect 338 1566 341 1623
rect 346 1596 349 1676
rect 354 1653 357 1763
rect 370 1746 373 2166
rect 378 2023 381 2186
rect 378 1983 381 2016
rect 378 1923 381 1966
rect 386 1943 389 2136
rect 386 1826 389 1936
rect 378 1823 389 1826
rect 378 1763 381 1816
rect 362 1743 373 1746
rect 394 1746 397 2276
rect 402 1826 405 2283
rect 418 2226 421 2293
rect 410 2223 421 2226
rect 410 2203 413 2223
rect 418 2136 421 2206
rect 410 2003 413 2136
rect 418 2133 429 2136
rect 418 2103 421 2126
rect 426 2026 429 2133
rect 434 2123 437 2226
rect 458 2216 461 2236
rect 450 2213 461 2216
rect 450 2156 453 2213
rect 450 2153 461 2156
rect 434 2036 437 2066
rect 442 2046 445 2136
rect 458 2116 461 2153
rect 466 2123 469 2216
rect 450 2113 461 2116
rect 450 2103 453 2113
rect 442 2043 453 2046
rect 434 2033 445 2036
rect 418 2013 421 2026
rect 426 2023 445 2026
rect 426 1993 429 2006
rect 410 1846 413 1986
rect 418 1856 421 1966
rect 434 1953 437 2016
rect 442 1993 445 2023
rect 450 2006 453 2043
rect 458 2033 461 2106
rect 466 2013 469 2116
rect 474 2113 477 2216
rect 482 2203 485 2226
rect 498 2156 501 2226
rect 482 2153 501 2156
rect 482 2113 485 2153
rect 490 2123 501 2126
rect 506 2103 509 2323
rect 522 2313 525 2346
rect 530 2213 533 2336
rect 538 2283 541 2326
rect 554 2263 557 2356
rect 586 2346 589 2423
rect 562 2333 565 2346
rect 586 2343 597 2346
rect 602 2343 605 2416
rect 634 2413 637 2453
rect 698 2446 701 2466
rect 694 2443 701 2446
rect 706 2443 709 2526
rect 722 2486 725 2543
rect 730 2533 733 2556
rect 746 2553 757 2556
rect 746 2523 749 2553
rect 770 2536 773 2633
rect 786 2603 789 2616
rect 818 2576 821 2643
rect 834 2613 837 2736
rect 850 2716 853 2726
rect 866 2723 869 2736
rect 874 2716 877 2736
rect 882 2723 885 2743
rect 850 2713 877 2716
rect 906 2706 909 2813
rect 930 2803 933 2906
rect 938 2903 949 2906
rect 970 2903 973 2926
rect 986 2923 997 2926
rect 938 2803 941 2816
rect 946 2813 949 2903
rect 954 2803 957 2816
rect 938 2733 941 2756
rect 962 2753 965 2896
rect 994 2843 997 2923
rect 1002 2916 1005 2926
rect 1010 2923 1013 2946
rect 1034 2916 1037 3016
rect 1046 2966 1049 3023
rect 1002 2913 1037 2916
rect 1042 2963 1049 2966
rect 1002 2883 1005 2913
rect 1042 2906 1045 2963
rect 1042 2903 1053 2906
rect 970 2803 973 2826
rect 1042 2823 1045 2846
rect 978 2723 981 2796
rect 1026 2783 1029 2816
rect 1042 2793 1045 2806
rect 1042 2706 1045 2726
rect 874 2703 909 2706
rect 1034 2703 1045 2706
rect 874 2626 877 2703
rect 874 2623 881 2626
rect 762 2533 773 2536
rect 802 2533 805 2576
rect 810 2573 821 2576
rect 762 2486 765 2533
rect 722 2483 733 2486
rect 762 2483 773 2486
rect 730 2466 733 2483
rect 730 2463 737 2466
rect 770 2463 773 2483
rect 514 2193 517 2206
rect 514 2113 517 2136
rect 522 2123 525 2146
rect 530 2133 533 2176
rect 482 2013 485 2026
rect 490 2006 493 2016
rect 450 2003 493 2006
rect 426 1943 445 1946
rect 426 1923 429 1943
rect 434 1923 437 1936
rect 442 1933 445 1943
rect 450 1916 453 2003
rect 498 1966 501 2066
rect 538 2053 541 2216
rect 546 2123 549 2186
rect 474 1963 501 1966
rect 446 1913 453 1916
rect 418 1853 437 1856
rect 410 1843 429 1846
rect 402 1823 421 1826
rect 402 1786 405 1816
rect 402 1783 413 1786
rect 394 1743 401 1746
rect 346 1593 357 1596
rect 338 1563 349 1566
rect 338 1533 341 1556
rect 338 1463 341 1526
rect 338 1396 341 1456
rect 346 1433 349 1563
rect 354 1513 357 1593
rect 362 1546 365 1743
rect 370 1553 373 1736
rect 386 1643 389 1736
rect 398 1646 401 1743
rect 410 1733 413 1783
rect 394 1643 401 1646
rect 378 1613 381 1636
rect 386 1583 389 1636
rect 362 1543 373 1546
rect 334 1393 341 1396
rect 322 1333 325 1366
rect 334 1316 337 1393
rect 298 1213 301 1226
rect 314 1216 317 1316
rect 334 1313 341 1316
rect 338 1293 341 1313
rect 306 1213 317 1216
rect 290 1123 293 1136
rect 282 1103 289 1106
rect 298 1103 301 1136
rect 286 1036 289 1103
rect 282 1033 289 1036
rect 282 1013 285 1033
rect 306 1016 309 1186
rect 314 1113 317 1213
rect 322 1083 325 1216
rect 330 1066 333 1266
rect 338 1103 341 1226
rect 346 1203 349 1426
rect 354 1413 357 1426
rect 354 1313 357 1346
rect 354 1183 357 1226
rect 362 1143 365 1536
rect 370 1136 373 1543
rect 378 1506 381 1566
rect 386 1523 389 1576
rect 378 1503 385 1506
rect 382 1436 385 1503
rect 378 1433 385 1436
rect 378 1403 381 1433
rect 386 1403 389 1416
rect 394 1386 397 1643
rect 402 1593 405 1626
rect 410 1543 413 1726
rect 418 1716 421 1823
rect 426 1813 429 1843
rect 426 1723 429 1786
rect 434 1783 437 1853
rect 446 1846 449 1913
rect 446 1843 453 1846
rect 418 1713 429 1716
rect 418 1613 421 1656
rect 402 1503 405 1536
rect 418 1533 421 1596
rect 426 1573 429 1713
rect 434 1613 437 1706
rect 442 1703 445 1826
rect 450 1803 453 1843
rect 450 1613 453 1786
rect 458 1763 461 1956
rect 466 1783 469 1816
rect 434 1586 437 1606
rect 442 1593 445 1606
rect 458 1603 461 1726
rect 434 1583 447 1586
rect 444 1566 447 1583
rect 442 1563 447 1566
rect 442 1556 445 1563
rect 458 1556 461 1566
rect 434 1553 445 1556
rect 450 1553 461 1556
rect 410 1523 421 1526
rect 434 1523 437 1553
rect 442 1516 445 1546
rect 450 1543 453 1553
rect 450 1523 453 1536
rect 386 1383 397 1386
rect 386 1343 389 1383
rect 402 1376 405 1476
rect 434 1446 437 1516
rect 442 1513 453 1516
rect 394 1373 405 1376
rect 410 1443 437 1446
rect 378 1316 381 1326
rect 386 1323 389 1336
rect 394 1323 397 1373
rect 410 1366 413 1443
rect 418 1413 421 1436
rect 434 1423 437 1443
rect 402 1363 413 1366
rect 418 1366 421 1406
rect 426 1373 429 1406
rect 434 1366 437 1416
rect 442 1403 445 1506
rect 450 1453 453 1513
rect 450 1383 453 1406
rect 418 1363 437 1366
rect 402 1316 405 1363
rect 418 1333 421 1346
rect 458 1326 461 1546
rect 378 1313 385 1316
rect 382 1246 385 1313
rect 382 1243 389 1246
rect 354 1133 373 1136
rect 346 1113 349 1126
rect 322 1063 333 1066
rect 306 1013 313 1016
rect 258 933 293 936
rect 242 893 249 896
rect 202 613 205 706
rect 210 683 213 713
rect 226 643 229 736
rect 234 713 237 726
rect 242 706 245 893
rect 250 813 253 826
rect 258 816 261 916
rect 282 913 285 926
rect 266 833 269 846
rect 274 823 277 836
rect 258 813 265 816
rect 234 703 245 706
rect 250 703 253 806
rect 262 746 265 813
rect 258 743 265 746
rect 194 493 197 526
rect 210 516 213 616
rect 218 613 221 636
rect 226 533 229 626
rect 234 616 237 703
rect 234 613 245 616
rect 206 513 213 516
rect 218 513 221 526
rect 234 523 237 606
rect 242 583 245 613
rect 250 583 253 636
rect 186 483 197 486
rect 126 443 133 446
rect 130 426 133 443
rect 130 423 137 426
rect 154 423 157 446
rect 162 443 169 446
rect 114 213 117 336
rect 122 203 125 416
rect 134 336 137 423
rect 130 333 137 336
rect 130 306 133 333
rect 146 323 149 416
rect 166 386 169 443
rect 194 413 197 483
rect 206 426 209 513
rect 242 506 245 576
rect 258 533 261 743
rect 282 733 285 896
rect 266 706 269 726
rect 266 703 277 706
rect 274 646 277 703
rect 266 643 277 646
rect 266 613 269 643
rect 290 636 293 933
rect 298 876 301 1006
rect 310 946 313 1013
rect 306 943 313 946
rect 306 886 309 943
rect 306 883 317 886
rect 298 873 309 876
rect 298 813 301 866
rect 298 733 301 746
rect 306 676 309 873
rect 314 813 317 883
rect 322 863 325 1063
rect 314 733 317 786
rect 314 693 317 716
rect 306 673 317 676
rect 290 633 317 636
rect 282 613 285 626
rect 290 613 293 626
rect 306 606 309 626
rect 274 603 309 606
rect 238 503 245 506
rect 202 423 209 426
rect 178 396 181 406
rect 202 403 205 423
rect 218 396 221 416
rect 178 393 221 396
rect 166 383 173 386
rect 170 333 173 383
rect 162 316 165 326
rect 202 316 205 336
rect 138 313 165 316
rect 194 313 205 316
rect 130 303 173 306
rect 90 173 93 196
rect 130 183 133 296
rect 154 143 157 216
rect 170 123 173 303
rect 194 246 197 313
rect 194 243 205 246
rect 194 203 197 226
rect 202 123 205 243
rect 210 206 213 393
rect 218 223 221 376
rect 226 323 229 496
rect 238 386 241 503
rect 238 383 245 386
rect 242 366 245 383
rect 250 373 253 526
rect 258 403 261 426
rect 242 363 253 366
rect 250 333 253 363
rect 234 323 253 326
rect 250 303 253 316
rect 258 273 261 336
rect 234 233 237 246
rect 210 203 217 206
rect 226 203 229 216
rect 214 116 217 203
rect 234 143 253 146
rect 226 126 229 136
rect 234 133 237 143
rect 226 123 237 126
rect 242 116 245 136
rect 250 123 253 143
rect 258 133 261 226
rect 266 123 269 586
rect 274 513 285 516
rect 274 203 277 416
rect 282 406 285 446
rect 290 423 293 596
rect 314 543 317 633
rect 322 593 325 856
rect 330 676 333 996
rect 338 903 341 1066
rect 346 1023 349 1036
rect 346 993 349 1006
rect 354 996 357 1133
rect 378 1123 381 1226
rect 386 1213 389 1243
rect 386 1113 389 1176
rect 362 1003 365 1026
rect 354 993 365 996
rect 346 903 349 916
rect 354 856 357 926
rect 362 893 365 993
rect 370 913 373 1046
rect 378 993 381 1016
rect 378 923 381 956
rect 386 906 389 1086
rect 346 853 357 856
rect 338 823 341 836
rect 338 733 341 816
rect 338 713 341 726
rect 330 673 341 676
rect 330 586 333 666
rect 322 583 333 586
rect 314 513 317 536
rect 322 523 325 583
rect 330 533 333 556
rect 338 523 341 673
rect 346 506 349 853
rect 354 713 357 816
rect 370 813 373 906
rect 382 903 389 906
rect 362 626 365 806
rect 370 706 373 806
rect 382 746 385 903
rect 394 773 397 1316
rect 402 1313 413 1316
rect 402 1213 405 1226
rect 402 1183 405 1206
rect 410 1173 413 1313
rect 418 1203 421 1216
rect 402 1123 412 1126
rect 402 1033 405 1123
rect 402 933 405 946
rect 382 743 389 746
rect 378 713 381 726
rect 370 703 377 706
rect 374 636 377 703
rect 374 633 381 636
rect 354 623 365 626
rect 354 603 357 623
rect 362 553 365 616
rect 378 613 381 633
rect 354 533 357 546
rect 338 503 349 506
rect 298 423 301 436
rect 338 426 341 503
rect 306 406 309 426
rect 314 413 317 426
rect 338 423 349 426
rect 282 403 289 406
rect 286 266 289 403
rect 306 403 341 406
rect 282 263 289 266
rect 282 243 285 263
rect 282 163 285 216
rect 298 213 301 396
rect 306 373 309 403
rect 322 313 325 336
rect 330 313 333 326
rect 346 323 349 423
rect 354 393 357 526
rect 354 236 357 336
rect 362 323 365 426
rect 370 403 373 566
rect 378 356 381 536
rect 374 353 381 356
rect 374 266 377 353
rect 322 223 325 236
rect 346 233 357 236
rect 274 123 277 136
rect 314 133 317 216
rect 346 203 349 233
rect 362 213 365 266
rect 374 263 381 266
rect 386 263 389 743
rect 394 663 397 746
rect 402 706 405 826
rect 410 753 413 1116
rect 418 906 421 1146
rect 426 1123 429 1286
rect 426 1006 429 1106
rect 434 1063 437 1326
rect 450 1323 461 1326
rect 442 1203 445 1226
rect 450 1206 453 1323
rect 466 1253 469 1736
rect 474 1263 477 1963
rect 498 1923 501 1956
rect 506 1943 509 2006
rect 514 1906 517 1936
rect 506 1903 517 1906
rect 482 1763 485 1816
rect 482 1613 485 1756
rect 490 1723 493 1846
rect 506 1826 509 1903
rect 506 1823 513 1826
rect 498 1783 501 1806
rect 510 1756 513 1823
rect 510 1753 517 1756
rect 506 1723 509 1736
rect 482 1533 485 1606
rect 482 1503 485 1526
rect 490 1503 493 1716
rect 498 1663 501 1716
rect 514 1713 517 1753
rect 522 1696 525 1926
rect 530 1776 533 2046
rect 538 2003 541 2026
rect 538 1813 541 1936
rect 546 1863 549 2116
rect 554 1923 557 2256
rect 562 2206 565 2326
rect 570 2323 573 2336
rect 594 2323 597 2343
rect 650 2333 653 2406
rect 666 2403 669 2416
rect 694 2386 697 2443
rect 706 2393 709 2416
rect 734 2386 737 2463
rect 746 2413 749 2446
rect 778 2403 781 2526
rect 794 2513 797 2526
rect 802 2403 805 2416
rect 694 2383 701 2386
rect 570 2223 597 2226
rect 562 2203 569 2206
rect 566 2086 569 2203
rect 562 2083 569 2086
rect 562 2023 565 2083
rect 562 1983 565 2016
rect 570 2003 573 2066
rect 562 1906 565 1976
rect 570 1923 573 1996
rect 578 1963 581 2216
rect 594 2213 597 2223
rect 610 2213 613 2246
rect 586 2143 589 2206
rect 586 2043 589 2136
rect 594 2123 597 2196
rect 602 2113 605 2136
rect 610 2123 613 2206
rect 586 1936 589 2006
rect 578 1933 589 1936
rect 578 1916 581 1933
rect 558 1903 565 1906
rect 570 1913 581 1916
rect 558 1836 561 1903
rect 558 1833 565 1836
rect 530 1773 541 1776
rect 506 1693 525 1696
rect 506 1603 509 1693
rect 514 1596 517 1636
rect 522 1613 525 1626
rect 530 1603 533 1766
rect 498 1563 501 1596
rect 506 1593 517 1596
rect 538 1593 541 1773
rect 546 1763 549 1816
rect 562 1813 565 1833
rect 554 1753 557 1806
rect 498 1493 501 1516
rect 506 1503 509 1593
rect 546 1586 549 1746
rect 538 1583 549 1586
rect 514 1523 517 1556
rect 522 1516 525 1546
rect 518 1513 525 1516
rect 498 1483 509 1486
rect 450 1203 461 1206
rect 450 1196 453 1203
rect 442 1193 453 1196
rect 466 1196 469 1226
rect 466 1193 477 1196
rect 434 1013 437 1036
rect 442 1023 445 1193
rect 450 1096 453 1156
rect 458 1116 461 1146
rect 466 1133 469 1186
rect 474 1123 477 1193
rect 482 1143 485 1416
rect 498 1383 501 1416
rect 498 1343 501 1356
rect 506 1333 509 1483
rect 518 1446 521 1513
rect 514 1443 521 1446
rect 514 1413 517 1443
rect 522 1403 525 1426
rect 530 1413 533 1516
rect 538 1473 541 1583
rect 530 1396 533 1406
rect 514 1393 533 1396
rect 514 1326 517 1393
rect 538 1376 541 1466
rect 546 1453 549 1566
rect 554 1506 557 1736
rect 562 1723 565 1736
rect 570 1693 573 1913
rect 586 1896 589 1916
rect 582 1893 589 1896
rect 582 1786 585 1893
rect 594 1853 597 2106
rect 602 2013 605 2086
rect 610 1993 613 2106
rect 602 1923 605 1936
rect 610 1906 613 1936
rect 606 1903 613 1906
rect 606 1836 609 1903
rect 606 1833 613 1836
rect 582 1783 589 1786
rect 578 1666 581 1766
rect 570 1663 581 1666
rect 562 1556 565 1646
rect 570 1563 573 1663
rect 586 1646 589 1783
rect 594 1723 597 1816
rect 602 1803 605 1816
rect 610 1813 613 1833
rect 618 1813 621 2296
rect 626 2213 629 2226
rect 626 2093 629 2126
rect 626 2026 629 2066
rect 634 2033 637 2326
rect 674 2323 677 2336
rect 642 2296 645 2316
rect 642 2293 653 2296
rect 650 2226 653 2293
rect 690 2246 693 2326
rect 698 2323 701 2383
rect 730 2383 737 2386
rect 722 2333 725 2346
rect 730 2323 733 2383
rect 738 2323 741 2336
rect 762 2313 765 2336
rect 794 2333 797 2396
rect 810 2323 813 2573
rect 818 2533 821 2556
rect 866 2546 869 2616
rect 878 2546 881 2623
rect 898 2603 901 2616
rect 938 2613 941 2696
rect 1034 2656 1037 2703
rect 1034 2653 1045 2656
rect 978 2576 981 2616
rect 1002 2603 1005 2616
rect 1042 2613 1045 2653
rect 1050 2596 1053 2903
rect 1058 2893 1061 3006
rect 1074 3003 1077 3043
rect 1082 3013 1085 3046
rect 1090 3003 1093 3206
rect 1098 3173 1101 3226
rect 1130 3223 1141 3226
rect 1114 3203 1125 3206
rect 1130 3163 1133 3223
rect 1146 3216 1149 3226
rect 1210 3223 1229 3226
rect 1138 3213 1149 3216
rect 1138 3183 1141 3213
rect 1146 3146 1149 3176
rect 1130 3143 1149 3146
rect 1098 3013 1101 3036
rect 1106 2973 1109 3136
rect 1114 3103 1117 3126
rect 1114 2966 1117 3016
rect 1122 2976 1125 3136
rect 1130 3106 1133 3143
rect 1138 3123 1141 3136
rect 1146 3133 1149 3143
rect 1154 3126 1157 3156
rect 1146 3123 1157 3126
rect 1162 3116 1165 3126
rect 1138 3113 1165 3116
rect 1170 3116 1173 3146
rect 1170 3113 1177 3116
rect 1186 3113 1189 3206
rect 1202 3193 1205 3216
rect 1210 3143 1213 3223
rect 1218 3213 1229 3216
rect 1234 3213 1237 3276
rect 1242 3156 1245 3236
rect 1250 3223 1253 3236
rect 1234 3133 1237 3156
rect 1242 3153 1285 3156
rect 1250 3133 1253 3146
rect 1266 3133 1269 3146
rect 1130 3103 1149 3106
rect 1130 3023 1133 3046
rect 1130 2993 1133 3006
rect 1138 2983 1141 3016
rect 1146 3003 1149 3103
rect 1162 3076 1165 3096
rect 1158 3073 1165 3076
rect 1158 3016 1161 3073
rect 1174 3066 1177 3113
rect 1218 3093 1221 3126
rect 1226 3083 1229 3126
rect 1170 3063 1177 3066
rect 1158 3013 1165 3016
rect 1162 2996 1165 3013
rect 1170 3006 1173 3063
rect 1186 3023 1237 3026
rect 1186 3013 1189 3023
rect 1170 3003 1197 3006
rect 1162 2993 1181 2996
rect 1202 2993 1205 3016
rect 1218 3013 1237 3016
rect 1122 2973 1133 2976
rect 1114 2963 1125 2966
rect 1122 2943 1125 2963
rect 1106 2923 1109 2936
rect 1130 2926 1133 2973
rect 1154 2946 1157 2966
rect 1154 2943 1161 2946
rect 1126 2923 1133 2926
rect 1058 2803 1061 2886
rect 1058 2723 1061 2786
rect 1066 2743 1069 2876
rect 1126 2866 1129 2923
rect 1138 2883 1141 2926
rect 1146 2873 1149 2926
rect 1158 2866 1161 2943
rect 1170 2906 1173 2936
rect 1178 2926 1181 2993
rect 1210 2973 1213 3006
rect 1234 2966 1237 3006
rect 1210 2963 1237 2966
rect 1186 2933 1197 2936
rect 1210 2933 1213 2963
rect 1178 2923 1197 2926
rect 1218 2916 1221 2926
rect 1234 2923 1237 2956
rect 1242 2926 1245 3126
rect 1266 3123 1277 3126
rect 1282 3116 1285 3153
rect 1274 3113 1285 3116
rect 1290 3113 1293 3216
rect 1306 3213 1309 3246
rect 1298 3193 1301 3206
rect 1314 3203 1317 3216
rect 1322 3206 1325 3276
rect 1330 3233 1349 3236
rect 1330 3213 1333 3233
rect 1322 3203 1333 3206
rect 1330 3156 1333 3203
rect 1338 3183 1341 3216
rect 1346 3213 1349 3233
rect 1354 3223 1357 3246
rect 1362 3203 1365 3266
rect 1418 3213 1421 3236
rect 1498 3223 1501 3236
rect 1578 3233 1605 3236
rect 1538 3223 1549 3226
rect 1402 3163 1405 3206
rect 1418 3156 1421 3206
rect 1426 3173 1429 3216
rect 1482 3213 1501 3216
rect 1538 3213 1549 3216
rect 1578 3213 1581 3233
rect 1634 3216 1637 3266
rect 1642 3233 1685 3236
rect 1642 3223 1645 3233
rect 1474 3186 1477 3206
rect 1490 3193 1493 3213
rect 1538 3206 1541 3213
rect 1474 3183 1509 3186
rect 1298 3153 1333 3156
rect 1298 3123 1301 3153
rect 1314 3133 1317 3146
rect 1330 3133 1333 3153
rect 1378 3153 1421 3156
rect 1258 2986 1261 3016
rect 1266 2996 1269 3056
rect 1274 3003 1277 3113
rect 1306 3083 1309 3126
rect 1282 3013 1285 3026
rect 1290 3013 1293 3066
rect 1322 3036 1325 3126
rect 1330 3123 1365 3126
rect 1370 3123 1373 3136
rect 1362 3106 1365 3123
rect 1318 3033 1325 3036
rect 1354 3103 1365 3106
rect 1354 3036 1357 3103
rect 1354 3033 1365 3036
rect 1282 2996 1285 3006
rect 1266 2993 1285 2996
rect 1250 2933 1253 2986
rect 1258 2983 1269 2986
rect 1258 2933 1261 2946
rect 1242 2923 1253 2926
rect 1266 2923 1269 2983
rect 1306 2943 1309 3026
rect 1194 2913 1221 2916
rect 1170 2903 1213 2906
rect 1082 2743 1085 2786
rect 1066 2693 1069 2736
rect 1090 2723 1093 2866
rect 1126 2863 1133 2866
rect 1130 2846 1133 2863
rect 1154 2863 1161 2866
rect 1130 2843 1141 2846
rect 1114 2763 1117 2806
rect 1138 2743 1141 2843
rect 1154 2826 1157 2863
rect 1150 2823 1157 2826
rect 1150 2756 1153 2823
rect 1162 2793 1165 2816
rect 1150 2753 1157 2756
rect 1114 2723 1117 2736
rect 922 2573 981 2576
rect 1042 2593 1053 2596
rect 858 2543 869 2546
rect 874 2543 881 2546
rect 858 2533 861 2543
rect 858 2413 861 2526
rect 866 2503 869 2536
rect 874 2493 877 2543
rect 914 2533 917 2556
rect 922 2523 925 2573
rect 1042 2546 1045 2593
rect 1042 2543 1053 2546
rect 938 2523 941 2536
rect 954 2446 957 2466
rect 954 2443 961 2446
rect 826 2333 829 2346
rect 850 2323 853 2366
rect 698 2253 701 2296
rect 690 2243 701 2246
rect 642 2223 653 2226
rect 642 2163 645 2223
rect 626 2023 637 2026
rect 626 2003 629 2016
rect 594 1653 597 1716
rect 586 1643 597 1646
rect 562 1553 573 1556
rect 570 1523 573 1553
rect 578 1543 581 1626
rect 586 1603 589 1616
rect 586 1536 589 1596
rect 594 1543 597 1643
rect 578 1533 589 1536
rect 554 1503 565 1506
rect 562 1436 565 1503
rect 498 1323 517 1326
rect 522 1373 541 1376
rect 458 1113 477 1116
rect 450 1093 461 1096
rect 458 1036 461 1093
rect 450 1033 461 1036
rect 442 1006 445 1016
rect 450 1013 453 1033
rect 466 1006 469 1016
rect 426 1003 445 1006
rect 450 1003 469 1006
rect 426 913 429 976
rect 418 903 429 906
rect 418 813 421 836
rect 418 743 421 806
rect 426 773 429 903
rect 434 803 437 996
rect 450 993 469 996
rect 450 943 453 993
rect 474 946 477 1113
rect 466 943 477 946
rect 466 926 469 943
rect 462 923 469 926
rect 442 913 453 916
rect 442 766 445 836
rect 450 813 453 913
rect 462 856 465 923
rect 462 853 469 856
rect 466 813 469 853
rect 474 806 477 926
rect 482 816 485 1136
rect 490 1093 493 1126
rect 498 1106 501 1323
rect 522 1306 525 1373
rect 514 1303 525 1306
rect 514 1246 517 1303
rect 514 1243 525 1246
rect 514 1213 517 1226
rect 506 1123 509 1206
rect 498 1103 505 1106
rect 490 1003 493 1066
rect 502 1016 505 1103
rect 498 1013 505 1016
rect 498 996 501 1013
rect 490 993 501 996
rect 490 833 493 993
rect 514 956 517 1136
rect 522 973 525 1243
rect 530 1033 533 1346
rect 538 1026 541 1336
rect 546 1046 549 1436
rect 554 1433 565 1436
rect 578 1433 581 1533
rect 554 1186 557 1433
rect 562 1413 573 1416
rect 562 1383 565 1406
rect 578 1366 581 1426
rect 586 1416 589 1526
rect 594 1463 597 1536
rect 586 1413 597 1416
rect 562 1363 581 1366
rect 562 1323 565 1363
rect 562 1203 565 1246
rect 554 1183 561 1186
rect 558 1076 561 1183
rect 554 1073 561 1076
rect 554 1053 557 1073
rect 546 1043 557 1046
rect 530 1023 541 1026
rect 498 953 517 956
rect 482 813 489 816
rect 426 763 445 766
rect 458 803 477 806
rect 410 723 421 726
rect 426 723 429 763
rect 458 756 461 803
rect 434 753 461 756
rect 402 703 409 706
rect 406 656 409 703
rect 402 653 409 656
rect 394 523 397 606
rect 402 543 405 653
rect 410 533 413 616
rect 394 423 397 436
rect 402 416 405 526
rect 418 473 421 686
rect 426 526 429 716
rect 434 613 437 753
rect 458 743 469 746
rect 458 736 461 743
rect 442 733 461 736
rect 442 716 445 733
rect 442 713 449 716
rect 446 636 449 713
rect 458 693 461 716
rect 442 633 449 636
rect 442 613 445 633
rect 450 566 453 616
rect 458 603 461 626
rect 466 613 469 726
rect 474 613 477 756
rect 486 746 489 813
rect 482 743 489 746
rect 482 606 485 743
rect 498 726 501 953
rect 506 833 509 936
rect 514 923 517 946
rect 506 813 509 826
rect 514 796 517 916
rect 522 806 525 936
rect 530 913 533 1023
rect 538 1013 549 1016
rect 538 816 541 1006
rect 546 983 549 1013
rect 546 823 549 976
rect 530 813 541 816
rect 522 803 541 806
rect 506 756 509 796
rect 514 793 533 796
rect 506 753 517 756
rect 490 723 501 726
rect 506 723 509 736
rect 490 703 493 723
rect 514 716 517 753
rect 498 713 517 716
rect 522 713 525 766
rect 466 603 485 606
rect 490 603 493 676
rect 442 563 453 566
rect 442 533 445 563
rect 466 533 469 603
rect 498 573 501 713
rect 506 696 509 706
rect 514 703 525 706
rect 506 693 517 696
rect 506 613 509 626
rect 474 543 509 546
rect 426 523 445 526
rect 474 523 477 543
rect 514 536 517 693
rect 522 583 525 703
rect 530 653 533 793
rect 538 723 541 803
rect 546 613 549 816
rect 554 706 557 1043
rect 562 953 565 1006
rect 562 913 565 946
rect 562 793 565 906
rect 570 753 573 1336
rect 578 1303 581 1336
rect 586 1323 589 1406
rect 594 1343 597 1413
rect 594 1323 597 1336
rect 594 1233 597 1286
rect 578 1213 581 1226
rect 586 1203 589 1216
rect 578 1043 581 1146
rect 586 1123 589 1176
rect 594 1133 597 1146
rect 594 1093 597 1126
rect 602 1086 605 1786
rect 610 1736 613 1806
rect 626 1763 629 1916
rect 634 1823 637 2023
rect 642 1903 645 2156
rect 650 2113 653 2206
rect 666 2193 669 2206
rect 674 2153 677 2206
rect 658 2133 669 2136
rect 682 2133 685 2146
rect 690 2133 693 2226
rect 650 1926 653 2026
rect 658 1993 661 2066
rect 666 2013 669 2126
rect 658 1933 661 1946
rect 650 1923 661 1926
rect 650 1903 653 1916
rect 658 1886 661 1923
rect 650 1883 661 1886
rect 610 1733 621 1736
rect 610 1683 613 1726
rect 610 1613 613 1666
rect 610 1333 613 1556
rect 618 1326 621 1733
rect 626 1713 629 1756
rect 634 1733 637 1816
rect 626 1633 629 1706
rect 626 1563 629 1616
rect 634 1556 637 1726
rect 642 1703 645 1816
rect 650 1723 653 1883
rect 666 1823 669 2006
rect 674 1996 677 2036
rect 682 2003 685 2026
rect 674 1993 685 1996
rect 682 1923 685 1993
rect 690 1916 693 2126
rect 698 2103 701 2243
rect 682 1913 693 1916
rect 682 1846 685 1913
rect 674 1843 685 1846
rect 674 1816 677 1843
rect 698 1826 701 2096
rect 706 1923 709 2306
rect 818 2303 821 2316
rect 714 2213 717 2256
rect 738 2213 741 2236
rect 746 2213 757 2216
rect 762 2213 765 2286
rect 850 2246 853 2316
rect 850 2243 861 2246
rect 802 2223 805 2236
rect 722 2126 725 2206
rect 722 2123 733 2126
rect 738 2123 741 2146
rect 746 2123 749 2166
rect 754 2133 757 2213
rect 778 2193 781 2206
rect 786 2186 789 2206
rect 802 2203 805 2216
rect 786 2183 797 2186
rect 714 1963 717 2116
rect 730 2036 733 2123
rect 778 2116 781 2146
rect 794 2126 797 2183
rect 810 2173 813 2206
rect 794 2123 813 2126
rect 762 2113 781 2116
rect 786 2113 805 2116
rect 722 2033 733 2036
rect 722 2013 725 2033
rect 730 1966 733 2006
rect 746 1983 749 1996
rect 746 1966 749 1976
rect 730 1963 749 1966
rect 714 1876 717 1936
rect 738 1926 741 1936
rect 730 1923 741 1926
rect 730 1906 733 1923
rect 730 1903 737 1906
rect 714 1873 725 1876
rect 658 1813 677 1816
rect 682 1823 709 1826
rect 658 1743 661 1813
rect 682 1806 685 1823
rect 690 1813 701 1816
rect 706 1813 709 1823
rect 714 1806 717 1866
rect 674 1803 685 1806
rect 666 1733 669 1746
rect 674 1693 677 1803
rect 698 1786 701 1806
rect 694 1783 701 1786
rect 706 1803 717 1806
rect 682 1656 685 1736
rect 650 1653 685 1656
rect 642 1603 645 1636
rect 650 1603 653 1653
rect 658 1576 661 1646
rect 666 1623 677 1626
rect 674 1593 677 1606
rect 682 1603 685 1653
rect 694 1646 697 1783
rect 706 1726 709 1803
rect 722 1726 725 1873
rect 734 1826 737 1903
rect 730 1823 737 1826
rect 730 1803 733 1823
rect 738 1733 741 1796
rect 706 1723 717 1726
rect 722 1723 733 1726
rect 746 1723 749 1963
rect 754 1903 757 2046
rect 762 1913 765 2113
rect 778 2043 797 2046
rect 770 1993 773 2016
rect 778 2013 781 2043
rect 794 2013 797 2026
rect 786 1986 789 2006
rect 782 1983 789 1986
rect 782 1936 785 1983
rect 794 1943 797 1956
rect 782 1933 789 1936
rect 786 1856 789 1933
rect 794 1856 797 1886
rect 802 1863 805 2113
rect 810 1983 813 2123
rect 818 2013 821 2196
rect 818 1973 821 2006
rect 826 2003 829 2146
rect 834 1996 837 2146
rect 842 2123 845 2216
rect 850 2173 853 2243
rect 858 2203 861 2226
rect 866 2146 869 2216
rect 858 2143 869 2146
rect 850 2033 853 2136
rect 858 2083 861 2143
rect 866 2113 869 2136
rect 842 2023 853 2026
rect 842 2013 853 2016
rect 826 1993 837 1996
rect 786 1853 805 1856
rect 770 1813 773 1826
rect 802 1823 805 1853
rect 810 1813 813 1926
rect 818 1913 821 1926
rect 826 1906 829 1993
rect 834 1923 837 1976
rect 818 1903 829 1906
rect 818 1866 821 1903
rect 826 1886 829 1896
rect 842 1893 845 1906
rect 850 1903 853 1916
rect 858 1903 861 2026
rect 866 1973 869 2106
rect 866 1933 869 1956
rect 874 1926 877 2436
rect 890 2403 893 2416
rect 938 2393 941 2416
rect 958 2376 961 2443
rect 970 2413 973 2516
rect 978 2486 981 2526
rect 1026 2503 1029 2536
rect 978 2483 1021 2486
rect 1010 2413 1013 2466
rect 1018 2416 1021 2483
rect 1050 2436 1053 2543
rect 1058 2533 1061 2556
rect 1082 2523 1085 2616
rect 1098 2586 1101 2606
rect 1114 2586 1117 2656
rect 1138 2613 1141 2736
rect 1146 2723 1149 2736
rect 1154 2706 1157 2753
rect 1150 2703 1157 2706
rect 1098 2583 1117 2586
rect 1150 2586 1153 2703
rect 1150 2583 1157 2586
rect 1154 2563 1157 2583
rect 1162 2566 1165 2746
rect 1170 2716 1173 2746
rect 1186 2723 1189 2746
rect 1194 2733 1197 2816
rect 1202 2726 1205 2816
rect 1210 2803 1213 2903
rect 1250 2823 1253 2923
rect 1290 2896 1293 2936
rect 1318 2896 1321 3033
rect 1330 2903 1333 3026
rect 1338 2963 1341 3006
rect 1346 2983 1349 3016
rect 1354 3003 1357 3016
rect 1362 2953 1365 3033
rect 1370 2973 1373 3016
rect 1378 3003 1381 3153
rect 1402 3133 1405 3146
rect 1410 3133 1413 3153
rect 1434 3133 1437 3156
rect 1402 3113 1405 3126
rect 1410 3073 1413 3126
rect 1474 3113 1477 3136
rect 1418 3013 1421 3026
rect 1426 3023 1437 3026
rect 1338 2923 1341 2946
rect 1282 2893 1293 2896
rect 1306 2893 1321 2896
rect 1282 2836 1285 2893
rect 1282 2833 1293 2836
rect 1250 2793 1253 2806
rect 1258 2776 1261 2816
rect 1266 2803 1269 2816
rect 1290 2786 1293 2833
rect 1306 2823 1309 2893
rect 1330 2816 1333 2886
rect 1370 2883 1373 2926
rect 1378 2856 1381 2926
rect 1386 2913 1389 2936
rect 1314 2813 1333 2816
rect 1354 2853 1381 2856
rect 1354 2813 1357 2853
rect 1394 2813 1397 2936
rect 1410 2926 1413 2976
rect 1418 2963 1421 3006
rect 1418 2933 1421 2946
rect 1402 2906 1405 2926
rect 1410 2923 1421 2926
rect 1402 2903 1409 2906
rect 1306 2796 1309 2806
rect 1314 2803 1317 2813
rect 1406 2806 1409 2903
rect 1306 2793 1341 2796
rect 1290 2783 1317 2786
rect 1234 2773 1277 2776
rect 1234 2743 1237 2773
rect 1242 2743 1253 2746
rect 1194 2723 1205 2726
rect 1194 2716 1197 2723
rect 1170 2713 1197 2716
rect 1242 2716 1245 2736
rect 1250 2726 1253 2743
rect 1258 2733 1261 2746
rect 1250 2723 1261 2726
rect 1274 2723 1277 2773
rect 1290 2763 1293 2783
rect 1314 2733 1317 2783
rect 1338 2723 1341 2793
rect 1370 2763 1373 2806
rect 1402 2803 1409 2806
rect 1394 2723 1397 2746
rect 1402 2743 1405 2803
rect 1242 2713 1253 2716
rect 1258 2713 1261 2723
rect 1402 2716 1405 2736
rect 1378 2713 1405 2716
rect 1210 2576 1213 2616
rect 1226 2603 1229 2616
rect 1250 2613 1253 2713
rect 1162 2563 1173 2566
rect 1098 2523 1101 2536
rect 1050 2433 1061 2436
rect 1018 2413 1029 2416
rect 954 2373 961 2376
rect 890 2343 933 2346
rect 890 2316 893 2343
rect 886 2313 893 2316
rect 886 2236 889 2313
rect 886 2233 893 2236
rect 882 1946 885 2216
rect 890 2203 893 2233
rect 898 2213 901 2336
rect 922 2326 925 2336
rect 930 2333 933 2343
rect 914 2323 925 2326
rect 906 2196 909 2266
rect 914 2223 917 2323
rect 922 2263 925 2316
rect 902 2193 909 2196
rect 890 2103 893 2176
rect 902 2136 905 2193
rect 914 2143 917 2216
rect 922 2143 925 2206
rect 938 2193 941 2326
rect 954 2306 957 2373
rect 978 2323 981 2406
rect 1026 2403 1029 2413
rect 954 2303 965 2306
rect 962 2236 965 2303
rect 954 2233 965 2236
rect 946 2156 949 2216
rect 938 2153 949 2156
rect 954 2156 957 2233
rect 986 2226 989 2336
rect 986 2223 993 2226
rect 954 2153 965 2156
rect 938 2136 941 2153
rect 946 2143 957 2146
rect 902 2133 909 2136
rect 890 1956 893 2096
rect 898 1973 901 2006
rect 906 1996 909 2133
rect 914 2006 917 2046
rect 922 2016 925 2136
rect 930 2063 933 2136
rect 938 2133 949 2136
rect 938 2083 941 2126
rect 922 2013 933 2016
rect 938 2013 941 2046
rect 914 2003 925 2006
rect 906 1993 941 1996
rect 890 1953 925 1956
rect 882 1943 893 1946
rect 826 1883 845 1886
rect 818 1863 825 1866
rect 754 1733 757 1806
rect 762 1803 789 1806
rect 706 1663 709 1716
rect 694 1643 701 1646
rect 698 1626 701 1643
rect 698 1623 709 1626
rect 626 1553 637 1556
rect 642 1573 661 1576
rect 626 1336 629 1553
rect 634 1533 637 1546
rect 642 1473 645 1573
rect 650 1456 653 1546
rect 634 1453 653 1456
rect 634 1413 637 1453
rect 642 1433 645 1446
rect 634 1366 637 1406
rect 642 1373 645 1426
rect 650 1393 653 1416
rect 634 1363 645 1366
rect 626 1333 637 1336
rect 610 1243 613 1326
rect 618 1323 629 1326
rect 610 1183 613 1226
rect 618 1143 621 1296
rect 626 1153 629 1323
rect 634 1263 637 1333
rect 642 1323 645 1363
rect 650 1333 653 1346
rect 642 1203 645 1226
rect 650 1223 653 1236
rect 650 1146 653 1216
rect 626 1143 653 1146
rect 594 1083 605 1086
rect 610 1133 621 1136
rect 578 973 581 1036
rect 594 936 597 1083
rect 610 1013 613 1133
rect 626 1126 629 1143
rect 618 1123 629 1126
rect 618 1023 621 1123
rect 642 1113 645 1126
rect 658 1076 661 1566
rect 690 1556 693 1616
rect 714 1603 717 1723
rect 722 1586 725 1716
rect 718 1583 725 1586
rect 690 1553 709 1556
rect 666 1503 669 1526
rect 666 1383 669 1426
rect 666 1293 669 1356
rect 674 1333 677 1536
rect 690 1526 693 1536
rect 698 1533 701 1546
rect 706 1533 709 1553
rect 718 1526 721 1583
rect 682 1523 693 1526
rect 698 1523 721 1526
rect 682 1313 685 1476
rect 690 1353 693 1416
rect 690 1236 693 1336
rect 698 1246 701 1523
rect 706 1503 709 1516
rect 714 1426 717 1506
rect 730 1473 733 1723
rect 738 1703 741 1716
rect 754 1696 757 1726
rect 738 1693 757 1696
rect 738 1523 741 1693
rect 714 1423 721 1426
rect 706 1403 709 1416
rect 706 1313 709 1396
rect 718 1346 721 1423
rect 730 1416 733 1456
rect 746 1443 749 1686
rect 762 1596 765 1803
rect 794 1746 797 1766
rect 770 1733 773 1746
rect 794 1743 801 1746
rect 786 1706 789 1736
rect 778 1703 789 1706
rect 770 1613 773 1626
rect 778 1613 781 1703
rect 798 1676 801 1743
rect 798 1673 805 1676
rect 758 1593 765 1596
rect 758 1526 761 1593
rect 754 1523 761 1526
rect 770 1523 773 1576
rect 754 1503 757 1523
rect 770 1503 773 1516
rect 738 1423 741 1436
rect 730 1413 741 1416
rect 746 1413 749 1436
rect 754 1423 765 1426
rect 770 1423 773 1436
rect 754 1413 765 1416
rect 738 1403 741 1413
rect 714 1343 721 1346
rect 738 1346 741 1376
rect 738 1343 749 1346
rect 698 1243 709 1246
rect 690 1233 701 1236
rect 666 1213 669 1226
rect 690 1213 693 1226
rect 666 1203 677 1206
rect 666 1093 669 1203
rect 658 1073 665 1076
rect 650 1036 653 1056
rect 586 933 597 936
rect 578 843 581 926
rect 586 903 589 933
rect 594 903 597 916
rect 626 913 629 1006
rect 634 903 637 1036
rect 646 1033 653 1036
rect 646 876 649 1033
rect 662 1026 665 1073
rect 674 1033 677 1146
rect 690 1123 693 1206
rect 698 1116 701 1233
rect 706 1163 709 1243
rect 690 1113 701 1116
rect 706 1113 709 1126
rect 658 1023 665 1026
rect 646 873 653 876
rect 578 813 581 836
rect 610 803 613 836
rect 618 783 621 816
rect 626 813 629 866
rect 642 833 645 856
rect 562 716 565 736
rect 578 733 605 736
rect 570 723 581 726
rect 562 713 581 716
rect 554 703 565 706
rect 482 533 517 536
rect 482 523 485 533
rect 442 503 445 523
rect 506 506 509 526
rect 514 523 517 533
rect 522 506 525 576
rect 498 503 509 506
rect 518 503 525 506
rect 442 423 469 426
rect 398 413 405 416
rect 398 346 401 413
rect 410 363 413 406
rect 418 396 421 416
rect 426 413 437 416
rect 442 413 445 423
rect 450 396 453 406
rect 418 393 453 396
rect 394 343 401 346
rect 394 293 397 343
rect 410 323 413 336
rect 418 333 421 393
rect 426 323 429 356
rect 378 243 381 263
rect 370 233 389 236
rect 214 113 245 116
rect 330 113 333 136
rect 338 123 341 136
rect 346 133 349 166
rect 378 163 381 226
rect 394 223 397 246
rect 434 223 437 336
rect 442 293 445 336
rect 458 323 461 416
rect 474 346 477 476
rect 498 456 501 503
rect 498 453 509 456
rect 506 433 509 453
rect 518 426 521 503
rect 506 423 521 426
rect 466 343 477 346
rect 354 123 357 156
rect 402 133 405 166
rect 410 123 413 216
rect 418 203 421 216
rect 426 213 445 216
rect 418 113 421 136
rect 426 113 429 213
rect 434 203 445 206
rect 466 203 469 343
rect 498 333 501 366
rect 490 323 501 326
rect 506 323 509 423
rect 530 416 533 606
rect 546 603 557 606
rect 562 596 565 703
rect 538 593 565 596
rect 538 423 541 593
rect 562 543 565 556
rect 546 533 565 536
rect 514 383 517 416
rect 530 413 541 416
rect 538 403 541 413
rect 546 393 549 496
rect 562 483 565 533
rect 578 523 581 713
rect 594 696 597 726
rect 586 693 597 696
rect 594 603 597 686
rect 562 386 565 466
rect 586 426 589 586
rect 602 493 605 733
rect 610 716 613 776
rect 626 746 629 806
rect 634 773 637 826
rect 618 743 637 746
rect 618 733 621 743
rect 610 713 617 716
rect 626 713 629 736
rect 634 716 637 743
rect 642 723 645 736
rect 634 713 645 716
rect 614 636 617 713
rect 610 633 617 636
rect 610 613 613 633
rect 634 616 637 626
rect 618 613 637 616
rect 634 583 637 606
rect 626 533 629 556
rect 626 493 629 526
rect 634 523 637 536
rect 642 506 645 626
rect 650 606 653 873
rect 658 683 661 1023
rect 666 933 669 956
rect 674 903 677 1026
rect 690 1016 693 1056
rect 682 1013 693 1016
rect 666 816 669 836
rect 674 823 677 866
rect 666 813 677 816
rect 666 633 669 776
rect 674 743 677 813
rect 682 736 685 986
rect 698 946 701 1026
rect 690 943 701 946
rect 690 913 693 926
rect 714 916 717 1343
rect 722 1313 725 1326
rect 730 1293 733 1326
rect 746 1313 749 1343
rect 754 1333 757 1406
rect 754 1306 757 1326
rect 762 1323 765 1413
rect 778 1406 781 1606
rect 794 1586 797 1666
rect 802 1603 805 1673
rect 810 1613 813 1796
rect 822 1746 825 1863
rect 818 1743 825 1746
rect 834 1743 837 1806
rect 794 1583 801 1586
rect 786 1533 789 1576
rect 786 1433 789 1526
rect 798 1486 801 1583
rect 810 1563 813 1596
rect 810 1513 813 1556
rect 794 1483 801 1486
rect 794 1426 797 1483
rect 774 1403 781 1406
rect 786 1423 797 1426
rect 774 1316 777 1403
rect 738 1303 757 1306
rect 762 1296 765 1316
rect 774 1313 781 1316
rect 722 1093 725 1216
rect 730 1013 733 1276
rect 698 883 701 916
rect 706 913 717 916
rect 722 913 725 926
rect 730 913 733 926
rect 706 896 709 913
rect 714 903 725 906
rect 706 893 717 896
rect 690 823 693 846
rect 698 743 709 746
rect 674 733 685 736
rect 674 613 677 733
rect 650 603 677 606
rect 638 503 645 506
rect 638 436 641 503
rect 650 446 653 546
rect 658 463 661 586
rect 666 513 669 526
rect 650 443 669 446
rect 618 433 629 436
rect 638 433 645 436
rect 586 423 597 426
rect 538 383 565 386
rect 570 386 573 406
rect 578 403 581 416
rect 570 383 577 386
rect 522 333 525 376
rect 538 316 541 383
rect 562 346 565 366
rect 514 313 541 316
rect 554 343 565 346
rect 514 223 517 313
rect 530 223 533 236
rect 554 226 557 343
rect 574 336 577 383
rect 594 366 597 423
rect 618 413 621 433
rect 626 403 629 426
rect 570 333 577 336
rect 586 363 597 366
rect 490 93 493 126
rect 498 123 501 186
rect 514 183 517 206
rect 506 116 509 136
rect 514 123 517 166
rect 522 133 525 216
rect 538 213 541 226
rect 554 223 565 226
rect 562 133 565 223
rect 570 206 573 333
rect 578 223 581 256
rect 586 216 589 363
rect 634 346 637 416
rect 642 403 645 433
rect 594 343 637 346
rect 594 333 597 343
rect 610 313 613 326
rect 586 213 597 216
rect 618 213 621 336
rect 642 333 645 346
rect 650 323 653 406
rect 658 393 661 416
rect 658 316 661 336
rect 642 303 645 316
rect 650 313 661 316
rect 650 213 653 313
rect 570 203 577 206
rect 574 126 577 203
rect 594 136 597 213
rect 666 203 669 443
rect 674 376 677 603
rect 682 533 685 726
rect 690 723 693 736
rect 714 733 717 893
rect 738 886 741 1166
rect 746 1116 749 1266
rect 754 1223 757 1296
rect 762 1293 769 1296
rect 766 1226 769 1293
rect 762 1223 769 1226
rect 762 1203 765 1223
rect 778 1206 781 1313
rect 786 1286 789 1423
rect 794 1403 797 1416
rect 802 1396 805 1416
rect 810 1403 813 1426
rect 802 1393 813 1396
rect 794 1303 797 1316
rect 786 1283 793 1286
rect 774 1203 781 1206
rect 774 1146 777 1203
rect 790 1196 793 1283
rect 754 1133 757 1146
rect 762 1143 777 1146
rect 786 1193 793 1196
rect 746 1113 753 1116
rect 750 1026 753 1113
rect 730 883 741 886
rect 746 1023 753 1026
rect 730 816 733 883
rect 730 813 741 816
rect 738 793 741 813
rect 722 723 725 736
rect 730 706 733 726
rect 722 703 733 706
rect 690 613 693 626
rect 698 616 701 636
rect 722 616 725 703
rect 738 693 741 736
rect 698 613 705 616
rect 690 583 693 606
rect 690 513 693 576
rect 702 546 705 613
rect 698 543 705 546
rect 714 613 725 616
rect 698 506 701 543
rect 682 503 701 506
rect 682 393 685 503
rect 706 486 709 526
rect 690 483 709 486
rect 674 373 681 376
rect 690 373 693 483
rect 714 476 717 613
rect 730 593 733 606
rect 698 473 717 476
rect 678 316 681 373
rect 698 333 701 473
rect 706 386 709 416
rect 722 413 725 466
rect 714 403 725 406
rect 730 403 733 516
rect 738 443 741 686
rect 722 396 725 403
rect 738 396 741 406
rect 722 393 741 396
rect 706 383 733 386
rect 714 333 725 336
rect 678 313 685 316
rect 682 246 685 313
rect 714 306 717 333
rect 722 316 725 326
rect 730 323 733 383
rect 746 363 749 1023
rect 754 933 757 1006
rect 754 803 757 846
rect 762 803 765 1143
rect 770 1133 781 1136
rect 770 1023 773 1086
rect 770 946 773 1006
rect 778 993 781 1006
rect 770 943 781 946
rect 770 883 773 943
rect 754 736 757 746
rect 770 736 773 816
rect 778 746 781 816
rect 786 803 789 1193
rect 794 1133 797 1166
rect 794 1093 797 1126
rect 802 1076 805 1386
rect 810 1303 813 1393
rect 818 1296 821 1743
rect 842 1733 845 1883
rect 850 1773 853 1816
rect 810 1293 821 1296
rect 810 1193 813 1293
rect 818 1223 821 1276
rect 798 1073 805 1076
rect 798 986 801 1073
rect 810 1013 813 1186
rect 818 1123 821 1216
rect 826 1206 829 1726
rect 842 1703 845 1716
rect 834 1613 837 1626
rect 850 1603 853 1646
rect 858 1596 861 1886
rect 866 1793 869 1926
rect 874 1923 881 1926
rect 878 1866 881 1923
rect 890 1916 893 1943
rect 906 1923 909 1936
rect 890 1913 909 1916
rect 874 1863 881 1866
rect 866 1743 869 1776
rect 874 1726 877 1863
rect 882 1813 885 1846
rect 890 1813 893 1856
rect 906 1846 909 1866
rect 902 1843 909 1846
rect 870 1723 877 1726
rect 870 1626 873 1723
rect 882 1626 885 1746
rect 890 1703 893 1806
rect 902 1756 905 1843
rect 914 1813 917 1926
rect 922 1843 925 1953
rect 902 1753 909 1756
rect 870 1623 877 1626
rect 882 1623 893 1626
rect 898 1623 901 1736
rect 906 1716 909 1753
rect 914 1733 917 1806
rect 922 1793 925 1826
rect 930 1813 933 1936
rect 922 1716 925 1736
rect 930 1723 933 1756
rect 938 1733 941 1993
rect 946 1906 949 2133
rect 962 2106 965 2153
rect 970 2123 973 2156
rect 954 2013 957 2106
rect 962 2103 969 2106
rect 966 2026 969 2103
rect 978 2093 981 2216
rect 990 2166 993 2223
rect 986 2163 993 2166
rect 986 2116 989 2163
rect 994 2133 997 2146
rect 1002 2136 1005 2326
rect 1010 2286 1013 2336
rect 1018 2313 1021 2356
rect 1026 2293 1029 2336
rect 1010 2283 1029 2286
rect 1034 2273 1037 2426
rect 1042 2413 1045 2426
rect 1042 2323 1045 2406
rect 1034 2226 1037 2236
rect 1010 2223 1037 2226
rect 1010 2213 1013 2223
rect 1010 2143 1013 2206
rect 1018 2203 1021 2216
rect 1034 2166 1037 2206
rect 1042 2203 1045 2266
rect 1058 2256 1061 2433
rect 1114 2413 1117 2426
rect 1130 2413 1133 2496
rect 1138 2406 1141 2526
rect 1170 2516 1173 2563
rect 1162 2513 1173 2516
rect 1162 2493 1165 2513
rect 1146 2423 1149 2456
rect 1090 2393 1093 2406
rect 1082 2333 1085 2366
rect 1082 2306 1085 2326
rect 1090 2323 1093 2356
rect 1098 2323 1101 2406
rect 1138 2403 1149 2406
rect 1186 2386 1189 2566
rect 1202 2536 1205 2576
rect 1210 2573 1237 2576
rect 1202 2533 1213 2536
rect 1194 2516 1197 2526
rect 1202 2523 1213 2526
rect 1218 2523 1221 2566
rect 1226 2533 1229 2546
rect 1234 2523 1237 2573
rect 1242 2516 1245 2526
rect 1194 2513 1245 2516
rect 1250 2503 1253 2576
rect 1290 2533 1293 2566
rect 1306 2556 1309 2616
rect 1330 2603 1333 2616
rect 1378 2613 1381 2713
rect 1418 2636 1421 2923
rect 1426 2913 1429 2986
rect 1442 2973 1445 3006
rect 1434 2813 1437 2936
rect 1450 2926 1453 3016
rect 1458 3003 1461 3066
rect 1466 2993 1469 3006
rect 1474 2953 1477 3016
rect 1458 2933 1461 2946
rect 1482 2936 1485 3116
rect 1490 3093 1493 3126
rect 1506 3113 1509 3183
rect 1514 3166 1517 3206
rect 1522 3203 1541 3206
rect 1514 3163 1525 3166
rect 1522 3133 1525 3163
rect 1522 3113 1525 3126
rect 1538 3123 1541 3136
rect 1546 3133 1549 3206
rect 1554 3173 1557 3206
rect 1578 3186 1581 3206
rect 1586 3193 1589 3216
rect 1634 3213 1645 3216
rect 1658 3206 1661 3226
rect 1658 3203 1669 3206
rect 1602 3186 1605 3196
rect 1578 3183 1605 3186
rect 1554 3136 1557 3166
rect 1554 3133 1565 3136
rect 1498 3103 1517 3106
rect 1554 3103 1557 3126
rect 1490 2943 1493 3016
rect 1498 3013 1501 3066
rect 1506 2946 1509 3056
rect 1514 3013 1517 3103
rect 1522 3003 1525 3046
rect 1530 3013 1533 3056
rect 1538 3006 1541 3086
rect 1530 3003 1541 3006
rect 1506 2943 1517 2946
rect 1482 2933 1501 2936
rect 1442 2896 1445 2926
rect 1450 2923 1461 2926
rect 1466 2923 1493 2926
rect 1458 2913 1461 2923
rect 1498 2906 1501 2933
rect 1490 2903 1501 2906
rect 1442 2893 1453 2896
rect 1450 2836 1453 2893
rect 1442 2833 1453 2836
rect 1490 2836 1493 2903
rect 1514 2896 1517 2943
rect 1530 2913 1533 3003
rect 1546 2973 1549 3006
rect 1538 2933 1549 2936
rect 1506 2893 1517 2896
rect 1490 2833 1501 2836
rect 1442 2816 1445 2833
rect 1442 2813 1477 2816
rect 1442 2746 1445 2813
rect 1490 2793 1493 2806
rect 1442 2743 1453 2746
rect 1458 2723 1477 2726
rect 1474 2713 1477 2723
rect 1410 2633 1421 2636
rect 1298 2553 1309 2556
rect 1410 2556 1413 2633
rect 1426 2586 1429 2616
rect 1442 2603 1445 2616
rect 1482 2613 1485 2736
rect 1498 2723 1501 2833
rect 1506 2746 1509 2893
rect 1538 2856 1541 2926
rect 1546 2903 1549 2933
rect 1514 2853 1541 2856
rect 1514 2786 1517 2853
rect 1514 2783 1525 2786
rect 1506 2743 1517 2746
rect 1522 2743 1525 2783
rect 1530 2763 1533 2806
rect 1426 2583 1437 2586
rect 1410 2553 1421 2556
rect 1202 2393 1205 2486
rect 1186 2383 1197 2386
rect 1106 2313 1109 2376
rect 1114 2306 1117 2336
rect 1154 2333 1157 2356
rect 1082 2303 1117 2306
rect 1122 2303 1125 2326
rect 1138 2323 1157 2326
rect 1146 2313 1157 2316
rect 1082 2286 1085 2303
rect 1050 2253 1061 2256
rect 1074 2283 1085 2286
rect 1042 2166 1045 2176
rect 1034 2163 1045 2166
rect 1002 2133 1013 2136
rect 1026 2133 1029 2156
rect 1042 2143 1045 2163
rect 1050 2153 1053 2253
rect 1074 2236 1077 2283
rect 1090 2276 1093 2296
rect 1090 2273 1101 2276
rect 1058 2223 1061 2236
rect 1074 2233 1085 2236
rect 986 2113 993 2116
rect 962 2023 969 2026
rect 954 1923 957 1986
rect 946 1903 953 1906
rect 950 1826 953 1903
rect 946 1823 953 1826
rect 946 1756 949 1823
rect 962 1813 965 2023
rect 970 1973 973 2006
rect 978 1953 981 2056
rect 990 2026 993 2113
rect 1002 2103 1005 2126
rect 1010 2096 1013 2133
rect 1018 2113 1021 2126
rect 986 2023 993 2026
rect 1002 2093 1013 2096
rect 970 1923 973 1936
rect 978 1823 981 1946
rect 986 1893 989 2023
rect 1002 2013 1005 2093
rect 1010 2023 1013 2046
rect 994 1983 997 2006
rect 1010 1973 1013 2016
rect 1018 1966 1021 2006
rect 1002 1963 1021 1966
rect 986 1853 989 1886
rect 970 1813 981 1816
rect 954 1763 957 1806
rect 946 1753 957 1756
rect 938 1723 949 1726
rect 938 1716 941 1723
rect 906 1713 913 1716
rect 922 1713 941 1716
rect 910 1626 913 1713
rect 930 1646 933 1666
rect 906 1623 913 1626
rect 842 1593 861 1596
rect 834 1483 837 1546
rect 842 1533 845 1593
rect 866 1543 869 1606
rect 842 1416 845 1426
rect 834 1413 845 1416
rect 834 1346 837 1413
rect 842 1363 845 1406
rect 850 1403 853 1536
rect 858 1483 861 1536
rect 866 1523 869 1536
rect 858 1403 861 1416
rect 834 1343 861 1346
rect 834 1333 853 1336
rect 834 1303 837 1333
rect 858 1313 861 1343
rect 866 1313 869 1476
rect 826 1203 837 1206
rect 798 983 805 986
rect 818 983 821 1086
rect 794 933 797 966
rect 794 903 797 926
rect 794 823 797 846
rect 802 813 805 983
rect 810 876 813 966
rect 818 883 821 916
rect 810 873 821 876
rect 778 743 797 746
rect 754 733 765 736
rect 770 733 781 736
rect 770 683 773 726
rect 754 513 757 676
rect 778 646 781 733
rect 786 693 789 726
rect 794 686 797 743
rect 762 643 781 646
rect 786 683 797 686
rect 762 613 765 643
rect 770 613 773 636
rect 786 616 789 683
rect 778 613 789 616
rect 762 583 765 606
rect 778 583 781 613
rect 762 523 765 566
rect 754 413 757 426
rect 762 406 765 446
rect 770 413 773 436
rect 762 403 773 406
rect 778 403 781 516
rect 786 453 789 606
rect 794 533 797 606
rect 802 486 805 746
rect 810 573 813 806
rect 818 703 821 873
rect 818 563 821 616
rect 826 603 829 1203
rect 834 996 837 1136
rect 842 1026 845 1306
rect 850 1123 853 1156
rect 858 1143 861 1216
rect 866 1193 869 1266
rect 858 1103 861 1126
rect 866 1096 869 1116
rect 850 1093 869 1096
rect 842 1023 853 1026
rect 842 1003 845 1016
rect 834 993 845 996
rect 834 923 837 946
rect 834 903 837 916
rect 834 573 837 896
rect 842 726 845 936
rect 850 923 853 1023
rect 874 1006 877 1623
rect 882 1473 885 1616
rect 882 1273 885 1416
rect 882 1233 885 1246
rect 882 1173 885 1226
rect 882 1123 885 1136
rect 890 1106 893 1623
rect 906 1603 909 1623
rect 922 1613 925 1646
rect 930 1643 937 1646
rect 898 1233 901 1536
rect 906 1506 909 1596
rect 914 1563 917 1606
rect 922 1556 925 1596
rect 934 1556 937 1643
rect 914 1553 925 1556
rect 930 1553 937 1556
rect 914 1523 917 1553
rect 922 1533 925 1546
rect 906 1503 917 1506
rect 914 1446 917 1503
rect 930 1453 933 1553
rect 938 1513 941 1536
rect 946 1523 949 1676
rect 954 1603 957 1753
rect 962 1723 965 1776
rect 970 1716 973 1746
rect 978 1733 981 1806
rect 986 1803 989 1826
rect 986 1726 989 1776
rect 994 1743 997 1936
rect 962 1713 973 1716
rect 978 1723 989 1726
rect 1002 1723 1005 1963
rect 1026 1956 1029 2086
rect 1042 2053 1045 2136
rect 1042 2013 1045 2026
rect 1010 1953 1029 1956
rect 1010 1836 1013 1953
rect 1042 1946 1045 1986
rect 1026 1943 1045 1946
rect 1018 1853 1021 1936
rect 1026 1923 1029 1943
rect 1042 1923 1045 1936
rect 1050 1916 1053 2126
rect 1058 2123 1061 2206
rect 1066 2203 1069 2216
rect 1066 2116 1069 2166
rect 1074 2153 1077 2216
rect 1082 2143 1085 2233
rect 1098 2226 1101 2273
rect 1094 2223 1101 2226
rect 1094 2136 1097 2223
rect 1106 2193 1109 2206
rect 1074 2133 1085 2136
rect 1090 2133 1097 2136
rect 1090 2116 1093 2133
rect 1106 2116 1109 2136
rect 1114 2133 1117 2216
rect 1122 2213 1133 2216
rect 1122 2163 1125 2206
rect 1130 2183 1133 2206
rect 1138 2176 1141 2226
rect 1130 2173 1141 2176
rect 1066 2113 1077 2116
rect 1058 2013 1061 2086
rect 1074 2026 1077 2113
rect 1086 2113 1093 2116
rect 1086 2036 1089 2113
rect 1086 2033 1093 2036
rect 1066 2023 1077 2026
rect 1034 1913 1053 1916
rect 1010 1833 1017 1836
rect 1014 1766 1017 1833
rect 1026 1813 1029 1846
rect 1010 1763 1017 1766
rect 1010 1743 1013 1763
rect 1026 1733 1029 1786
rect 1034 1773 1037 1913
rect 1042 1803 1045 1886
rect 1042 1766 1045 1796
rect 1050 1773 1053 1856
rect 1058 1766 1061 1936
rect 1066 1923 1069 2023
rect 1090 2013 1093 2033
rect 1098 2013 1101 2116
rect 1106 2113 1113 2116
rect 1110 2046 1113 2113
rect 1122 2083 1125 2126
rect 1106 2043 1113 2046
rect 1106 2006 1109 2043
rect 1082 2003 1109 2006
rect 1074 1883 1077 1966
rect 1106 1963 1109 2003
rect 1082 1926 1085 1946
rect 1098 1926 1101 1946
rect 1082 1923 1093 1926
rect 1098 1923 1105 1926
rect 1090 1876 1093 1923
rect 1074 1873 1093 1876
rect 1034 1736 1037 1766
rect 1042 1763 1061 1766
rect 1066 1756 1069 1856
rect 1050 1753 1069 1756
rect 1034 1733 1045 1736
rect 1018 1723 1037 1726
rect 914 1443 933 1446
rect 906 1423 909 1436
rect 906 1333 909 1346
rect 914 1313 917 1406
rect 898 1143 901 1186
rect 886 1103 893 1106
rect 886 1016 889 1103
rect 886 1013 893 1016
rect 898 1013 901 1116
rect 906 1083 909 1276
rect 922 1256 925 1406
rect 914 1253 925 1256
rect 914 1063 917 1253
rect 906 1013 909 1056
rect 866 1003 877 1006
rect 866 956 869 1003
rect 866 953 877 956
rect 858 883 861 916
rect 866 913 869 936
rect 874 896 877 953
rect 882 943 885 996
rect 870 893 877 896
rect 850 743 853 826
rect 858 803 861 846
rect 870 796 873 893
rect 882 823 885 896
rect 890 853 893 1013
rect 906 936 909 1006
rect 914 983 917 1006
rect 906 933 913 936
rect 898 843 901 926
rect 910 856 913 933
rect 906 853 913 856
rect 906 833 909 853
rect 870 793 877 796
rect 842 723 849 726
rect 846 626 849 723
rect 858 703 861 736
rect 866 733 869 776
rect 866 693 869 726
rect 874 676 877 793
rect 882 763 885 806
rect 870 673 877 676
rect 842 623 849 626
rect 810 503 813 546
rect 826 523 829 556
rect 794 483 805 486
rect 738 316 741 346
rect 722 313 741 316
rect 746 306 749 336
rect 714 303 749 306
rect 754 323 765 326
rect 754 286 757 323
rect 770 316 773 403
rect 674 243 685 246
rect 746 283 757 286
rect 762 313 773 316
rect 674 183 677 243
rect 746 236 749 283
rect 746 233 757 236
rect 682 223 709 226
rect 522 123 533 126
rect 538 116 541 126
rect 506 113 541 116
rect 570 123 577 126
rect 586 133 597 136
rect 570 53 573 123
rect 586 113 589 133
rect 666 123 669 156
rect 682 133 685 176
rect 690 163 693 216
rect 706 213 709 223
rect 754 213 757 233
rect 698 203 709 206
rect 722 193 725 206
rect 722 143 741 146
rect 722 133 725 143
rect 722 113 725 126
rect 730 116 733 136
rect 738 123 741 143
rect 746 116 749 176
rect 754 123 757 166
rect 762 153 765 313
rect 786 273 789 416
rect 794 403 797 483
rect 818 476 821 496
rect 834 493 837 536
rect 842 486 845 623
rect 814 473 821 476
rect 826 483 845 486
rect 802 393 805 456
rect 814 386 817 473
rect 814 383 821 386
rect 810 333 813 366
rect 818 323 821 383
rect 826 333 829 483
rect 834 323 837 416
rect 850 396 853 606
rect 858 603 861 626
rect 870 596 873 673
rect 882 623 885 726
rect 882 606 885 616
rect 890 613 893 806
rect 914 803 917 816
rect 898 703 901 716
rect 906 673 909 736
rect 906 606 909 626
rect 914 623 917 726
rect 882 603 909 606
rect 870 593 877 596
rect 858 523 861 546
rect 866 513 869 536
rect 866 413 869 446
rect 874 413 877 593
rect 906 533 909 603
rect 882 463 885 526
rect 914 516 917 606
rect 922 533 925 1246
rect 930 1183 933 1443
rect 938 1413 941 1426
rect 938 1393 941 1406
rect 930 1123 933 1166
rect 938 1116 941 1336
rect 946 1223 949 1446
rect 954 1333 957 1506
rect 962 1403 965 1713
rect 970 1613 973 1646
rect 962 1383 965 1396
rect 946 1173 949 1216
rect 934 1113 941 1116
rect 934 1026 937 1113
rect 930 1023 937 1026
rect 930 983 933 1023
rect 946 996 949 1166
rect 954 1106 957 1296
rect 962 1243 965 1336
rect 970 1293 973 1606
rect 978 1553 981 1723
rect 1034 1703 1037 1723
rect 986 1596 989 1696
rect 994 1603 997 1656
rect 1002 1623 1021 1626
rect 1018 1616 1021 1623
rect 1002 1603 1005 1616
rect 1010 1596 1013 1616
rect 1018 1613 1029 1616
rect 986 1593 1013 1596
rect 1002 1546 1005 1566
rect 994 1543 1005 1546
rect 978 1533 997 1536
rect 978 1503 981 1533
rect 1002 1526 1005 1543
rect 986 1493 989 1516
rect 978 1236 981 1416
rect 986 1413 989 1456
rect 994 1423 997 1526
rect 1002 1523 1009 1526
rect 1006 1456 1009 1523
rect 1002 1453 1009 1456
rect 986 1383 989 1406
rect 986 1263 989 1336
rect 962 1233 981 1236
rect 962 1213 965 1233
rect 994 1226 997 1416
rect 1002 1403 1005 1453
rect 1010 1413 1013 1436
rect 1018 1406 1021 1556
rect 1026 1453 1029 1606
rect 1034 1546 1037 1606
rect 1042 1563 1045 1733
rect 1034 1543 1045 1546
rect 1010 1403 1021 1406
rect 978 1223 997 1226
rect 978 1213 981 1223
rect 962 1126 965 1186
rect 970 1133 973 1206
rect 978 1143 981 1166
rect 962 1123 973 1126
rect 954 1103 965 1106
rect 962 1036 965 1103
rect 938 993 949 996
rect 954 1033 965 1036
rect 938 966 941 993
rect 930 963 941 966
rect 930 926 933 963
rect 938 933 941 956
rect 930 923 941 926
rect 946 923 949 986
rect 930 823 933 866
rect 930 583 933 756
rect 938 723 941 923
rect 946 803 949 886
rect 954 733 957 1033
rect 978 1003 981 1016
rect 962 933 965 966
rect 962 763 965 916
rect 970 893 973 996
rect 986 976 989 1216
rect 994 1123 997 1223
rect 994 1013 997 1036
rect 994 983 997 1006
rect 986 973 993 976
rect 978 846 981 936
rect 990 866 993 973
rect 990 863 997 866
rect 970 843 981 846
rect 970 796 973 843
rect 986 813 989 846
rect 970 793 989 796
rect 994 793 997 863
rect 1002 823 1005 1346
rect 1010 1173 1013 1403
rect 1026 1386 1029 1426
rect 1022 1383 1029 1386
rect 1022 1336 1025 1383
rect 1034 1343 1037 1526
rect 1022 1333 1029 1336
rect 1018 1203 1021 1306
rect 1026 1263 1029 1333
rect 1042 1326 1045 1543
rect 1050 1506 1053 1753
rect 1058 1733 1061 1746
rect 1058 1676 1061 1696
rect 1058 1673 1065 1676
rect 1062 1576 1065 1673
rect 1074 1606 1077 1873
rect 1102 1856 1105 1923
rect 1098 1853 1105 1856
rect 1114 1853 1117 2026
rect 1122 2006 1125 2016
rect 1130 2013 1133 2173
rect 1138 2073 1141 2126
rect 1146 2116 1149 2313
rect 1162 2306 1165 2336
rect 1158 2303 1165 2306
rect 1158 2236 1161 2303
rect 1194 2286 1197 2383
rect 1218 2326 1221 2346
rect 1214 2323 1221 2326
rect 1194 2283 1205 2286
rect 1154 2233 1161 2236
rect 1154 2203 1157 2233
rect 1154 2133 1157 2146
rect 1162 2123 1165 2216
rect 1146 2113 1153 2116
rect 1150 2066 1153 2113
rect 1146 2063 1153 2066
rect 1146 2013 1149 2063
rect 1162 2013 1165 2096
rect 1170 2006 1173 2276
rect 1122 2003 1133 2006
rect 1122 1923 1125 1986
rect 1130 1926 1133 2003
rect 1154 1983 1157 2006
rect 1162 2003 1173 2006
rect 1138 1933 1141 1946
rect 1130 1923 1141 1926
rect 1098 1833 1101 1853
rect 1122 1836 1125 1916
rect 1138 1913 1141 1923
rect 1146 1906 1149 1946
rect 1118 1833 1125 1836
rect 1130 1903 1149 1906
rect 1082 1783 1085 1826
rect 1098 1823 1109 1826
rect 1090 1746 1093 1816
rect 1118 1786 1121 1833
rect 1130 1793 1133 1903
rect 1138 1846 1141 1866
rect 1146 1856 1149 1903
rect 1154 1896 1157 1926
rect 1162 1923 1165 2003
rect 1154 1893 1165 1896
rect 1154 1863 1157 1886
rect 1146 1853 1157 1856
rect 1138 1843 1149 1846
rect 1146 1813 1149 1843
rect 1154 1813 1157 1853
rect 1162 1806 1165 1893
rect 1118 1783 1125 1786
rect 1090 1743 1101 1746
rect 1082 1613 1085 1736
rect 1098 1723 1101 1743
rect 1090 1626 1093 1676
rect 1114 1663 1117 1726
rect 1114 1636 1117 1656
rect 1098 1633 1117 1636
rect 1090 1623 1101 1626
rect 1090 1606 1093 1616
rect 1074 1603 1093 1606
rect 1098 1603 1101 1623
rect 1106 1603 1109 1633
rect 1114 1623 1117 1633
rect 1058 1573 1065 1576
rect 1058 1523 1061 1573
rect 1066 1533 1069 1556
rect 1082 1526 1085 1536
rect 1090 1533 1093 1586
rect 1050 1503 1061 1506
rect 1058 1456 1061 1503
rect 1074 1493 1077 1526
rect 1082 1523 1093 1526
rect 1090 1513 1093 1523
rect 1050 1453 1061 1456
rect 1050 1433 1053 1453
rect 1038 1323 1045 1326
rect 1038 1236 1041 1323
rect 1050 1303 1053 1406
rect 1066 1356 1069 1416
rect 1074 1366 1077 1476
rect 1098 1473 1101 1536
rect 1082 1413 1085 1426
rect 1090 1403 1093 1436
rect 1106 1433 1109 1526
rect 1114 1516 1117 1576
rect 1122 1533 1125 1783
rect 1130 1676 1133 1726
rect 1138 1693 1141 1736
rect 1146 1723 1149 1806
rect 1154 1803 1165 1806
rect 1154 1706 1157 1746
rect 1150 1703 1157 1706
rect 1130 1673 1137 1676
rect 1134 1576 1137 1673
rect 1150 1616 1153 1703
rect 1150 1613 1157 1616
rect 1146 1583 1149 1596
rect 1134 1573 1141 1576
rect 1114 1513 1121 1516
rect 1118 1426 1121 1513
rect 1074 1363 1081 1366
rect 1058 1353 1069 1356
rect 1058 1303 1061 1353
rect 1066 1313 1069 1346
rect 1038 1233 1045 1236
rect 1042 1216 1045 1233
rect 1034 1213 1045 1216
rect 1050 1213 1053 1256
rect 1026 1143 1029 1206
rect 1010 1033 1013 1136
rect 1034 1126 1037 1176
rect 1030 1123 1037 1126
rect 1018 1023 1021 1056
rect 1030 1026 1033 1123
rect 1042 1093 1045 1126
rect 1050 1123 1053 1166
rect 1058 1153 1061 1246
rect 1066 1213 1069 1276
rect 1078 1226 1081 1363
rect 1090 1333 1093 1346
rect 1074 1223 1081 1226
rect 1074 1206 1077 1223
rect 1090 1213 1093 1326
rect 1066 1203 1077 1206
rect 1030 1023 1037 1026
rect 1010 913 1013 1016
rect 1018 923 1021 946
rect 986 746 989 793
rect 986 743 1005 746
rect 1010 743 1013 826
rect 1018 813 1021 916
rect 1018 786 1021 806
rect 1026 803 1029 1006
rect 1034 913 1037 1023
rect 1034 803 1037 826
rect 1042 786 1045 1086
rect 1058 1076 1061 1146
rect 1066 1083 1069 1203
rect 1074 1183 1077 1196
rect 1074 1133 1085 1136
rect 1090 1133 1093 1196
rect 1018 783 1029 786
rect 978 716 981 736
rect 1026 716 1029 783
rect 962 713 981 716
rect 1018 713 1029 716
rect 1038 783 1045 786
rect 1050 1073 1061 1076
rect 938 613 941 676
rect 962 646 965 713
rect 954 643 965 646
rect 954 623 957 643
rect 954 556 957 616
rect 954 553 973 556
rect 930 543 957 546
rect 930 533 933 543
rect 938 533 949 536
rect 954 533 957 543
rect 910 513 917 516
rect 910 446 913 513
rect 882 423 893 426
rect 842 393 853 396
rect 770 146 773 246
rect 842 226 845 393
rect 850 323 853 376
rect 858 333 861 346
rect 866 316 869 406
rect 882 386 885 423
rect 890 403 893 416
rect 898 413 901 446
rect 910 443 917 446
rect 914 426 917 443
rect 922 433 925 526
rect 938 506 941 526
rect 946 523 957 526
rect 934 503 941 506
rect 934 446 937 503
rect 954 476 957 523
rect 970 486 973 553
rect 986 533 989 626
rect 1010 613 1013 696
rect 1002 563 1005 606
rect 946 473 957 476
rect 962 483 973 486
rect 946 453 949 473
rect 962 466 965 483
rect 954 463 965 466
rect 934 443 941 446
rect 914 423 933 426
rect 906 406 909 416
rect 898 403 909 406
rect 882 383 893 386
rect 874 333 877 366
rect 890 326 893 383
rect 862 313 869 316
rect 826 223 845 226
rect 778 183 781 206
rect 762 143 773 146
rect 762 123 765 143
rect 802 133 805 216
rect 810 176 813 216
rect 826 203 829 216
rect 850 203 853 266
rect 810 173 821 176
rect 730 113 749 116
rect 818 116 821 173
rect 862 156 865 313
rect 862 153 869 156
rect 826 143 845 146
rect 826 123 829 143
rect 834 116 837 136
rect 842 133 845 143
rect 858 123 861 136
rect 866 123 869 153
rect 874 123 877 326
rect 882 323 893 326
rect 882 303 885 323
rect 906 216 909 266
rect 914 223 917 336
rect 930 246 933 423
rect 938 413 941 443
rect 922 243 933 246
rect 922 233 925 243
rect 930 223 933 236
rect 890 133 893 216
rect 906 213 925 216
rect 938 183 941 336
rect 946 316 949 426
rect 954 363 957 463
rect 970 456 973 466
rect 962 453 973 456
rect 962 413 965 453
rect 986 446 989 526
rect 1002 513 1005 526
rect 1010 456 1013 586
rect 1018 536 1021 713
rect 1038 696 1041 783
rect 1026 693 1041 696
rect 1050 696 1053 1073
rect 1058 1033 1061 1066
rect 1058 1003 1061 1016
rect 1074 993 1077 1133
rect 1082 1123 1093 1126
rect 1082 1023 1085 1116
rect 1098 1046 1101 1416
rect 1106 1413 1109 1426
rect 1114 1423 1121 1426
rect 1106 1373 1109 1406
rect 1106 1113 1109 1336
rect 1094 1043 1101 1046
rect 1058 943 1085 946
rect 1058 923 1061 943
rect 1066 893 1069 936
rect 1074 906 1077 926
rect 1082 923 1085 943
rect 1094 926 1097 1043
rect 1106 936 1109 1036
rect 1114 1033 1117 1423
rect 1130 1413 1133 1566
rect 1138 1516 1141 1573
rect 1138 1513 1145 1516
rect 1154 1513 1157 1613
rect 1142 1446 1145 1513
rect 1142 1443 1149 1446
rect 1138 1406 1141 1426
rect 1130 1403 1141 1406
rect 1122 1323 1125 1376
rect 1130 1303 1133 1403
rect 1122 1176 1125 1226
rect 1138 1213 1141 1346
rect 1146 1273 1149 1443
rect 1138 1176 1141 1196
rect 1146 1183 1149 1206
rect 1122 1173 1133 1176
rect 1138 1173 1149 1176
rect 1122 1133 1125 1166
rect 1130 1086 1133 1173
rect 1122 1083 1133 1086
rect 1122 1016 1125 1083
rect 1118 1013 1125 1016
rect 1118 956 1121 1013
rect 1130 963 1133 1066
rect 1118 953 1125 956
rect 1106 933 1113 936
rect 1094 923 1101 926
rect 1074 903 1093 906
rect 1058 823 1061 836
rect 1058 753 1061 806
rect 1066 786 1069 826
rect 1074 803 1077 816
rect 1066 783 1077 786
rect 1058 733 1061 746
rect 1058 703 1061 726
rect 1066 706 1069 736
rect 1074 723 1077 783
rect 1082 716 1085 896
rect 1090 783 1093 903
rect 1098 836 1101 923
rect 1110 886 1113 933
rect 1106 883 1113 886
rect 1106 853 1109 883
rect 1098 833 1105 836
rect 1090 723 1093 756
rect 1102 736 1105 833
rect 1098 733 1105 736
rect 1082 713 1093 716
rect 1066 703 1085 706
rect 1050 693 1069 696
rect 1026 633 1029 693
rect 1026 553 1029 616
rect 1018 533 1029 536
rect 1018 463 1021 526
rect 1026 496 1029 533
rect 1034 513 1037 646
rect 1042 623 1045 686
rect 1042 613 1053 616
rect 1058 576 1061 626
rect 1026 493 1033 496
rect 1010 453 1021 456
rect 986 443 997 446
rect 970 393 973 406
rect 978 383 981 416
rect 994 413 997 443
rect 986 346 989 406
rect 954 343 989 346
rect 954 323 957 343
rect 962 323 965 336
rect 986 333 989 343
rect 978 316 981 326
rect 994 323 997 356
rect 946 313 981 316
rect 1002 293 1005 406
rect 1010 393 1013 416
rect 1018 286 1021 453
rect 1030 376 1033 493
rect 1042 396 1045 576
rect 1050 573 1061 576
rect 1050 533 1053 573
rect 1066 566 1069 693
rect 1074 613 1077 656
rect 1058 563 1069 566
rect 1058 533 1061 563
rect 1074 533 1077 556
rect 1050 496 1053 516
rect 1050 493 1061 496
rect 1058 426 1061 493
rect 1050 423 1061 426
rect 1050 403 1053 423
rect 1042 393 1053 396
rect 1030 373 1037 376
rect 1014 283 1021 286
rect 1014 236 1017 283
rect 1034 276 1037 373
rect 1050 316 1053 393
rect 1050 313 1061 316
rect 1026 273 1037 276
rect 1026 253 1029 273
rect 946 223 949 236
rect 954 223 957 236
rect 1014 233 1021 236
rect 986 213 989 226
rect 818 113 837 116
rect 898 73 901 146
rect 1002 133 1005 226
rect 1010 173 1013 216
rect 1018 203 1021 233
rect 1050 223 1053 306
rect 1050 166 1053 216
rect 1058 203 1061 313
rect 1074 226 1077 516
rect 1082 513 1085 646
rect 1090 636 1093 713
rect 1098 676 1101 733
rect 1106 683 1109 716
rect 1098 673 1109 676
rect 1106 653 1109 673
rect 1090 633 1101 636
rect 1098 586 1101 633
rect 1114 606 1117 866
rect 1122 813 1125 953
rect 1130 913 1133 936
rect 1122 743 1125 806
rect 1122 723 1125 736
rect 1122 613 1125 706
rect 1130 623 1133 836
rect 1138 693 1141 1136
rect 1146 1123 1149 1173
rect 1154 1136 1157 1426
rect 1162 1193 1165 1803
rect 1170 1723 1173 1976
rect 1170 1613 1173 1666
rect 1178 1546 1181 2266
rect 1186 2223 1189 2236
rect 1186 2193 1189 2206
rect 1194 2173 1197 2206
rect 1202 2196 1205 2283
rect 1214 2246 1217 2323
rect 1234 2316 1237 2496
rect 1266 2493 1269 2526
rect 1250 2393 1253 2416
rect 1242 2343 1253 2346
rect 1242 2333 1245 2343
rect 1214 2243 1221 2246
rect 1210 2213 1213 2226
rect 1202 2193 1209 2196
rect 1186 2103 1189 2116
rect 1194 2086 1197 2136
rect 1206 2116 1209 2193
rect 1186 2083 1197 2086
rect 1202 2113 1209 2116
rect 1186 2003 1189 2083
rect 1194 2013 1197 2026
rect 1202 2006 1205 2113
rect 1218 2096 1221 2243
rect 1226 2213 1229 2316
rect 1234 2313 1245 2316
rect 1266 2313 1269 2376
rect 1274 2333 1277 2416
rect 1282 2413 1285 2526
rect 1298 2523 1301 2553
rect 1314 2513 1317 2536
rect 1362 2486 1365 2526
rect 1410 2503 1413 2536
rect 1418 2486 1421 2553
rect 1426 2533 1429 2556
rect 1362 2483 1381 2486
rect 1290 2413 1293 2426
rect 1314 2403 1317 2426
rect 1354 2413 1357 2426
rect 1338 2393 1341 2406
rect 1362 2393 1365 2406
rect 1242 2236 1245 2313
rect 1234 2233 1245 2236
rect 1234 2213 1237 2233
rect 1226 2203 1237 2206
rect 1194 2003 1205 2006
rect 1210 2093 1221 2096
rect 1186 1756 1189 1946
rect 1194 1923 1197 2003
rect 1194 1793 1197 1856
rect 1186 1753 1197 1756
rect 1186 1733 1189 1746
rect 1186 1663 1189 1726
rect 1194 1716 1197 1753
rect 1202 1733 1205 1936
rect 1210 1896 1213 2093
rect 1218 2013 1221 2086
rect 1218 1916 1221 1926
rect 1226 1923 1229 2146
rect 1234 2036 1237 2203
rect 1242 2093 1245 2216
rect 1250 2183 1253 2216
rect 1258 2133 1261 2146
rect 1258 2116 1261 2126
rect 1266 2123 1269 2306
rect 1282 2253 1309 2256
rect 1282 2236 1285 2253
rect 1278 2233 1285 2236
rect 1278 2156 1281 2233
rect 1278 2153 1285 2156
rect 1282 2116 1285 2153
rect 1258 2113 1285 2116
rect 1290 2066 1293 2216
rect 1298 2146 1301 2246
rect 1306 2223 1309 2253
rect 1306 2163 1309 2206
rect 1298 2143 1309 2146
rect 1298 2113 1301 2136
rect 1306 2133 1309 2143
rect 1286 2063 1293 2066
rect 1234 2033 1253 2036
rect 1234 1943 1237 2016
rect 1242 1996 1245 2006
rect 1250 2003 1253 2033
rect 1258 2013 1261 2026
rect 1286 2016 1289 2063
rect 1242 1993 1253 1996
rect 1218 1913 1229 1916
rect 1210 1893 1221 1896
rect 1218 1836 1221 1893
rect 1218 1833 1229 1836
rect 1218 1813 1221 1826
rect 1210 1793 1213 1806
rect 1226 1796 1229 1833
rect 1234 1823 1237 1926
rect 1250 1916 1253 1993
rect 1266 1983 1269 2006
rect 1274 1926 1277 2016
rect 1286 2013 1293 2016
rect 1282 1963 1285 1996
rect 1246 1913 1253 1916
rect 1246 1846 1249 1913
rect 1258 1906 1261 1926
rect 1274 1923 1285 1926
rect 1258 1903 1269 1906
rect 1242 1843 1249 1846
rect 1242 1813 1245 1843
rect 1226 1793 1237 1796
rect 1210 1733 1213 1776
rect 1194 1713 1201 1716
rect 1210 1713 1213 1726
rect 1198 1636 1201 1713
rect 1218 1703 1221 1736
rect 1194 1633 1201 1636
rect 1186 1603 1189 1626
rect 1194 1613 1197 1633
rect 1210 1623 1221 1626
rect 1194 1576 1197 1606
rect 1202 1603 1205 1616
rect 1210 1613 1221 1616
rect 1194 1573 1205 1576
rect 1170 1543 1181 1546
rect 1170 1506 1173 1543
rect 1186 1536 1189 1546
rect 1178 1533 1189 1536
rect 1194 1533 1197 1566
rect 1202 1543 1205 1573
rect 1170 1503 1181 1506
rect 1170 1403 1173 1496
rect 1178 1423 1181 1503
rect 1186 1416 1189 1526
rect 1202 1493 1205 1536
rect 1210 1533 1213 1556
rect 1218 1506 1221 1613
rect 1226 1603 1229 1786
rect 1234 1583 1237 1793
rect 1242 1643 1245 1806
rect 1250 1786 1253 1826
rect 1258 1793 1261 1826
rect 1266 1803 1269 1903
rect 1250 1783 1261 1786
rect 1274 1783 1277 1916
rect 1282 1903 1285 1923
rect 1282 1793 1285 1896
rect 1250 1623 1253 1736
rect 1258 1713 1261 1783
rect 1290 1776 1293 2013
rect 1286 1773 1293 1776
rect 1266 1723 1269 1766
rect 1274 1723 1277 1746
rect 1258 1686 1261 1706
rect 1258 1683 1269 1686
rect 1266 1636 1269 1683
rect 1286 1666 1289 1773
rect 1298 1683 1301 2056
rect 1306 2013 1309 2046
rect 1314 2003 1317 2336
rect 1330 2326 1333 2336
rect 1338 2333 1341 2366
rect 1370 2356 1373 2416
rect 1378 2406 1381 2483
rect 1410 2483 1421 2486
rect 1386 2423 1389 2436
rect 1410 2406 1413 2483
rect 1426 2413 1429 2526
rect 1434 2523 1437 2583
rect 1466 2513 1469 2536
rect 1490 2476 1493 2526
rect 1466 2473 1493 2476
rect 1378 2403 1389 2406
rect 1394 2393 1397 2406
rect 1410 2403 1421 2406
rect 1418 2356 1421 2403
rect 1370 2353 1421 2356
rect 1322 2323 1341 2326
rect 1330 2203 1333 2296
rect 1338 2233 1341 2316
rect 1346 2293 1349 2336
rect 1370 2333 1373 2346
rect 1362 2323 1373 2326
rect 1354 2246 1357 2316
rect 1378 2303 1381 2336
rect 1354 2243 1381 2246
rect 1322 2173 1325 2196
rect 1330 2193 1341 2196
rect 1306 1773 1309 1936
rect 1314 1923 1317 1946
rect 1314 1763 1317 1906
rect 1286 1663 1293 1666
rect 1258 1633 1269 1636
rect 1258 1616 1261 1633
rect 1250 1613 1261 1616
rect 1242 1576 1245 1606
rect 1250 1576 1253 1613
rect 1210 1503 1221 1506
rect 1210 1446 1213 1503
rect 1178 1413 1189 1416
rect 1194 1443 1213 1446
rect 1170 1333 1173 1386
rect 1178 1326 1181 1413
rect 1186 1373 1189 1406
rect 1178 1323 1189 1326
rect 1154 1133 1165 1136
rect 1154 1116 1157 1126
rect 1146 1113 1157 1116
rect 1146 863 1149 1113
rect 1162 1106 1165 1133
rect 1154 1103 1165 1106
rect 1154 913 1157 1103
rect 1170 1093 1173 1256
rect 1162 1013 1165 1036
rect 1162 983 1165 1006
rect 1170 1003 1173 1016
rect 1178 986 1181 1306
rect 1186 1213 1189 1226
rect 1186 1123 1189 1196
rect 1186 1066 1189 1116
rect 1194 1073 1197 1443
rect 1210 1416 1213 1436
rect 1218 1423 1221 1496
rect 1234 1486 1237 1576
rect 1242 1573 1253 1576
rect 1226 1483 1237 1486
rect 1202 1303 1205 1416
rect 1210 1413 1221 1416
rect 1218 1403 1221 1413
rect 1210 1243 1213 1366
rect 1202 1186 1205 1236
rect 1202 1183 1209 1186
rect 1206 1126 1209 1183
rect 1206 1123 1213 1126
rect 1202 1066 1205 1116
rect 1186 1063 1205 1066
rect 1186 1023 1189 1036
rect 1194 1013 1197 1063
rect 1210 1033 1213 1123
rect 1218 1113 1221 1386
rect 1194 996 1197 1006
rect 1174 983 1181 986
rect 1186 993 1197 996
rect 1154 756 1157 806
rect 1162 796 1165 966
rect 1174 926 1177 983
rect 1186 933 1189 993
rect 1174 923 1181 926
rect 1170 803 1173 826
rect 1178 813 1181 923
rect 1162 793 1189 796
rect 1146 753 1157 756
rect 1146 713 1149 753
rect 1154 743 1173 746
rect 1090 583 1101 586
rect 1110 603 1117 606
rect 1090 563 1093 583
rect 1110 536 1113 603
rect 1122 576 1125 606
rect 1122 573 1133 576
rect 1106 533 1113 536
rect 1122 533 1125 566
rect 1130 533 1133 573
rect 1090 406 1093 456
rect 1098 433 1101 526
rect 1086 403 1093 406
rect 1086 316 1089 403
rect 1098 383 1101 416
rect 1106 343 1109 533
rect 1146 526 1149 686
rect 1154 533 1157 743
rect 1170 736 1173 743
rect 1162 716 1165 736
rect 1170 733 1181 736
rect 1186 723 1189 793
rect 1194 733 1197 916
rect 1202 843 1205 1016
rect 1226 1013 1229 1483
rect 1234 1393 1237 1476
rect 1242 1413 1245 1566
rect 1234 1006 1237 1336
rect 1242 1266 1245 1406
rect 1250 1283 1253 1573
rect 1258 1566 1261 1596
rect 1266 1583 1269 1606
rect 1258 1563 1277 1566
rect 1282 1563 1285 1646
rect 1290 1573 1293 1663
rect 1298 1623 1301 1656
rect 1298 1566 1301 1616
rect 1306 1583 1309 1696
rect 1314 1573 1317 1736
rect 1290 1563 1301 1566
rect 1258 1373 1261 1556
rect 1274 1546 1277 1563
rect 1266 1473 1269 1546
rect 1274 1543 1285 1546
rect 1290 1543 1293 1563
rect 1298 1543 1317 1546
rect 1266 1383 1269 1456
rect 1258 1336 1261 1366
rect 1258 1333 1269 1336
rect 1274 1333 1277 1536
rect 1282 1486 1285 1543
rect 1290 1523 1293 1536
rect 1298 1526 1301 1536
rect 1298 1523 1317 1526
rect 1282 1483 1293 1486
rect 1282 1343 1285 1426
rect 1266 1323 1269 1333
rect 1258 1313 1269 1316
rect 1242 1263 1249 1266
rect 1246 1196 1249 1263
rect 1258 1203 1261 1313
rect 1274 1306 1277 1326
rect 1266 1303 1277 1306
rect 1266 1213 1269 1303
rect 1274 1203 1277 1266
rect 1246 1193 1261 1196
rect 1218 1003 1237 1006
rect 1210 983 1213 996
rect 1210 923 1213 976
rect 1210 893 1213 916
rect 1218 913 1221 1003
rect 1226 896 1229 936
rect 1234 923 1237 996
rect 1222 893 1229 896
rect 1222 826 1225 893
rect 1210 823 1225 826
rect 1162 713 1169 716
rect 1202 713 1205 786
rect 1166 636 1169 713
rect 1162 633 1169 636
rect 1162 613 1165 633
rect 1170 603 1173 616
rect 1114 506 1117 526
rect 1122 523 1133 526
rect 1138 513 1141 526
rect 1146 523 1157 526
rect 1114 503 1125 506
rect 1122 426 1125 503
rect 1114 423 1125 426
rect 1114 403 1117 423
rect 1098 323 1101 336
rect 1106 323 1109 336
rect 1122 333 1125 396
rect 1130 333 1133 356
rect 1114 323 1125 326
rect 1122 316 1125 323
rect 1138 316 1141 426
rect 1154 396 1157 523
rect 1170 433 1173 536
rect 1178 416 1181 706
rect 1202 616 1205 676
rect 1194 613 1205 616
rect 1186 516 1189 566
rect 1194 526 1197 613
rect 1202 593 1205 606
rect 1202 533 1205 586
rect 1194 523 1205 526
rect 1186 513 1197 516
rect 1186 423 1197 426
rect 1178 413 1197 416
rect 1202 413 1205 523
rect 1210 453 1213 823
rect 1218 813 1229 816
rect 1218 763 1221 806
rect 1218 683 1221 736
rect 1226 703 1229 813
rect 1218 593 1221 616
rect 1226 603 1229 676
rect 1234 586 1237 916
rect 1230 583 1237 586
rect 1218 473 1221 526
rect 1230 456 1233 583
rect 1242 566 1245 1136
rect 1250 843 1253 1126
rect 1250 733 1253 806
rect 1250 703 1253 726
rect 1250 573 1253 606
rect 1242 563 1253 566
rect 1242 533 1245 556
rect 1250 526 1253 563
rect 1242 523 1253 526
rect 1242 473 1245 523
rect 1258 513 1261 1193
rect 1266 1133 1269 1156
rect 1266 1093 1269 1116
rect 1266 993 1269 1036
rect 1274 993 1277 1146
rect 1282 1063 1285 1326
rect 1290 1253 1293 1483
rect 1298 1423 1301 1523
rect 1306 1426 1309 1456
rect 1314 1433 1317 1476
rect 1306 1423 1316 1426
rect 1298 1403 1301 1416
rect 1313 1413 1316 1423
rect 1290 1203 1293 1226
rect 1298 1203 1301 1326
rect 1290 1106 1293 1196
rect 1298 1123 1301 1196
rect 1290 1103 1297 1106
rect 1294 1036 1297 1103
rect 1290 1033 1297 1036
rect 1290 1013 1293 1033
rect 1306 1016 1309 1396
rect 1314 1383 1317 1406
rect 1314 1146 1317 1366
rect 1322 1306 1325 2136
rect 1330 2103 1333 2126
rect 1338 2113 1341 2136
rect 1330 2013 1333 2036
rect 1338 1993 1341 2076
rect 1346 1953 1349 2216
rect 1354 2213 1357 2243
rect 1362 2193 1365 2206
rect 1354 2123 1357 2136
rect 1362 2086 1365 2136
rect 1370 2123 1373 2236
rect 1378 2213 1381 2243
rect 1394 2226 1397 2353
rect 1390 2223 1397 2226
rect 1390 2156 1393 2223
rect 1390 2153 1397 2156
rect 1362 2083 1373 2086
rect 1354 1996 1357 2066
rect 1362 2013 1365 2036
rect 1370 2013 1373 2083
rect 1378 2073 1381 2136
rect 1386 2053 1389 2136
rect 1386 2006 1389 2016
rect 1370 2003 1389 2006
rect 1354 1993 1373 1996
rect 1354 1936 1357 1946
rect 1330 1823 1333 1926
rect 1338 1893 1341 1936
rect 1346 1933 1357 1936
rect 1338 1813 1341 1836
rect 1330 1793 1333 1806
rect 1330 1693 1333 1726
rect 1330 1603 1333 1616
rect 1330 1543 1333 1566
rect 1338 1553 1341 1736
rect 1346 1703 1349 1916
rect 1354 1883 1357 1926
rect 1362 1803 1365 1966
rect 1370 1913 1373 1993
rect 1378 1903 1381 1996
rect 1370 1813 1373 1896
rect 1378 1846 1381 1876
rect 1386 1853 1389 1996
rect 1378 1843 1389 1846
rect 1370 1796 1373 1806
rect 1378 1803 1381 1836
rect 1386 1813 1389 1843
rect 1354 1733 1357 1796
rect 1370 1793 1381 1796
rect 1354 1713 1357 1726
rect 1370 1703 1373 1786
rect 1378 1696 1381 1793
rect 1386 1713 1389 1796
rect 1362 1693 1381 1696
rect 1346 1613 1349 1626
rect 1346 1546 1349 1586
rect 1338 1543 1349 1546
rect 1338 1533 1341 1543
rect 1354 1533 1357 1666
rect 1362 1623 1365 1693
rect 1330 1413 1333 1526
rect 1362 1516 1365 1616
rect 1370 1563 1373 1636
rect 1378 1596 1381 1626
rect 1386 1603 1389 1626
rect 1378 1593 1389 1596
rect 1370 1543 1373 1556
rect 1378 1533 1381 1546
rect 1386 1533 1389 1593
rect 1354 1513 1365 1516
rect 1354 1426 1357 1513
rect 1370 1473 1373 1526
rect 1354 1423 1361 1426
rect 1338 1403 1341 1416
rect 1346 1403 1349 1416
rect 1330 1323 1333 1336
rect 1338 1323 1341 1346
rect 1346 1306 1349 1376
rect 1322 1303 1329 1306
rect 1326 1216 1329 1303
rect 1322 1213 1329 1216
rect 1338 1303 1349 1306
rect 1322 1193 1325 1213
rect 1338 1166 1341 1303
rect 1358 1296 1361 1423
rect 1354 1293 1361 1296
rect 1346 1213 1349 1226
rect 1338 1163 1349 1166
rect 1314 1143 1341 1146
rect 1330 1096 1333 1116
rect 1322 1093 1333 1096
rect 1322 1036 1325 1093
rect 1322 1033 1333 1036
rect 1302 1013 1309 1016
rect 1330 1013 1333 1033
rect 1266 613 1269 936
rect 1274 933 1277 956
rect 1274 913 1277 926
rect 1282 856 1285 1006
rect 1290 943 1293 1006
rect 1302 936 1305 1013
rect 1298 933 1305 936
rect 1298 883 1301 933
rect 1314 923 1317 996
rect 1322 986 1325 1006
rect 1322 983 1333 986
rect 1322 966 1325 983
rect 1322 963 1329 966
rect 1326 896 1329 963
rect 1322 893 1329 896
rect 1322 876 1325 893
rect 1314 873 1325 876
rect 1282 853 1309 856
rect 1274 803 1277 816
rect 1282 813 1293 816
rect 1298 813 1301 846
rect 1290 746 1293 806
rect 1290 743 1301 746
rect 1306 743 1309 853
rect 1274 713 1277 726
rect 1274 623 1277 686
rect 1282 633 1285 736
rect 1314 673 1317 873
rect 1282 606 1285 626
rect 1278 603 1285 606
rect 1266 533 1269 586
rect 1278 546 1281 603
rect 1278 543 1285 546
rect 1282 526 1285 543
rect 1266 523 1285 526
rect 1266 476 1269 523
rect 1258 473 1269 476
rect 1230 453 1237 456
rect 1226 413 1229 436
rect 1154 393 1161 396
rect 1086 313 1093 316
rect 1122 313 1141 316
rect 1090 293 1093 313
rect 1138 293 1141 306
rect 1074 223 1093 226
rect 1098 213 1101 246
rect 1010 163 1053 166
rect 1010 133 1013 163
rect 1026 133 1029 156
rect 938 116 941 126
rect 914 113 941 116
rect 954 63 957 126
rect 962 113 965 126
rect 1018 103 1021 126
rect 1026 123 1037 126
rect 1034 83 1037 123
rect 1042 93 1045 136
rect 1058 123 1061 196
rect 1090 176 1093 206
rect 1138 196 1141 216
rect 1146 203 1149 386
rect 1158 336 1161 393
rect 1154 333 1161 336
rect 1154 296 1157 333
rect 1162 296 1165 316
rect 1154 293 1165 296
rect 1154 263 1157 293
rect 1154 196 1157 206
rect 1138 193 1157 196
rect 1082 173 1093 176
rect 1106 103 1109 116
rect 1114 113 1117 136
rect 1122 133 1125 186
rect 1138 133 1141 166
rect 1162 133 1165 286
rect 1170 213 1173 406
rect 1194 403 1197 413
rect 1202 383 1205 406
rect 1234 383 1237 453
rect 1242 413 1245 446
rect 1178 306 1181 346
rect 1250 343 1253 406
rect 1258 336 1261 473
rect 1266 396 1269 466
rect 1266 393 1277 396
rect 1274 346 1277 393
rect 1242 333 1261 336
rect 1266 343 1277 346
rect 1242 326 1245 333
rect 1186 323 1245 326
rect 1178 303 1189 306
rect 1186 246 1189 303
rect 1178 243 1189 246
rect 1178 153 1181 243
rect 1186 223 1205 226
rect 1186 206 1189 223
rect 1186 203 1193 206
rect 1190 146 1193 203
rect 1210 193 1213 306
rect 1186 143 1193 146
rect 1162 103 1165 126
rect 1170 73 1173 126
rect 1186 123 1189 143
rect 1202 63 1205 136
rect 1218 133 1221 316
rect 1242 313 1261 316
rect 1242 213 1245 313
rect 1250 293 1253 306
rect 1250 203 1253 226
rect 1242 133 1245 166
rect 1210 103 1213 126
rect 1258 116 1261 216
rect 1266 203 1269 343
rect 1274 213 1277 326
rect 1282 243 1285 306
rect 1282 203 1285 226
rect 1290 183 1293 616
rect 1298 586 1301 666
rect 1306 596 1309 616
rect 1314 613 1317 666
rect 1306 593 1317 596
rect 1298 583 1309 586
rect 1306 506 1309 583
rect 1322 513 1325 816
rect 1330 803 1333 816
rect 1338 773 1341 1143
rect 1346 1133 1349 1163
rect 1346 1113 1349 1126
rect 1346 1073 1349 1106
rect 1346 923 1349 976
rect 1330 613 1333 726
rect 1346 713 1349 916
rect 1354 723 1357 1293
rect 1362 1213 1365 1246
rect 1362 1103 1365 1206
rect 1370 1163 1373 1456
rect 1386 1453 1389 1526
rect 1378 1366 1381 1436
rect 1378 1363 1385 1366
rect 1382 1256 1385 1363
rect 1378 1253 1385 1256
rect 1378 1123 1381 1253
rect 1386 1223 1389 1236
rect 1370 1026 1373 1106
rect 1378 1053 1381 1116
rect 1370 1023 1381 1026
rect 1362 923 1365 996
rect 1370 923 1373 1016
rect 1378 943 1381 1023
rect 1386 1013 1389 1206
rect 1362 746 1365 906
rect 1378 813 1381 846
rect 1370 763 1373 806
rect 1386 803 1389 926
rect 1362 743 1373 746
rect 1362 706 1365 736
rect 1358 703 1365 706
rect 1358 636 1361 703
rect 1370 663 1373 743
rect 1394 736 1397 2153
rect 1402 2106 1405 2216
rect 1410 2133 1413 2216
rect 1418 2203 1421 2236
rect 1426 2213 1429 2306
rect 1442 2263 1445 2426
rect 1466 2403 1469 2473
rect 1498 2466 1501 2516
rect 1506 2476 1509 2736
rect 1514 2726 1517 2743
rect 1514 2723 1525 2726
rect 1522 2636 1525 2723
rect 1538 2713 1541 2726
rect 1554 2673 1557 3006
rect 1562 3003 1565 3133
rect 1594 3093 1597 3126
rect 1602 3123 1613 3126
rect 1618 3106 1621 3146
rect 1642 3143 1661 3146
rect 1610 3103 1621 3106
rect 1578 3023 1581 3036
rect 1562 2886 1565 2936
rect 1570 2903 1573 3016
rect 1586 3013 1597 3016
rect 1602 3013 1605 3026
rect 1594 2996 1597 3006
rect 1610 3003 1613 3103
rect 1618 3076 1621 3103
rect 1626 3083 1629 3126
rect 1634 3116 1637 3136
rect 1634 3113 1645 3116
rect 1618 3073 1629 3076
rect 1618 3013 1621 3066
rect 1626 3036 1629 3073
rect 1642 3066 1645 3113
rect 1634 3063 1645 3066
rect 1634 3043 1637 3063
rect 1658 3046 1661 3143
rect 1674 3123 1677 3216
rect 1682 3213 1685 3233
rect 1826 3233 1845 3236
rect 1690 3203 1693 3216
rect 1698 3193 1709 3196
rect 1682 3103 1685 3126
rect 1658 3043 1669 3046
rect 1626 3033 1637 3036
rect 1618 2996 1621 3006
rect 1626 3003 1629 3016
rect 1634 3006 1637 3033
rect 1642 3013 1645 3036
rect 1634 3003 1653 3006
rect 1594 2993 1621 2996
rect 1658 2993 1661 3016
rect 1666 3003 1669 3043
rect 1602 2933 1605 2946
rect 1610 2933 1621 2936
rect 1610 2916 1613 2926
rect 1626 2923 1629 2956
rect 1658 2933 1661 2966
rect 1674 2926 1677 2956
rect 1682 2936 1685 3086
rect 1706 3043 1709 3126
rect 1706 3013 1709 3036
rect 1714 3003 1717 3136
rect 1722 3113 1725 3126
rect 1730 3123 1733 3166
rect 1754 3133 1757 3216
rect 1770 3213 1773 3226
rect 1786 3213 1797 3216
rect 1818 3213 1821 3226
rect 1762 3193 1765 3206
rect 1794 3193 1797 3213
rect 1826 3203 1829 3233
rect 1778 3143 1781 3156
rect 1786 3133 1789 3166
rect 1818 3143 1829 3146
rect 1834 3136 1837 3216
rect 1842 3183 1845 3226
rect 1850 3213 1853 3266
rect 1826 3133 1837 3136
rect 1826 3126 1829 3133
rect 1722 3013 1725 3096
rect 1738 3013 1741 3106
rect 1722 2946 1725 3006
rect 1746 2956 1749 3046
rect 1754 3023 1757 3036
rect 1754 2963 1757 3006
rect 1746 2953 1757 2956
rect 1706 2943 1725 2946
rect 1682 2933 1701 2936
rect 1706 2933 1709 2943
rect 1586 2913 1613 2916
rect 1634 2903 1637 2926
rect 1562 2883 1573 2886
rect 1570 2836 1573 2883
rect 1666 2866 1669 2926
rect 1674 2923 1685 2926
rect 1562 2833 1573 2836
rect 1658 2863 1669 2866
rect 1562 2813 1565 2833
rect 1658 2823 1661 2863
rect 1698 2846 1701 2933
rect 1714 2863 1717 2926
rect 1698 2843 1709 2846
rect 1610 2793 1613 2816
rect 1618 2803 1621 2816
rect 1642 2803 1645 2816
rect 1658 2766 1661 2806
rect 1518 2633 1525 2636
rect 1518 2576 1521 2633
rect 1530 2603 1533 2616
rect 1546 2603 1549 2616
rect 1570 2613 1573 2736
rect 1586 2733 1589 2766
rect 1634 2763 1661 2766
rect 1674 2763 1677 2806
rect 1706 2796 1709 2843
rect 1722 2813 1725 2936
rect 1730 2933 1733 2946
rect 1738 2813 1741 2936
rect 1754 2913 1757 2953
rect 1762 2896 1765 3066
rect 1770 3003 1773 3026
rect 1778 2983 1781 3126
rect 1802 3123 1829 3126
rect 1826 3093 1829 3123
rect 1850 3116 1853 3126
rect 1858 3123 1861 3246
rect 1874 3193 1877 3216
rect 1866 3116 1869 3136
rect 1850 3113 1869 3116
rect 1874 3096 1877 3126
rect 1882 3116 1885 3226
rect 1914 3216 1917 3226
rect 1922 3223 1925 3236
rect 1898 3213 1917 3216
rect 1898 3146 1901 3213
rect 1946 3206 1949 3236
rect 1906 3203 1949 3206
rect 1922 3183 1925 3196
rect 1930 3146 1933 3176
rect 1954 3153 1957 3226
rect 1970 3223 1981 3226
rect 1986 3223 2037 3226
rect 1978 3216 1981 3223
rect 1970 3186 1973 3216
rect 1978 3213 1997 3216
rect 1994 3193 1997 3213
rect 1962 3183 1973 3186
rect 1970 3163 1973 3183
rect 1898 3143 1933 3146
rect 1914 3133 1925 3136
rect 1930 3133 1933 3143
rect 1986 3133 1989 3146
rect 1994 3133 1997 3186
rect 2002 3163 2005 3216
rect 2034 3186 2037 3223
rect 2042 3216 2045 3226
rect 2050 3223 2077 3226
rect 2042 3213 2053 3216
rect 2042 3193 2045 3206
rect 2050 3203 2053 3213
rect 2034 3183 2045 3186
rect 2026 3133 2029 3166
rect 2034 3133 2037 3156
rect 1930 3123 1965 3126
rect 1930 3116 1933 3123
rect 1882 3113 1933 3116
rect 1858 3093 1877 3096
rect 1786 2963 1789 3016
rect 1810 3013 1813 3036
rect 1818 3003 1821 3056
rect 1858 3053 1861 3093
rect 1882 3086 1885 3106
rect 1866 3083 1885 3086
rect 1850 3033 1861 3036
rect 1858 3023 1861 3033
rect 1826 3003 1829 3016
rect 1834 2983 1837 3006
rect 1842 2993 1845 3016
rect 1858 2976 1861 3006
rect 1866 3003 1869 3083
rect 1874 3013 1877 3066
rect 1898 3013 1909 3016
rect 1906 2986 1909 3013
rect 1914 2996 1917 3016
rect 1922 3003 1925 3056
rect 1938 3016 1941 3026
rect 1954 3023 1957 3036
rect 1962 3023 1965 3096
rect 1930 3013 1941 3016
rect 1946 3013 1973 3016
rect 1946 3003 1949 3013
rect 1914 2993 1965 2996
rect 1906 2983 1917 2986
rect 1802 2973 1861 2976
rect 1778 2933 1789 2936
rect 1802 2933 1805 2973
rect 1818 2933 1821 2966
rect 1754 2893 1765 2896
rect 1698 2793 1709 2796
rect 1634 2723 1637 2763
rect 1514 2573 1521 2576
rect 1514 2523 1517 2573
rect 1554 2503 1557 2536
rect 1586 2533 1589 2566
rect 1570 2523 1581 2526
rect 1594 2523 1597 2606
rect 1570 2486 1573 2523
rect 1602 2516 1605 2526
rect 1562 2483 1573 2486
rect 1586 2513 1605 2516
rect 1506 2473 1517 2476
rect 1482 2463 1501 2466
rect 1458 2333 1461 2346
rect 1466 2333 1469 2396
rect 1482 2393 1485 2463
rect 1458 2303 1461 2316
rect 1442 2226 1445 2236
rect 1442 2223 1453 2226
rect 1434 2213 1445 2216
rect 1450 2213 1453 2223
rect 1426 2203 1437 2206
rect 1426 2123 1429 2146
rect 1402 2103 1413 2106
rect 1410 2026 1413 2103
rect 1434 2076 1437 2156
rect 1442 2146 1445 2206
rect 1474 2146 1477 2366
rect 1490 2323 1493 2346
rect 1506 2333 1509 2416
rect 1514 2363 1517 2473
rect 1562 2426 1565 2483
rect 1586 2466 1589 2513
rect 1610 2503 1613 2536
rect 1634 2533 1637 2556
rect 1554 2423 1565 2426
rect 1578 2463 1589 2466
rect 1554 2406 1557 2423
rect 1550 2403 1557 2406
rect 1538 2333 1541 2346
rect 1550 2316 1553 2403
rect 1514 2286 1517 2306
rect 1442 2143 1461 2146
rect 1474 2143 1485 2146
rect 1402 2023 1413 2026
rect 1426 2073 1437 2076
rect 1426 2026 1429 2073
rect 1442 2026 1445 2066
rect 1450 2033 1453 2136
rect 1458 2123 1461 2143
rect 1466 2073 1469 2136
rect 1474 2113 1477 2136
rect 1482 2056 1485 2143
rect 1458 2053 1485 2056
rect 1426 2023 1437 2026
rect 1442 2023 1453 2026
rect 1402 1963 1405 2023
rect 1402 1713 1405 1956
rect 1418 1926 1421 1996
rect 1426 1953 1429 2006
rect 1434 1963 1437 2023
rect 1450 2006 1453 2023
rect 1446 2003 1453 2006
rect 1446 1946 1449 2003
rect 1410 1923 1421 1926
rect 1434 1943 1449 1946
rect 1434 1923 1437 1943
rect 1410 1803 1413 1923
rect 1418 1913 1429 1916
rect 1434 1896 1437 1916
rect 1430 1893 1437 1896
rect 1442 1893 1445 1926
rect 1430 1826 1433 1893
rect 1418 1733 1421 1826
rect 1426 1823 1433 1826
rect 1402 1703 1421 1706
rect 1402 1503 1405 1616
rect 1410 1533 1413 1696
rect 1410 1476 1413 1516
rect 1406 1473 1413 1476
rect 1406 1396 1409 1473
rect 1418 1443 1421 1703
rect 1426 1603 1429 1823
rect 1434 1803 1437 1816
rect 1442 1736 1445 1856
rect 1450 1823 1453 1936
rect 1458 1853 1461 2053
rect 1474 2013 1477 2036
rect 1482 2013 1485 2046
rect 1466 1993 1469 2006
rect 1466 1913 1469 1926
rect 1474 1883 1477 2006
rect 1482 1876 1485 1926
rect 1466 1873 1485 1876
rect 1450 1793 1453 1816
rect 1458 1783 1461 1816
rect 1466 1793 1469 1873
rect 1474 1803 1477 1816
rect 1482 1803 1485 1836
rect 1490 1826 1493 2226
rect 1498 1903 1501 2286
rect 1510 2283 1517 2286
rect 1510 2216 1513 2283
rect 1510 2213 1517 2216
rect 1506 2163 1509 2196
rect 1506 2133 1509 2156
rect 1514 2123 1517 2213
rect 1506 2066 1509 2086
rect 1506 2063 1513 2066
rect 1510 1996 1513 2063
rect 1506 1993 1513 1996
rect 1506 1903 1509 1993
rect 1498 1833 1501 1896
rect 1490 1823 1501 1826
rect 1490 1803 1493 1816
rect 1498 1786 1501 1823
rect 1494 1783 1501 1786
rect 1442 1733 1461 1736
rect 1434 1693 1437 1716
rect 1442 1703 1445 1726
rect 1434 1636 1437 1656
rect 1434 1633 1441 1636
rect 1426 1533 1429 1556
rect 1426 1436 1429 1526
rect 1438 1506 1441 1633
rect 1450 1603 1453 1716
rect 1458 1653 1461 1733
rect 1466 1683 1469 1706
rect 1458 1606 1461 1646
rect 1466 1623 1469 1666
rect 1474 1613 1477 1766
rect 1494 1726 1497 1783
rect 1506 1733 1509 1896
rect 1514 1813 1517 1976
rect 1482 1643 1485 1726
rect 1490 1723 1497 1726
rect 1490 1696 1493 1723
rect 1498 1703 1501 1716
rect 1490 1693 1501 1696
rect 1490 1613 1493 1686
rect 1498 1626 1501 1693
rect 1514 1653 1517 1806
rect 1514 1633 1517 1646
rect 1498 1623 1509 1626
rect 1506 1613 1509 1623
rect 1458 1603 1465 1606
rect 1450 1523 1453 1556
rect 1462 1516 1465 1603
rect 1482 1583 1485 1606
rect 1474 1533 1477 1576
rect 1506 1523 1509 1536
rect 1458 1513 1465 1516
rect 1438 1503 1445 1506
rect 1442 1436 1445 1503
rect 1458 1443 1461 1513
rect 1482 1493 1485 1516
rect 1490 1483 1493 1506
rect 1506 1496 1509 1516
rect 1502 1493 1509 1496
rect 1418 1433 1429 1436
rect 1434 1433 1445 1436
rect 1418 1396 1421 1433
rect 1426 1403 1429 1426
rect 1406 1393 1413 1396
rect 1418 1393 1429 1396
rect 1402 1323 1405 1336
rect 1402 1203 1405 1266
rect 1402 1063 1405 1136
rect 1410 1133 1413 1393
rect 1410 1013 1413 1126
rect 1418 1023 1421 1386
rect 1426 1236 1429 1393
rect 1434 1253 1437 1433
rect 1458 1423 1469 1426
rect 1442 1403 1445 1416
rect 1450 1413 1461 1416
rect 1466 1413 1469 1423
rect 1458 1386 1461 1406
rect 1450 1383 1461 1386
rect 1466 1383 1469 1406
rect 1482 1403 1485 1456
rect 1442 1333 1445 1346
rect 1442 1236 1445 1286
rect 1450 1253 1453 1383
rect 1426 1233 1437 1236
rect 1442 1233 1449 1236
rect 1426 1213 1429 1226
rect 1426 1083 1429 1126
rect 1434 1093 1437 1233
rect 1446 1146 1449 1233
rect 1446 1143 1453 1146
rect 1442 1123 1445 1136
rect 1450 1076 1453 1143
rect 1458 1106 1461 1256
rect 1466 1213 1469 1336
rect 1474 1333 1485 1336
rect 1490 1326 1493 1416
rect 1502 1346 1505 1493
rect 1514 1483 1517 1626
rect 1522 1496 1525 2316
rect 1550 2313 1557 2316
rect 1530 2213 1533 2276
rect 1530 2143 1533 2206
rect 1538 2153 1541 2196
rect 1530 2036 1533 2126
rect 1538 2103 1541 2136
rect 1546 2123 1549 2296
rect 1554 2186 1557 2313
rect 1562 2303 1565 2376
rect 1570 2333 1573 2416
rect 1578 2413 1581 2463
rect 1594 2393 1597 2406
rect 1594 2356 1597 2376
rect 1626 2363 1629 2526
rect 1642 2523 1645 2616
rect 1658 2603 1661 2616
rect 1682 2613 1685 2696
rect 1698 2603 1701 2793
rect 1722 2743 1725 2806
rect 1754 2746 1757 2893
rect 1770 2746 1773 2926
rect 1778 2923 1789 2926
rect 1778 2913 1781 2923
rect 1810 2916 1813 2926
rect 1826 2923 1829 2956
rect 1786 2913 1813 2916
rect 1850 2826 1853 2936
rect 1866 2903 1869 2966
rect 1898 2933 1901 2946
rect 1914 2933 1917 2983
rect 1922 2933 1925 2986
rect 1834 2823 1853 2826
rect 1906 2826 1909 2926
rect 1930 2923 1933 2976
rect 1938 2923 1941 2956
rect 1954 2933 1957 2946
rect 1962 2913 1965 2993
rect 1978 2983 1981 3116
rect 2018 3113 2021 3126
rect 2042 3123 2045 3183
rect 2058 3153 2061 3216
rect 2074 3213 2077 3223
rect 2082 3203 2085 3236
rect 2090 3213 2093 3246
rect 2106 3203 2109 3226
rect 2178 3223 2181 3246
rect 2114 3173 2117 3206
rect 2122 3183 2125 3216
rect 2130 3193 2133 3206
rect 2138 3203 2141 3216
rect 2170 3213 2181 3216
rect 2178 3193 2181 3206
rect 2186 3203 2189 3236
rect 2258 3213 2261 3236
rect 2202 3203 2213 3206
rect 2218 3186 2221 3206
rect 2266 3203 2269 3216
rect 2322 3213 2325 3226
rect 2330 3213 2333 3246
rect 2282 3193 2285 3206
rect 2322 3193 2325 3206
rect 2210 3183 2221 3186
rect 2058 3143 2117 3146
rect 2058 3123 2061 3143
rect 2066 3133 2077 3136
rect 2082 3133 2085 3143
rect 2090 3133 2109 3136
rect 2074 3126 2077 3133
rect 2090 3126 2093 3133
rect 2066 3113 2069 3126
rect 2074 3123 2093 3126
rect 2098 3106 2101 3126
rect 2094 3103 2101 3106
rect 1906 2823 1917 2826
rect 1802 2763 1805 2806
rect 1754 2743 1765 2746
rect 1770 2743 1805 2746
rect 1730 2693 1733 2736
rect 1738 2713 1741 2726
rect 1762 2723 1765 2743
rect 1722 2613 1741 2616
rect 1666 2503 1669 2536
rect 1682 2533 1709 2536
rect 1714 2533 1717 2566
rect 1682 2486 1685 2533
rect 1674 2483 1685 2486
rect 1594 2353 1601 2356
rect 1578 2323 1581 2336
rect 1586 2306 1589 2336
rect 1578 2303 1589 2306
rect 1562 2213 1565 2276
rect 1578 2236 1581 2303
rect 1598 2296 1601 2353
rect 1610 2333 1613 2346
rect 1642 2343 1645 2416
rect 1674 2386 1677 2483
rect 1690 2413 1693 2526
rect 1706 2516 1709 2533
rect 1722 2523 1725 2613
rect 1730 2516 1733 2536
rect 1738 2523 1741 2606
rect 1754 2603 1757 2616
rect 1786 2606 1789 2736
rect 1802 2613 1805 2686
rect 1786 2603 1797 2606
rect 1794 2546 1797 2603
rect 1834 2586 1837 2823
rect 1850 2803 1853 2816
rect 1866 2813 1885 2816
rect 1842 2723 1845 2736
rect 1858 2656 1861 2736
rect 1866 2733 1869 2813
rect 1890 2803 1893 2816
rect 1898 2746 1901 2816
rect 1906 2803 1917 2806
rect 1946 2763 1949 2846
rect 1970 2776 1973 2926
rect 1978 2916 1981 2936
rect 1978 2913 1985 2916
rect 1982 2836 1985 2913
rect 1978 2833 1985 2836
rect 1978 2813 1981 2833
rect 1986 2803 1989 2816
rect 1954 2773 1973 2776
rect 1882 2743 1901 2746
rect 1954 2743 1957 2773
rect 1890 2683 1893 2736
rect 1898 2713 1901 2726
rect 1962 2656 1965 2736
rect 1978 2733 1981 2786
rect 1970 2713 1973 2726
rect 1994 2656 1997 3036
rect 2002 3023 2037 3026
rect 2002 3013 2005 3023
rect 2010 2963 2013 3016
rect 2018 2983 2021 3006
rect 2002 2933 2005 2946
rect 2010 2933 2021 2936
rect 2026 2916 2029 3016
rect 2034 3003 2037 3023
rect 2042 2973 2045 3046
rect 2066 3003 2069 3016
rect 2082 3003 2085 3096
rect 2094 3036 2097 3103
rect 2106 3053 2109 3133
rect 2094 3033 2101 3036
rect 2090 2956 2093 3016
rect 2098 3003 2101 3033
rect 2090 2953 2097 2956
rect 2002 2913 2029 2916
rect 2034 2913 2037 2926
rect 2058 2843 2061 2936
rect 2082 2923 2085 2946
rect 2094 2896 2097 2953
rect 2106 2913 2109 3046
rect 2114 3006 2117 3143
rect 2122 3093 2125 3136
rect 2130 3133 2133 3146
rect 2178 3133 2181 3166
rect 2210 3163 2213 3183
rect 2218 3173 2229 3176
rect 2338 3173 2341 3226
rect 2154 3123 2165 3126
rect 2170 3116 2173 3126
rect 2146 3113 2173 3116
rect 2122 3013 2125 3036
rect 2114 3003 2125 3006
rect 2090 2893 2097 2896
rect 2090 2876 2093 2893
rect 2066 2873 2093 2876
rect 2058 2816 2061 2836
rect 2066 2823 2069 2873
rect 2130 2846 2133 3056
rect 2146 2983 2149 3006
rect 2154 3003 2157 3026
rect 2162 3023 2173 3026
rect 2178 3016 2181 3036
rect 2170 3013 2181 3016
rect 2186 3013 2189 3056
rect 2170 2963 2173 3013
rect 2194 2983 2197 2996
rect 2138 2923 2141 2936
rect 2026 2783 2029 2816
rect 2034 2746 2037 2816
rect 2042 2803 2045 2816
rect 2050 2813 2069 2816
rect 2026 2743 2037 2746
rect 2050 2743 2053 2813
rect 2058 2803 2069 2806
rect 2074 2803 2077 2826
rect 2114 2803 2117 2846
rect 2130 2843 2141 2846
rect 2138 2826 2141 2843
rect 2146 2833 2149 2926
rect 2138 2823 2149 2826
rect 2146 2776 2149 2823
rect 2154 2813 2157 2936
rect 2178 2926 2181 2936
rect 2170 2923 2181 2926
rect 2170 2856 2173 2923
rect 2178 2903 2181 2916
rect 2162 2853 2173 2856
rect 2162 2813 2165 2853
rect 2186 2846 2189 2936
rect 2202 2893 2205 3116
rect 2210 3113 2213 3126
rect 2226 3113 2229 3173
rect 2234 3133 2237 3146
rect 2274 3133 2277 3166
rect 2330 3156 2333 3166
rect 2330 3153 2349 3156
rect 2282 3133 2285 3146
rect 2218 3003 2221 3106
rect 2250 3103 2253 3126
rect 2210 2923 2213 2976
rect 2218 2933 2221 2956
rect 2226 2933 2229 3096
rect 2266 3056 2269 3126
rect 2282 3113 2285 3126
rect 2306 3123 2309 3136
rect 2330 3133 2333 3153
rect 2322 3106 2325 3126
rect 2314 3103 2325 3106
rect 2258 3053 2269 3056
rect 2234 3013 2237 3036
rect 2258 3023 2261 3053
rect 2274 3026 2277 3076
rect 2314 3046 2317 3103
rect 2314 3043 2325 3046
rect 2270 3023 2277 3026
rect 2322 3023 2325 3043
rect 2250 3013 2261 3016
rect 2250 3006 2253 3013
rect 2234 3003 2253 3006
rect 2234 2933 2237 2946
rect 2226 2903 2229 2926
rect 2242 2896 2245 2966
rect 2258 2956 2261 3006
rect 2270 2966 2273 3023
rect 2270 2963 2277 2966
rect 2250 2953 2261 2956
rect 2250 2913 2253 2926
rect 2274 2923 2277 2963
rect 2282 2933 2285 3016
rect 2290 3013 2309 3016
rect 2330 3013 2333 3036
rect 2290 2993 2293 3013
rect 2298 3003 2325 3006
rect 2338 3003 2341 3146
rect 2346 3043 2349 3153
rect 2354 3146 2357 3216
rect 2362 3153 2365 3206
rect 2370 3193 2373 3216
rect 2378 3176 2381 3206
rect 2410 3186 2413 3216
rect 2426 3203 2429 3236
rect 2506 3233 2533 3236
rect 2434 3193 2437 3226
rect 2442 3223 2469 3226
rect 2442 3203 2445 3223
rect 2410 3183 2429 3186
rect 2370 3173 2381 3176
rect 2354 3143 2365 3146
rect 2346 3013 2349 3026
rect 2242 2893 2253 2896
rect 2290 2893 2293 2976
rect 2298 2933 2301 3003
rect 2322 2936 2325 2996
rect 2354 2953 2357 3136
rect 2362 3063 2365 3143
rect 2370 3123 2373 3173
rect 2394 3133 2413 3136
rect 2378 3113 2381 3126
rect 2386 3103 2389 3126
rect 2394 3103 2397 3133
rect 2410 3106 2413 3116
rect 2418 3113 2421 3176
rect 2426 3106 2429 3183
rect 2442 3153 2453 3156
rect 2410 3103 2429 3106
rect 2370 3003 2373 3046
rect 2378 2976 2381 3086
rect 2386 3076 2389 3096
rect 2386 3073 2397 3076
rect 2370 2973 2381 2976
rect 2306 2933 2317 2936
rect 2322 2933 2333 2936
rect 2182 2843 2189 2846
rect 2182 2776 2185 2843
rect 2194 2813 2197 2826
rect 2234 2823 2237 2856
rect 2250 2836 2253 2893
rect 2306 2853 2309 2926
rect 2322 2883 2325 2926
rect 2330 2856 2333 2933
rect 2338 2923 2341 2936
rect 2354 2913 2357 2926
rect 2322 2853 2333 2856
rect 2250 2833 2261 2836
rect 2210 2803 2213 2816
rect 2218 2813 2237 2816
rect 2146 2773 2153 2776
rect 2098 2763 2141 2766
rect 2042 2726 2045 2736
rect 2050 2733 2093 2736
rect 2098 2733 2101 2763
rect 2042 2723 2069 2726
rect 1858 2653 1885 2656
rect 1962 2653 1989 2656
rect 1994 2653 2029 2656
rect 1826 2583 1837 2586
rect 1794 2543 1805 2546
rect 1706 2513 1733 2516
rect 1746 2503 1749 2536
rect 1706 2393 1709 2436
rect 1674 2383 1685 2386
rect 1658 2333 1669 2336
rect 1674 2333 1677 2356
rect 1682 2326 1685 2383
rect 1746 2366 1749 2386
rect 1754 2373 1757 2416
rect 1786 2413 1789 2526
rect 1802 2436 1805 2543
rect 1810 2533 1813 2556
rect 1826 2536 1829 2583
rect 1842 2543 1845 2616
rect 1858 2603 1861 2616
rect 1882 2613 1885 2653
rect 1826 2533 1837 2536
rect 1834 2446 1837 2533
rect 1858 2523 1869 2526
rect 1834 2443 1841 2446
rect 1794 2433 1805 2436
rect 1770 2376 1773 2396
rect 1762 2373 1773 2376
rect 1746 2363 1757 2366
rect 1698 2333 1701 2346
rect 1594 2293 1601 2296
rect 1578 2233 1589 2236
rect 1554 2183 1565 2186
rect 1554 2043 1557 2176
rect 1530 2033 1541 2036
rect 1530 2003 1533 2026
rect 1530 1933 1533 1946
rect 1538 1896 1541 2033
rect 1546 2013 1549 2036
rect 1562 2026 1565 2183
rect 1570 2123 1573 2136
rect 1578 2133 1581 2216
rect 1586 2206 1589 2233
rect 1594 2213 1597 2293
rect 1586 2203 1597 2206
rect 1602 2203 1605 2226
rect 1618 2216 1621 2306
rect 1634 2263 1637 2326
rect 1642 2323 1685 2326
rect 1738 2323 1741 2346
rect 1754 2333 1757 2363
rect 1762 2323 1765 2373
rect 1778 2323 1781 2336
rect 1786 2333 1789 2356
rect 1794 2323 1797 2433
rect 1810 2403 1813 2416
rect 1838 2376 1841 2443
rect 1826 2333 1829 2376
rect 1834 2373 1841 2376
rect 1834 2326 1837 2373
rect 1842 2333 1845 2356
rect 1610 2213 1621 2216
rect 1626 2213 1629 2236
rect 1634 2213 1637 2226
rect 1586 2133 1589 2156
rect 1594 2123 1597 2203
rect 1602 2056 1605 2136
rect 1610 2126 1613 2196
rect 1618 2163 1621 2206
rect 1626 2143 1629 2206
rect 1634 2133 1637 2146
rect 1610 2123 1621 2126
rect 1618 2056 1621 2123
rect 1578 2053 1605 2056
rect 1610 2053 1621 2056
rect 1558 2023 1565 2026
rect 1558 1956 1561 2023
rect 1570 2013 1573 2026
rect 1578 2006 1581 2053
rect 1570 2003 1581 2006
rect 1594 1996 1597 2016
rect 1602 2013 1605 2026
rect 1558 1953 1565 1956
rect 1546 1933 1557 1936
rect 1546 1913 1549 1933
rect 1538 1893 1545 1896
rect 1530 1803 1533 1886
rect 1542 1826 1545 1893
rect 1554 1883 1557 1926
rect 1562 1896 1565 1953
rect 1570 1913 1573 1996
rect 1578 1993 1597 1996
rect 1602 1993 1605 2006
rect 1578 1923 1581 1993
rect 1610 1986 1613 2053
rect 1626 2013 1629 2036
rect 1618 2003 1629 2006
rect 1634 2003 1637 2106
rect 1610 1983 1617 1986
rect 1562 1893 1569 1896
rect 1538 1823 1545 1826
rect 1554 1823 1557 1846
rect 1566 1826 1569 1893
rect 1562 1823 1569 1826
rect 1530 1723 1533 1736
rect 1530 1696 1533 1716
rect 1538 1713 1541 1823
rect 1546 1783 1549 1806
rect 1530 1693 1537 1696
rect 1534 1616 1537 1693
rect 1534 1613 1541 1616
rect 1546 1613 1549 1716
rect 1530 1513 1533 1606
rect 1538 1573 1541 1613
rect 1554 1593 1557 1806
rect 1522 1493 1529 1496
rect 1514 1373 1517 1466
rect 1526 1426 1529 1493
rect 1522 1423 1529 1426
rect 1502 1343 1509 1346
rect 1474 1323 1493 1326
rect 1474 1303 1477 1323
rect 1498 1306 1501 1326
rect 1490 1303 1501 1306
rect 1474 1216 1477 1256
rect 1490 1236 1493 1303
rect 1490 1233 1501 1236
rect 1498 1216 1501 1233
rect 1474 1213 1501 1216
rect 1466 1173 1469 1206
rect 1482 1146 1485 1196
rect 1490 1153 1493 1206
rect 1498 1146 1501 1206
rect 1482 1143 1501 1146
rect 1466 1123 1469 1136
rect 1458 1103 1465 1106
rect 1434 1073 1453 1076
rect 1434 1013 1437 1073
rect 1434 956 1437 1006
rect 1442 1003 1445 1066
rect 1462 1036 1465 1103
rect 1458 1033 1465 1036
rect 1450 1013 1453 1026
rect 1434 953 1441 956
rect 1402 753 1405 916
rect 1418 913 1421 926
rect 1410 853 1413 906
rect 1410 776 1413 836
rect 1426 786 1429 946
rect 1438 906 1441 953
rect 1450 923 1453 1006
rect 1438 903 1445 906
rect 1442 846 1445 903
rect 1442 843 1453 846
rect 1450 803 1453 843
rect 1458 796 1461 1033
rect 1466 963 1469 1016
rect 1474 1013 1477 1026
rect 1482 1003 1485 1126
rect 1490 1003 1493 1086
rect 1498 973 1501 1106
rect 1506 1096 1509 1343
rect 1514 1313 1517 1336
rect 1522 1296 1525 1423
rect 1538 1413 1541 1426
rect 1518 1293 1525 1296
rect 1518 1216 1521 1293
rect 1518 1213 1525 1216
rect 1514 1113 1517 1196
rect 1506 1093 1513 1096
rect 1510 1026 1513 1093
rect 1506 1023 1513 1026
rect 1474 933 1477 946
rect 1482 926 1485 966
rect 1506 926 1509 1023
rect 1514 943 1517 1006
rect 1466 913 1469 926
rect 1474 923 1485 926
rect 1474 813 1477 923
rect 1498 913 1501 926
rect 1506 923 1513 926
rect 1482 823 1493 826
rect 1482 796 1485 823
rect 1490 803 1493 816
rect 1498 803 1501 896
rect 1510 846 1513 923
rect 1506 843 1513 846
rect 1450 793 1461 796
rect 1474 793 1485 796
rect 1426 783 1437 786
rect 1410 773 1421 776
rect 1394 733 1413 736
rect 1418 733 1421 773
rect 1410 726 1413 733
rect 1378 723 1397 726
rect 1410 723 1421 726
rect 1358 633 1365 636
rect 1338 623 1349 626
rect 1346 616 1349 623
rect 1338 603 1341 616
rect 1346 613 1357 616
rect 1306 503 1317 506
rect 1298 403 1301 456
rect 1314 393 1317 503
rect 1330 393 1333 576
rect 1338 503 1341 536
rect 1362 426 1365 633
rect 1370 613 1373 626
rect 1370 573 1373 606
rect 1378 533 1381 723
rect 1386 673 1389 716
rect 1394 713 1413 716
rect 1394 703 1397 713
rect 1402 703 1413 706
rect 1418 696 1421 723
rect 1434 696 1437 783
rect 1450 723 1453 793
rect 1466 723 1469 736
rect 1394 693 1421 696
rect 1426 693 1437 696
rect 1466 693 1469 716
rect 1386 603 1389 646
rect 1394 583 1397 693
rect 1426 673 1429 693
rect 1474 676 1477 793
rect 1482 743 1485 786
rect 1466 673 1477 676
rect 1402 623 1437 626
rect 1378 443 1381 526
rect 1386 463 1389 526
rect 1402 523 1405 623
rect 1418 573 1421 616
rect 1426 536 1429 606
rect 1434 596 1437 606
rect 1442 603 1445 626
rect 1450 596 1453 646
rect 1434 593 1453 596
rect 1466 546 1469 673
rect 1482 656 1485 726
rect 1498 703 1501 736
rect 1478 653 1485 656
rect 1478 586 1481 653
rect 1490 593 1493 676
rect 1498 613 1501 626
rect 1478 583 1485 586
rect 1466 543 1477 546
rect 1410 513 1413 536
rect 1422 533 1429 536
rect 1362 423 1397 426
rect 1362 413 1365 423
rect 1298 253 1301 336
rect 1306 316 1309 346
rect 1314 323 1317 336
rect 1306 313 1317 316
rect 1306 203 1309 216
rect 1258 113 1269 116
rect 1290 103 1293 136
rect 1298 133 1301 146
rect 1314 133 1317 313
rect 1330 223 1333 356
rect 1354 323 1357 406
rect 1362 243 1365 386
rect 1370 353 1373 406
rect 1378 373 1381 416
rect 1386 236 1389 416
rect 1394 333 1397 423
rect 1410 416 1413 476
rect 1422 466 1425 533
rect 1422 463 1429 466
rect 1402 413 1413 416
rect 1402 383 1405 406
rect 1418 396 1421 446
rect 1414 393 1421 396
rect 1322 173 1325 206
rect 1330 116 1333 216
rect 1338 203 1341 216
rect 1346 213 1349 236
rect 1386 233 1397 236
rect 1402 233 1405 326
rect 1414 296 1417 393
rect 1426 333 1429 463
rect 1434 456 1437 526
rect 1442 513 1445 536
rect 1450 523 1453 536
rect 1434 453 1453 456
rect 1434 403 1437 416
rect 1442 413 1445 446
rect 1450 386 1453 453
rect 1442 383 1453 386
rect 1442 326 1445 383
rect 1430 323 1445 326
rect 1414 293 1421 296
rect 1354 193 1357 226
rect 1394 213 1397 233
rect 1410 203 1413 226
rect 1418 203 1421 293
rect 1430 216 1433 323
rect 1458 316 1461 476
rect 1466 443 1469 526
rect 1466 333 1469 426
rect 1442 293 1445 316
rect 1450 313 1461 316
rect 1426 213 1433 216
rect 1426 196 1429 213
rect 1418 193 1429 196
rect 1330 113 1365 116
rect 1370 83 1373 146
rect 1394 133 1397 146
rect 1402 133 1405 166
rect 1418 126 1421 193
rect 1442 146 1445 216
rect 1450 193 1453 313
rect 1474 296 1477 543
rect 1482 533 1485 583
rect 1482 503 1485 526
rect 1498 503 1501 606
rect 1506 436 1509 843
rect 1514 803 1517 826
rect 1514 723 1517 776
rect 1522 683 1525 1213
rect 1530 1193 1533 1406
rect 1530 1083 1533 1106
rect 1530 1013 1533 1066
rect 1538 1026 1541 1336
rect 1546 1043 1549 1546
rect 1562 1443 1565 1823
rect 1570 1793 1573 1806
rect 1578 1783 1581 1816
rect 1570 1703 1573 1726
rect 1578 1633 1581 1736
rect 1570 1583 1573 1626
rect 1578 1523 1581 1606
rect 1570 1493 1581 1496
rect 1554 1423 1557 1436
rect 1562 1413 1565 1426
rect 1554 1393 1557 1406
rect 1562 1403 1573 1406
rect 1578 1403 1581 1493
rect 1554 1326 1557 1386
rect 1562 1333 1565 1376
rect 1570 1363 1573 1403
rect 1586 1373 1589 1906
rect 1594 1893 1597 1916
rect 1594 1743 1597 1816
rect 1602 1813 1605 1966
rect 1614 1856 1617 1983
rect 1626 1916 1629 1926
rect 1634 1923 1637 1966
rect 1626 1913 1637 1916
rect 1610 1853 1617 1856
rect 1602 1753 1605 1806
rect 1610 1733 1613 1853
rect 1618 1823 1621 1836
rect 1602 1656 1605 1726
rect 1610 1713 1613 1726
rect 1594 1653 1605 1656
rect 1594 1613 1597 1653
rect 1618 1643 1621 1816
rect 1626 1813 1629 1866
rect 1594 1543 1597 1606
rect 1610 1603 1613 1616
rect 1626 1613 1629 1766
rect 1634 1663 1637 1913
rect 1554 1323 1565 1326
rect 1570 1323 1581 1326
rect 1554 1133 1557 1306
rect 1554 1113 1557 1126
rect 1538 1023 1545 1026
rect 1530 833 1533 1006
rect 1542 956 1545 1023
rect 1538 953 1545 956
rect 1538 866 1541 953
rect 1554 946 1557 1086
rect 1562 963 1565 1323
rect 1570 1203 1573 1226
rect 1570 1133 1573 1146
rect 1570 1083 1573 1126
rect 1554 943 1561 946
rect 1546 883 1549 936
rect 1558 876 1561 943
rect 1554 873 1561 876
rect 1538 863 1545 866
rect 1542 806 1545 863
rect 1554 813 1557 873
rect 1570 813 1573 1006
rect 1542 803 1557 806
rect 1562 803 1573 806
rect 1530 733 1533 786
rect 1546 736 1549 756
rect 1542 733 1549 736
rect 1530 673 1533 726
rect 1542 626 1545 733
rect 1514 533 1517 626
rect 1530 613 1533 626
rect 1542 623 1549 626
rect 1546 606 1549 623
rect 1522 603 1549 606
rect 1554 596 1557 803
rect 1578 786 1581 1316
rect 1586 1303 1589 1336
rect 1586 1223 1589 1246
rect 1586 1163 1589 1216
rect 1594 1123 1597 1516
rect 1602 1473 1605 1526
rect 1618 1513 1621 1606
rect 1634 1603 1637 1636
rect 1626 1533 1629 1566
rect 1634 1496 1637 1576
rect 1626 1493 1637 1496
rect 1602 1383 1605 1446
rect 1626 1416 1629 1493
rect 1626 1413 1637 1416
rect 1626 1346 1629 1396
rect 1602 1323 1605 1346
rect 1622 1343 1629 1346
rect 1610 1316 1613 1336
rect 1602 1313 1613 1316
rect 1602 1203 1605 1313
rect 1610 1146 1613 1276
rect 1622 1266 1625 1343
rect 1634 1283 1637 1413
rect 1622 1263 1629 1266
rect 1618 1213 1621 1246
rect 1610 1143 1617 1146
rect 1586 1113 1597 1116
rect 1586 1053 1589 1113
rect 1586 833 1589 1046
rect 1562 783 1581 786
rect 1562 716 1565 783
rect 1570 723 1573 776
rect 1586 753 1589 806
rect 1594 746 1597 1086
rect 1602 1003 1605 1136
rect 1614 1056 1617 1143
rect 1626 1123 1629 1263
rect 1634 1213 1637 1276
rect 1614 1053 1629 1056
rect 1610 1003 1613 1016
rect 1618 983 1621 1006
rect 1610 943 1613 966
rect 1626 943 1629 1053
rect 1634 936 1637 1206
rect 1582 743 1597 746
rect 1602 743 1605 936
rect 1610 773 1613 926
rect 1618 783 1621 936
rect 1626 933 1637 936
rect 1626 853 1629 933
rect 1634 913 1637 926
rect 1626 826 1629 846
rect 1626 823 1633 826
rect 1630 776 1633 823
rect 1642 813 1645 2323
rect 1698 2296 1701 2316
rect 1810 2306 1813 2326
rect 1834 2323 1845 2326
rect 1850 2316 1853 2476
rect 1874 2433 1877 2536
rect 1882 2466 1885 2526
rect 1890 2503 1893 2536
rect 1898 2523 1901 2606
rect 1906 2533 1909 2566
rect 1946 2533 1949 2616
rect 1962 2603 1965 2616
rect 1986 2613 1989 2653
rect 1986 2543 2005 2546
rect 1962 2533 1973 2536
rect 1914 2523 1925 2526
rect 1962 2483 1965 2533
rect 1970 2523 1981 2526
rect 1882 2463 1893 2466
rect 1858 2346 1861 2416
rect 1890 2413 1893 2463
rect 1906 2403 1909 2416
rect 1954 2376 1957 2416
rect 1986 2413 1989 2543
rect 1994 2496 1997 2536
rect 2002 2523 2005 2543
rect 2018 2503 2021 2536
rect 1994 2493 2005 2496
rect 2002 2403 2005 2493
rect 2026 2446 2029 2653
rect 2034 2533 2037 2586
rect 2042 2533 2045 2616
rect 2066 2603 2069 2616
rect 2090 2613 2093 2733
rect 2114 2613 2117 2736
rect 2138 2723 2141 2763
rect 2150 2716 2153 2773
rect 2146 2713 2153 2716
rect 2162 2773 2185 2776
rect 2146 2696 2149 2713
rect 2138 2693 2149 2696
rect 2138 2636 2141 2693
rect 2130 2633 2141 2636
rect 2050 2493 2053 2536
rect 2114 2533 2117 2556
rect 2130 2526 2133 2633
rect 2162 2626 2165 2773
rect 2218 2743 2221 2813
rect 2250 2806 2253 2826
rect 2226 2803 2237 2806
rect 2242 2803 2253 2806
rect 2258 2766 2261 2833
rect 2282 2803 2285 2846
rect 2306 2803 2309 2816
rect 2322 2776 2325 2853
rect 2370 2826 2373 2973
rect 2394 2966 2397 3073
rect 2410 3013 2413 3036
rect 2418 3013 2421 3103
rect 2426 3013 2429 3026
rect 2434 3006 2437 3146
rect 2450 3133 2453 3153
rect 2458 3143 2461 3216
rect 2466 3166 2469 3223
rect 2474 3186 2477 3226
rect 2506 3213 2509 3233
rect 2514 3223 2525 3226
rect 2474 3183 2493 3186
rect 2466 3163 2473 3166
rect 2442 3013 2445 3126
rect 2450 3086 2453 3126
rect 2458 3093 2461 3126
rect 2470 3106 2473 3163
rect 2482 3123 2485 3136
rect 2490 3133 2493 3183
rect 2466 3103 2473 3106
rect 2466 3086 2469 3103
rect 2490 3096 2493 3126
rect 2498 3103 2501 3206
rect 2514 3203 2517 3223
rect 2522 3153 2525 3216
rect 2530 3213 2533 3233
rect 2530 3146 2533 3206
rect 2522 3143 2549 3146
rect 2554 3143 2557 3206
rect 2570 3163 2573 3226
rect 2450 3083 2469 3086
rect 2482 3093 2493 3096
rect 2522 3093 2525 3143
rect 2546 3136 2549 3143
rect 2530 3123 2533 3136
rect 2538 3126 2541 3136
rect 2546 3133 2557 3136
rect 2538 3123 2565 3126
rect 2562 3106 2565 3123
rect 2554 3103 2565 3106
rect 2482 3066 2485 3093
rect 2474 3063 2485 3066
rect 2490 3066 2493 3086
rect 2490 3063 2501 3066
rect 2458 3013 2461 3036
rect 2474 3016 2477 3063
rect 2498 3016 2501 3063
rect 2554 3036 2557 3103
rect 2554 3033 2565 3036
rect 2474 3013 2485 3016
rect 2426 3003 2437 3006
rect 2378 2963 2397 2966
rect 2378 2933 2381 2963
rect 2394 2943 2429 2946
rect 2394 2923 2397 2943
rect 2402 2893 2405 2936
rect 2362 2813 2365 2826
rect 2370 2823 2389 2826
rect 2410 2823 2413 2926
rect 2418 2923 2421 2936
rect 2426 2933 2429 2943
rect 2442 2926 2445 3006
rect 2458 2983 2461 3006
rect 2482 2946 2485 3013
rect 2450 2943 2485 2946
rect 2490 3013 2501 3016
rect 2490 2933 2493 3013
rect 2530 3003 2533 3016
rect 2546 2973 2549 3006
rect 2506 2936 2509 2956
rect 2502 2933 2509 2936
rect 2426 2903 2429 2926
rect 2442 2923 2469 2926
rect 2466 2843 2469 2923
rect 2474 2883 2477 2926
rect 2502 2836 2505 2933
rect 2370 2803 2373 2816
rect 2322 2773 2333 2776
rect 2258 2763 2301 2766
rect 2162 2623 2169 2626
rect 2138 2543 2141 2596
rect 2146 2533 2149 2616
rect 2066 2456 2069 2496
rect 2066 2453 2073 2456
rect 2026 2443 2037 2446
rect 1954 2373 2013 2376
rect 1858 2343 1893 2346
rect 1890 2333 1893 2343
rect 1802 2303 1813 2306
rect 1682 2293 1701 2296
rect 1658 2256 1661 2276
rect 1658 2253 1669 2256
rect 1650 2203 1653 2246
rect 1666 2196 1669 2253
rect 1658 2193 1669 2196
rect 1658 2146 1661 2193
rect 1682 2186 1685 2293
rect 1706 2193 1709 2296
rect 1802 2226 1805 2303
rect 1826 2273 1829 2316
rect 1850 2313 1869 2316
rect 1746 2223 1765 2226
rect 1802 2223 1813 2226
rect 1818 2223 1821 2236
rect 1746 2216 1749 2223
rect 1714 2203 1717 2216
rect 1682 2183 1701 2186
rect 1650 2143 1661 2146
rect 1650 2083 1653 2143
rect 1650 2013 1653 2026
rect 1650 1943 1653 2006
rect 1650 1833 1653 1936
rect 1650 1813 1653 1826
rect 1650 1733 1653 1756
rect 1650 1693 1653 1726
rect 1658 1713 1661 2136
rect 1666 2113 1669 2136
rect 1666 1933 1669 2006
rect 1666 1903 1669 1926
rect 1674 1883 1677 2146
rect 1682 2013 1685 2026
rect 1690 2006 1693 2086
rect 1698 2076 1701 2183
rect 1722 2163 1725 2216
rect 1738 2213 1749 2216
rect 1730 2183 1733 2206
rect 1746 2193 1749 2206
rect 1754 2173 1757 2216
rect 1762 2213 1765 2223
rect 1762 2156 1765 2206
rect 1746 2143 1749 2156
rect 1758 2153 1765 2156
rect 1698 2073 1709 2076
rect 1698 2023 1701 2066
rect 1706 2033 1709 2073
rect 1682 2003 1693 2006
rect 1682 1923 1685 2003
rect 1698 1936 1701 2016
rect 1706 2003 1709 2026
rect 1690 1933 1701 1936
rect 1690 1906 1693 1933
rect 1686 1903 1693 1906
rect 1686 1836 1689 1903
rect 1698 1883 1701 1926
rect 1706 1873 1709 1946
rect 1714 1923 1717 2126
rect 1722 2033 1725 2136
rect 1722 2013 1725 2026
rect 1730 2006 1733 2106
rect 1738 2083 1741 2136
rect 1746 2113 1749 2126
rect 1758 2066 1761 2153
rect 1754 2063 1761 2066
rect 1738 2013 1741 2046
rect 1722 1953 1725 2006
rect 1730 2003 1741 2006
rect 1746 2003 1749 2056
rect 1738 1956 1741 2003
rect 1730 1953 1741 1956
rect 1722 1923 1725 1936
rect 1730 1903 1733 1953
rect 1738 1933 1741 1946
rect 1746 1926 1749 1976
rect 1738 1923 1749 1926
rect 1754 1923 1757 2063
rect 1762 1993 1765 2056
rect 1770 1983 1773 2176
rect 1778 2133 1781 2216
rect 1802 2186 1805 2206
rect 1794 2183 1805 2186
rect 1794 2136 1797 2183
rect 1794 2133 1805 2136
rect 1786 2043 1789 2116
rect 1666 1813 1669 1836
rect 1686 1833 1693 1836
rect 1674 1783 1677 1806
rect 1666 1696 1669 1736
rect 1682 1713 1685 1816
rect 1666 1693 1677 1696
rect 1650 1493 1653 1646
rect 1658 1616 1661 1666
rect 1674 1636 1677 1693
rect 1690 1646 1693 1833
rect 1698 1756 1701 1836
rect 1714 1803 1717 1866
rect 1722 1813 1725 1836
rect 1730 1806 1733 1846
rect 1722 1803 1733 1806
rect 1698 1753 1709 1756
rect 1698 1733 1701 1746
rect 1698 1663 1701 1726
rect 1706 1713 1709 1753
rect 1690 1643 1701 1646
rect 1674 1633 1685 1636
rect 1658 1613 1677 1616
rect 1658 1593 1661 1606
rect 1658 1543 1661 1566
rect 1674 1506 1677 1526
rect 1666 1503 1677 1506
rect 1666 1436 1669 1503
rect 1666 1433 1677 1436
rect 1650 1413 1669 1416
rect 1650 1303 1653 1396
rect 1658 1293 1661 1406
rect 1650 1203 1653 1226
rect 1658 1126 1661 1216
rect 1666 1213 1669 1413
rect 1674 1326 1677 1433
rect 1682 1423 1685 1633
rect 1690 1623 1693 1636
rect 1698 1573 1701 1643
rect 1690 1503 1693 1536
rect 1698 1513 1701 1526
rect 1706 1496 1709 1656
rect 1714 1616 1717 1746
rect 1722 1733 1725 1803
rect 1722 1703 1725 1726
rect 1730 1723 1733 1776
rect 1730 1633 1733 1646
rect 1722 1623 1733 1626
rect 1738 1623 1741 1923
rect 1746 1803 1749 1886
rect 1714 1613 1725 1616
rect 1714 1533 1717 1596
rect 1698 1493 1709 1496
rect 1682 1343 1685 1356
rect 1674 1323 1681 1326
rect 1690 1323 1693 1436
rect 1698 1393 1701 1493
rect 1698 1333 1701 1346
rect 1678 1246 1681 1323
rect 1674 1243 1681 1246
rect 1666 1133 1669 1146
rect 1650 1123 1661 1126
rect 1650 1083 1653 1123
rect 1666 1116 1669 1126
rect 1658 1113 1669 1116
rect 1650 823 1653 1006
rect 1658 816 1661 1113
rect 1666 1013 1669 1096
rect 1666 943 1669 966
rect 1666 893 1669 936
rect 1650 813 1661 816
rect 1650 806 1653 813
rect 1626 773 1633 776
rect 1642 803 1653 806
rect 1562 713 1573 716
rect 1538 593 1557 596
rect 1530 473 1533 526
rect 1498 433 1509 436
rect 1466 293 1477 296
rect 1466 236 1469 293
rect 1466 233 1477 236
rect 1458 203 1461 216
rect 1466 203 1469 216
rect 1474 193 1477 233
rect 1482 213 1485 406
rect 1498 386 1501 433
rect 1514 423 1525 426
rect 1530 393 1533 406
rect 1538 403 1541 593
rect 1562 586 1565 686
rect 1570 663 1573 713
rect 1546 583 1565 586
rect 1546 413 1549 583
rect 1498 383 1549 386
rect 1490 353 1517 356
rect 1490 333 1493 353
rect 1498 333 1501 346
rect 1514 336 1517 353
rect 1514 333 1525 336
rect 1490 306 1493 326
rect 1506 323 1517 326
rect 1490 303 1501 306
rect 1490 186 1493 296
rect 1498 213 1501 303
rect 1474 183 1493 186
rect 1442 143 1453 146
rect 1410 123 1421 126
rect 1426 93 1429 136
rect 1434 83 1437 126
rect 1450 96 1453 143
rect 1474 133 1477 183
rect 1482 143 1501 146
rect 1498 133 1501 143
rect 1498 113 1501 126
rect 1442 93 1453 96
rect 1442 73 1445 93
rect 1506 83 1509 206
rect 1514 203 1517 323
rect 1522 283 1525 326
rect 1530 303 1533 336
rect 1538 323 1541 346
rect 1546 293 1549 383
rect 1554 346 1557 526
rect 1562 513 1565 536
rect 1562 363 1565 466
rect 1570 453 1573 656
rect 1582 626 1585 743
rect 1594 723 1597 736
rect 1618 716 1621 726
rect 1626 723 1629 773
rect 1642 733 1645 803
rect 1666 746 1669 826
rect 1650 743 1669 746
rect 1618 713 1645 716
rect 1650 666 1653 743
rect 1658 703 1661 736
rect 1658 683 1661 696
rect 1578 623 1585 626
rect 1594 653 1605 656
rect 1578 576 1581 623
rect 1586 593 1589 606
rect 1578 573 1585 576
rect 1570 383 1573 406
rect 1582 346 1585 573
rect 1594 533 1597 653
rect 1618 633 1621 666
rect 1626 663 1653 666
rect 1666 663 1669 736
rect 1602 613 1605 626
rect 1602 513 1605 526
rect 1610 523 1613 626
rect 1618 593 1621 626
rect 1618 463 1621 536
rect 1626 473 1629 663
rect 1634 633 1637 656
rect 1634 623 1645 626
rect 1634 513 1637 623
rect 1650 613 1653 626
rect 1642 533 1645 546
rect 1650 516 1653 536
rect 1646 513 1653 516
rect 1594 413 1597 456
rect 1610 406 1613 416
rect 1602 403 1613 406
rect 1554 343 1561 346
rect 1558 286 1561 343
rect 1578 343 1585 346
rect 1554 283 1561 286
rect 1530 203 1533 226
rect 1538 196 1541 236
rect 1514 193 1541 196
rect 1514 133 1517 193
rect 1546 173 1549 216
rect 1554 203 1557 283
rect 1570 266 1573 336
rect 1566 263 1573 266
rect 1566 186 1569 263
rect 1566 183 1573 186
rect 1570 163 1573 183
rect 1570 123 1573 146
rect 1578 133 1581 343
rect 1602 333 1605 346
rect 1586 213 1589 326
rect 1618 323 1621 406
rect 1602 216 1605 236
rect 1602 213 1613 216
rect 1602 163 1605 206
rect 1618 203 1621 276
rect 1562 43 1565 116
rect 1586 103 1589 126
rect 1602 113 1605 136
rect 1618 103 1621 116
rect 1626 93 1629 456
rect 1634 403 1637 436
rect 1634 306 1637 366
rect 1646 356 1649 513
rect 1658 436 1661 536
rect 1666 506 1669 616
rect 1674 523 1677 1243
rect 1682 1203 1685 1226
rect 1690 1196 1693 1286
rect 1698 1203 1701 1256
rect 1690 1193 1701 1196
rect 1682 1133 1685 1146
rect 1682 1093 1685 1126
rect 1682 1023 1685 1056
rect 1690 943 1693 1136
rect 1698 1133 1701 1193
rect 1682 906 1685 926
rect 1682 903 1689 906
rect 1686 756 1689 903
rect 1698 843 1701 1126
rect 1706 853 1709 1486
rect 1730 1453 1733 1623
rect 1746 1606 1749 1736
rect 1754 1733 1757 1916
rect 1762 1743 1765 1946
rect 1770 1933 1773 1956
rect 1770 1843 1773 1926
rect 1770 1823 1773 1836
rect 1770 1736 1773 1816
rect 1778 1786 1781 2026
rect 1786 1923 1789 1996
rect 1794 1983 1797 2066
rect 1802 2043 1805 2133
rect 1802 1963 1805 2006
rect 1810 1946 1813 2223
rect 1818 2133 1821 2216
rect 1850 2203 1853 2306
rect 1818 2113 1821 2126
rect 1826 2056 1829 2166
rect 1834 2143 1853 2146
rect 1834 2123 1837 2143
rect 1842 2086 1845 2136
rect 1850 2133 1853 2143
rect 1850 2103 1853 2126
rect 1842 2083 1853 2086
rect 1826 2053 1837 2056
rect 1818 1993 1821 2016
rect 1810 1943 1821 1946
rect 1794 1933 1813 1936
rect 1786 1823 1789 1906
rect 1778 1783 1789 1786
rect 1762 1733 1773 1736
rect 1762 1716 1765 1726
rect 1778 1723 1781 1776
rect 1786 1763 1789 1783
rect 1742 1603 1749 1606
rect 1742 1466 1745 1603
rect 1754 1513 1757 1716
rect 1762 1713 1773 1716
rect 1742 1463 1749 1466
rect 1746 1443 1749 1463
rect 1730 1406 1733 1416
rect 1714 1403 1733 1406
rect 1714 1336 1717 1396
rect 1714 1333 1725 1336
rect 1714 1123 1717 1326
rect 1722 1133 1725 1333
rect 1730 1306 1733 1376
rect 1738 1313 1741 1406
rect 1746 1333 1749 1416
rect 1754 1396 1757 1506
rect 1762 1416 1765 1696
rect 1770 1523 1773 1713
rect 1778 1706 1781 1716
rect 1786 1713 1789 1736
rect 1778 1703 1789 1706
rect 1778 1526 1781 1646
rect 1794 1613 1797 1933
rect 1802 1693 1805 1926
rect 1810 1833 1813 1846
rect 1818 1826 1821 1943
rect 1826 1923 1829 2046
rect 1834 2013 1837 2053
rect 1842 1993 1845 2046
rect 1850 2013 1853 2083
rect 1858 2033 1861 2256
rect 1858 2006 1861 2026
rect 1850 2003 1861 2006
rect 1842 1946 1845 1966
rect 1838 1943 1845 1946
rect 1850 1963 1861 1966
rect 1826 1846 1829 1916
rect 1838 1866 1841 1943
rect 1838 1863 1845 1866
rect 1826 1843 1837 1846
rect 1810 1823 1821 1826
rect 1810 1676 1813 1823
rect 1834 1813 1837 1843
rect 1818 1773 1821 1806
rect 1842 1803 1845 1863
rect 1850 1796 1853 1963
rect 1858 1893 1861 1916
rect 1858 1833 1861 1886
rect 1866 1843 1869 2313
rect 1874 2306 1877 2326
rect 1898 2316 1901 2336
rect 1898 2313 1909 2316
rect 1922 2313 1933 2316
rect 1874 2303 1881 2306
rect 1878 2136 1881 2303
rect 1890 2203 1893 2286
rect 1906 2246 1909 2313
rect 1898 2243 1909 2246
rect 1898 2166 1901 2243
rect 1938 2233 1941 2326
rect 1954 2273 1957 2316
rect 1978 2303 1981 2336
rect 1986 2333 1989 2356
rect 2010 2333 2013 2373
rect 2018 2333 2021 2356
rect 2034 2346 2037 2443
rect 2050 2403 2053 2416
rect 2070 2396 2073 2453
rect 2082 2413 2085 2526
rect 2106 2523 2133 2526
rect 2154 2523 2157 2616
rect 2166 2556 2169 2623
rect 2178 2613 2189 2616
rect 2178 2603 2181 2613
rect 2194 2563 2197 2726
rect 2234 2723 2237 2736
rect 2202 2633 2221 2636
rect 2202 2603 2205 2633
rect 2218 2603 2221 2633
rect 2250 2613 2253 2736
rect 2266 2733 2269 2756
rect 2298 2696 2301 2763
rect 2330 2756 2333 2773
rect 2330 2753 2337 2756
rect 2314 2723 2317 2746
rect 2290 2693 2301 2696
rect 2162 2553 2169 2556
rect 2098 2403 2101 2436
rect 2026 2343 2037 2346
rect 2066 2393 2073 2396
rect 2026 2326 2029 2343
rect 2066 2326 2069 2393
rect 1994 2323 2045 2326
rect 2010 2283 2013 2316
rect 1978 2226 1981 2246
rect 1914 2223 1973 2226
rect 1978 2223 1989 2226
rect 1914 2213 1917 2223
rect 1890 2163 1901 2166
rect 1878 2133 1885 2136
rect 1874 1836 1877 2126
rect 1882 2056 1885 2133
rect 1890 2126 1893 2163
rect 1906 2136 1909 2206
rect 1922 2146 1925 2206
rect 1930 2173 1933 2216
rect 1954 2163 1957 2206
rect 1970 2173 1973 2206
rect 1986 2166 1989 2223
rect 2002 2176 2005 2256
rect 2042 2246 2045 2323
rect 2058 2323 2069 2326
rect 2058 2253 2061 2323
rect 2074 2316 2077 2376
rect 2082 2323 2085 2356
rect 2122 2346 2125 2416
rect 2106 2343 2125 2346
rect 2106 2333 2109 2343
rect 2130 2336 2133 2523
rect 2162 2493 2165 2553
rect 2170 2523 2173 2536
rect 2178 2413 2181 2526
rect 2186 2503 2189 2536
rect 2210 2533 2213 2556
rect 2202 2493 2205 2526
rect 2266 2523 2269 2636
rect 2290 2616 2293 2693
rect 2334 2686 2337 2753
rect 2354 2733 2357 2746
rect 2378 2743 2381 2816
rect 2330 2683 2337 2686
rect 2286 2613 2293 2616
rect 2286 2556 2289 2613
rect 2286 2553 2293 2556
rect 2114 2326 2117 2336
rect 2106 2323 2117 2326
rect 2122 2333 2133 2336
rect 2138 2333 2141 2406
rect 2194 2403 2197 2436
rect 2234 2426 2237 2446
rect 2226 2423 2237 2426
rect 2226 2366 2229 2423
rect 2242 2376 2245 2416
rect 2274 2413 2277 2526
rect 2282 2523 2285 2536
rect 2290 2443 2293 2553
rect 2298 2533 2301 2606
rect 2314 2563 2317 2616
rect 2330 2556 2333 2683
rect 2346 2633 2349 2726
rect 2338 2613 2365 2616
rect 2370 2606 2373 2656
rect 2386 2633 2389 2823
rect 2394 2813 2413 2816
rect 2410 2783 2413 2806
rect 2418 2803 2421 2826
rect 2474 2803 2477 2836
rect 2502 2833 2509 2836
rect 2498 2783 2501 2816
rect 2394 2723 2397 2736
rect 2418 2666 2421 2756
rect 2466 2723 2469 2746
rect 2498 2666 2501 2726
rect 2506 2696 2509 2833
rect 2514 2813 2517 2936
rect 2538 2933 2541 2946
rect 2546 2933 2549 2966
rect 2554 2936 2557 3016
rect 2562 3006 2565 3033
rect 2570 3013 2573 3036
rect 2578 3013 2581 3176
rect 2586 3096 2589 3206
rect 2634 3193 2637 3216
rect 2706 3206 2709 3216
rect 2698 3203 2709 3206
rect 2714 3203 2717 3216
rect 2722 3213 2725 3226
rect 2738 3223 2741 3236
rect 2762 3213 2789 3216
rect 2794 3213 2797 3266
rect 2802 3213 2813 3216
rect 2858 3213 2861 3236
rect 2866 3223 2877 3226
rect 2594 3103 2597 3126
rect 2602 3123 2605 3156
rect 2586 3093 2597 3096
rect 2594 3056 2597 3093
rect 2618 3073 2621 3166
rect 2626 3143 2653 3146
rect 2626 3133 2629 3143
rect 2626 3113 2629 3126
rect 2634 3123 2637 3136
rect 2682 3123 2685 3136
rect 2690 3123 2693 3136
rect 2698 3106 2701 3203
rect 2706 3133 2709 3196
rect 2762 3193 2765 3206
rect 2770 3183 2773 3206
rect 2786 3203 2789 3213
rect 2778 3193 2789 3196
rect 2794 3193 2797 3206
rect 2738 3143 2781 3146
rect 2738 3133 2741 3143
rect 2690 3103 2701 3106
rect 2714 3103 2717 3126
rect 2594 3053 2605 3056
rect 2562 3003 2573 3006
rect 2554 2933 2565 2936
rect 2522 2923 2541 2926
rect 2562 2916 2565 2933
rect 2570 2923 2573 3003
rect 2578 2973 2581 3006
rect 2602 2976 2605 3053
rect 2642 3003 2645 3016
rect 2650 3003 2653 3026
rect 2594 2973 2605 2976
rect 2594 2933 2597 2973
rect 2538 2913 2565 2916
rect 2554 2813 2557 2826
rect 2538 2733 2541 2756
rect 2570 2723 2573 2806
rect 2578 2793 2581 2926
rect 2618 2923 2621 2946
rect 2626 2916 2629 2986
rect 2642 2976 2645 2996
rect 2622 2913 2629 2916
rect 2638 2973 2645 2976
rect 2602 2813 2605 2826
rect 2602 2743 2605 2806
rect 2610 2793 2613 2896
rect 2622 2846 2625 2913
rect 2638 2906 2641 2973
rect 2658 2966 2661 3036
rect 2690 2996 2693 3103
rect 2714 3003 2717 3096
rect 2738 3033 2741 3126
rect 2746 3123 2749 3136
rect 2754 2996 2757 3016
rect 2762 3013 2765 3136
rect 2770 3123 2773 3136
rect 2778 3133 2781 3143
rect 2794 3123 2797 3136
rect 2810 3123 2813 3186
rect 2850 3133 2853 3206
rect 2866 3136 2869 3223
rect 2882 3216 2885 3226
rect 2874 3213 2885 3216
rect 2874 3203 2877 3213
rect 2890 3146 2893 3216
rect 2898 3173 2901 3236
rect 2914 3203 2917 3266
rect 3306 3253 3349 3256
rect 2938 3223 2973 3226
rect 2922 3146 2925 3216
rect 2954 3213 2973 3216
rect 2994 3213 2997 3236
rect 3018 3233 3069 3236
rect 2970 3156 2973 3206
rect 2978 3193 2981 3206
rect 2986 3203 2997 3206
rect 2970 3153 2997 3156
rect 2890 3143 2925 3146
rect 2866 3133 2877 3136
rect 2866 3106 2869 3126
rect 2858 3103 2869 3106
rect 2858 3026 2861 3103
rect 2794 3013 2797 3026
rect 2834 3023 2861 3026
rect 2690 2993 2701 2996
rect 2698 2976 2701 2993
rect 2674 2973 2701 2976
rect 2746 2993 2757 2996
rect 2658 2963 2665 2966
rect 2662 2916 2665 2963
rect 2658 2913 2665 2916
rect 2638 2903 2645 2906
rect 2642 2886 2645 2903
rect 2658 2893 2661 2913
rect 2634 2883 2645 2886
rect 2674 2846 2677 2973
rect 2682 2923 2685 2966
rect 2690 2933 2693 2946
rect 2714 2933 2717 2956
rect 2746 2946 2749 2993
rect 2746 2943 2757 2946
rect 2618 2843 2625 2846
rect 2650 2843 2677 2846
rect 2618 2776 2621 2843
rect 2614 2773 2621 2776
rect 2614 2706 2617 2773
rect 2626 2713 2629 2826
rect 2650 2793 2653 2843
rect 2682 2816 2685 2856
rect 2674 2813 2685 2816
rect 2698 2826 2701 2926
rect 2746 2906 2749 2926
rect 2742 2903 2749 2906
rect 2742 2826 2745 2903
rect 2698 2823 2733 2826
rect 2742 2823 2749 2826
rect 2650 2733 2653 2756
rect 2674 2733 2677 2813
rect 2614 2703 2621 2706
rect 2506 2693 2517 2696
rect 2394 2663 2421 2666
rect 2474 2663 2501 2666
rect 2354 2603 2373 2606
rect 2394 2603 2397 2663
rect 2410 2653 2437 2656
rect 2354 2583 2357 2603
rect 2306 2523 2309 2556
rect 2314 2553 2333 2556
rect 2290 2403 2293 2436
rect 2314 2396 2317 2553
rect 2322 2503 2325 2536
rect 2370 2533 2373 2546
rect 2346 2456 2349 2526
rect 2362 2463 2365 2526
rect 2370 2516 2373 2526
rect 2378 2523 2381 2566
rect 2386 2516 2389 2526
rect 2370 2513 2389 2516
rect 2402 2493 2405 2616
rect 2410 2603 2413 2653
rect 2418 2546 2421 2636
rect 2426 2603 2429 2616
rect 2434 2603 2437 2653
rect 2474 2613 2477 2663
rect 2514 2636 2517 2693
rect 2506 2633 2517 2636
rect 2442 2596 2445 2606
rect 2414 2543 2421 2546
rect 2434 2593 2445 2596
rect 2414 2496 2417 2543
rect 2426 2503 2429 2536
rect 2434 2506 2437 2593
rect 2490 2553 2493 2616
rect 2498 2596 2501 2606
rect 2506 2603 2509 2633
rect 2514 2613 2557 2616
rect 2562 2613 2565 2636
rect 2514 2603 2517 2613
rect 2522 2596 2525 2606
rect 2498 2593 2533 2596
rect 2498 2536 2501 2566
rect 2442 2533 2469 2536
rect 2490 2533 2501 2536
rect 2522 2533 2525 2576
rect 2530 2536 2533 2593
rect 2530 2533 2549 2536
rect 2554 2533 2557 2613
rect 2562 2603 2581 2606
rect 2442 2513 2445 2533
rect 2450 2523 2557 2526
rect 2554 2516 2557 2523
rect 2554 2513 2565 2516
rect 2570 2506 2573 2556
rect 2586 2546 2589 2646
rect 2594 2553 2597 2616
rect 2586 2543 2597 2546
rect 2434 2503 2453 2506
rect 2414 2493 2421 2496
rect 2346 2453 2373 2456
rect 2306 2393 2317 2396
rect 2242 2373 2269 2376
rect 2226 2363 2253 2366
rect 2066 2313 2077 2316
rect 2042 2243 2053 2246
rect 2010 2186 2013 2216
rect 2026 2213 2029 2226
rect 2034 2193 2037 2206
rect 2010 2183 2037 2186
rect 2002 2173 2029 2176
rect 1978 2163 1989 2166
rect 1922 2143 1941 2146
rect 1906 2133 1925 2136
rect 1890 2123 1909 2126
rect 1882 2053 1901 2056
rect 1882 1963 1885 2006
rect 1882 1923 1885 1946
rect 1890 1933 1893 1996
rect 1866 1833 1877 1836
rect 1826 1793 1853 1796
rect 1806 1673 1813 1676
rect 1786 1536 1789 1606
rect 1806 1556 1809 1673
rect 1818 1616 1821 1736
rect 1826 1723 1829 1793
rect 1858 1776 1861 1826
rect 1854 1773 1861 1776
rect 1826 1623 1829 1666
rect 1834 1636 1837 1736
rect 1842 1663 1845 1756
rect 1854 1716 1857 1773
rect 1854 1713 1861 1716
rect 1834 1633 1845 1636
rect 1818 1613 1837 1616
rect 1806 1553 1813 1556
rect 1786 1533 1805 1536
rect 1778 1523 1797 1526
rect 1770 1483 1773 1516
rect 1778 1423 1781 1436
rect 1762 1413 1781 1416
rect 1754 1393 1761 1396
rect 1730 1303 1749 1306
rect 1730 1203 1733 1226
rect 1738 1156 1741 1236
rect 1730 1153 1741 1156
rect 1730 1126 1733 1153
rect 1738 1133 1741 1146
rect 1730 1123 1741 1126
rect 1746 1116 1749 1303
rect 1758 1266 1761 1393
rect 1770 1276 1773 1376
rect 1778 1323 1781 1413
rect 1786 1333 1789 1523
rect 1794 1503 1797 1516
rect 1778 1293 1781 1316
rect 1794 1313 1797 1426
rect 1802 1413 1805 1533
rect 1802 1313 1805 1396
rect 1786 1283 1789 1306
rect 1770 1273 1781 1276
rect 1730 1113 1749 1116
rect 1754 1263 1761 1266
rect 1714 913 1717 1076
rect 1722 1003 1725 1026
rect 1722 823 1725 946
rect 1706 803 1717 806
rect 1706 773 1709 796
rect 1682 753 1689 756
rect 1682 733 1685 753
rect 1698 743 1701 766
rect 1698 686 1701 726
rect 1714 703 1717 803
rect 1690 683 1701 686
rect 1690 626 1693 683
rect 1682 623 1693 626
rect 1682 603 1685 623
rect 1706 613 1709 626
rect 1714 623 1717 696
rect 1682 513 1685 526
rect 1666 503 1673 506
rect 1670 446 1673 503
rect 1670 443 1677 446
rect 1658 433 1669 436
rect 1658 403 1661 426
rect 1666 403 1669 433
rect 1646 353 1653 356
rect 1642 323 1645 336
rect 1634 303 1641 306
rect 1638 236 1641 303
rect 1650 266 1653 353
rect 1658 333 1661 376
rect 1674 313 1677 443
rect 1690 403 1693 536
rect 1706 426 1709 606
rect 1722 533 1725 816
rect 1730 803 1733 1113
rect 1754 1036 1757 1263
rect 1762 1223 1765 1246
rect 1770 1206 1773 1266
rect 1778 1226 1781 1273
rect 1786 1243 1805 1246
rect 1786 1233 1789 1243
rect 1778 1223 1789 1226
rect 1794 1223 1797 1236
rect 1802 1233 1805 1243
rect 1786 1216 1789 1223
rect 1766 1203 1773 1206
rect 1766 1136 1769 1203
rect 1778 1173 1781 1216
rect 1786 1213 1793 1216
rect 1790 1146 1793 1213
rect 1802 1153 1805 1226
rect 1790 1143 1797 1146
rect 1762 1133 1769 1136
rect 1762 1083 1765 1133
rect 1770 1076 1773 1126
rect 1778 1123 1789 1126
rect 1770 1073 1789 1076
rect 1754 1033 1781 1036
rect 1738 996 1741 1016
rect 1746 1013 1749 1026
rect 1738 993 1749 996
rect 1730 593 1733 706
rect 1738 696 1741 986
rect 1746 973 1749 993
rect 1746 713 1749 966
rect 1738 693 1745 696
rect 1742 606 1745 693
rect 1738 603 1745 606
rect 1738 583 1741 603
rect 1754 536 1757 986
rect 1762 893 1765 926
rect 1762 703 1765 806
rect 1770 803 1773 1026
rect 1778 956 1781 1033
rect 1786 963 1789 1073
rect 1794 983 1797 1143
rect 1802 1023 1805 1126
rect 1778 953 1789 956
rect 1778 733 1781 946
rect 1786 906 1789 953
rect 1794 923 1797 956
rect 1786 903 1793 906
rect 1790 826 1793 903
rect 1786 823 1793 826
rect 1770 693 1773 716
rect 1778 686 1781 726
rect 1762 683 1781 686
rect 1762 623 1765 683
rect 1786 676 1789 823
rect 1794 683 1797 806
rect 1802 706 1805 1006
rect 1810 923 1813 1553
rect 1818 1533 1821 1606
rect 1826 1583 1829 1606
rect 1818 1456 1821 1516
rect 1834 1473 1837 1536
rect 1818 1453 1837 1456
rect 1818 1423 1821 1453
rect 1826 1416 1829 1446
rect 1834 1423 1837 1453
rect 1826 1413 1837 1416
rect 1842 1413 1845 1633
rect 1850 1623 1853 1696
rect 1850 1593 1853 1616
rect 1858 1586 1861 1713
rect 1850 1583 1861 1586
rect 1850 1513 1853 1583
rect 1866 1576 1869 1833
rect 1874 1823 1885 1826
rect 1874 1743 1877 1823
rect 1890 1813 1893 1906
rect 1874 1633 1877 1726
rect 1882 1696 1885 1736
rect 1890 1723 1893 1746
rect 1898 1723 1901 2053
rect 1906 2013 1909 2123
rect 1922 2116 1925 2133
rect 1938 2123 1941 2143
rect 1914 2103 1917 2116
rect 1922 2113 1941 2116
rect 1938 2106 1941 2113
rect 1922 2023 1925 2036
rect 1930 2026 1933 2106
rect 1938 2103 1949 2106
rect 1938 2033 1941 2066
rect 1930 2023 1941 2026
rect 1946 2023 1949 2103
rect 1954 2023 1957 2116
rect 1962 2093 1965 2126
rect 1978 2113 1981 2163
rect 1994 2133 1997 2146
rect 2002 2123 2005 2166
rect 1914 2013 1933 2016
rect 1906 1943 1909 2006
rect 1906 1893 1909 1926
rect 1914 1903 1917 2013
rect 1938 2006 1941 2023
rect 1930 2003 1941 2006
rect 1922 1933 1925 1966
rect 1906 1813 1909 1826
rect 1906 1746 1909 1766
rect 1914 1753 1917 1856
rect 1922 1746 1925 1926
rect 1930 1813 1933 2003
rect 1938 1883 1941 1966
rect 1906 1743 1917 1746
rect 1922 1743 1933 1746
rect 1914 1736 1917 1743
rect 1914 1733 1925 1736
rect 1906 1723 1917 1726
rect 1882 1693 1889 1696
rect 1886 1636 1889 1693
rect 1898 1663 1901 1716
rect 1906 1683 1909 1723
rect 1882 1633 1889 1636
rect 1882 1616 1885 1633
rect 1858 1573 1869 1576
rect 1874 1613 1885 1616
rect 1890 1613 1901 1616
rect 1858 1543 1861 1573
rect 1874 1526 1877 1613
rect 1882 1583 1885 1606
rect 1890 1533 1893 1613
rect 1906 1606 1909 1636
rect 1914 1613 1917 1646
rect 1898 1603 1909 1606
rect 1866 1523 1877 1526
rect 1866 1456 1869 1523
rect 1866 1453 1877 1456
rect 1858 1423 1861 1436
rect 1818 1053 1821 1406
rect 1826 1043 1829 1406
rect 1834 1313 1837 1413
rect 1842 1396 1845 1406
rect 1842 1393 1869 1396
rect 1834 1156 1837 1286
rect 1858 1256 1861 1336
rect 1866 1333 1869 1393
rect 1874 1373 1877 1453
rect 1882 1346 1885 1526
rect 1890 1353 1893 1436
rect 1874 1336 1877 1346
rect 1882 1343 1893 1346
rect 1874 1333 1885 1336
rect 1866 1323 1877 1326
rect 1890 1316 1893 1343
rect 1886 1313 1893 1316
rect 1842 1223 1845 1256
rect 1858 1253 1869 1256
rect 1866 1246 1869 1253
rect 1858 1223 1861 1246
rect 1866 1243 1877 1246
rect 1842 1163 1845 1216
rect 1866 1206 1869 1243
rect 1858 1203 1869 1206
rect 1834 1153 1845 1156
rect 1810 733 1813 856
rect 1818 716 1821 1026
rect 1826 963 1829 1026
rect 1834 993 1837 1146
rect 1842 986 1845 1153
rect 1850 1013 1853 1176
rect 1858 1146 1861 1203
rect 1874 1183 1877 1226
rect 1886 1206 1889 1313
rect 1898 1213 1901 1603
rect 1922 1586 1925 1733
rect 1930 1703 1933 1743
rect 1930 1633 1933 1696
rect 1938 1683 1941 1806
rect 1930 1616 1933 1626
rect 1938 1623 1941 1636
rect 1930 1613 1941 1616
rect 1930 1593 1933 1606
rect 1938 1603 1941 1613
rect 1914 1583 1925 1586
rect 1906 1406 1909 1576
rect 1914 1503 1917 1583
rect 1914 1413 1917 1436
rect 1906 1403 1917 1406
rect 1906 1333 1909 1346
rect 1914 1326 1917 1403
rect 1906 1323 1917 1326
rect 1886 1203 1893 1206
rect 1858 1143 1877 1146
rect 1834 983 1845 986
rect 1826 853 1829 916
rect 1826 763 1829 806
rect 1834 776 1837 983
rect 1842 823 1845 946
rect 1850 943 1853 1006
rect 1858 1003 1861 1143
rect 1866 996 1869 1136
rect 1862 993 1869 996
rect 1850 843 1853 936
rect 1862 876 1865 993
rect 1874 923 1877 1143
rect 1882 1123 1885 1166
rect 1890 1093 1893 1203
rect 1882 1023 1885 1036
rect 1882 993 1885 1006
rect 1858 873 1865 876
rect 1842 793 1845 806
rect 1850 783 1853 826
rect 1834 773 1841 776
rect 1826 723 1829 746
rect 1818 713 1829 716
rect 1802 703 1821 706
rect 1786 673 1813 676
rect 1770 613 1773 626
rect 1778 623 1789 626
rect 1746 533 1757 536
rect 1746 523 1749 533
rect 1762 526 1765 606
rect 1778 526 1781 623
rect 1794 613 1797 626
rect 1794 583 1797 606
rect 1810 603 1813 673
rect 1818 573 1821 703
rect 1826 566 1829 713
rect 1838 616 1841 773
rect 1858 766 1861 873
rect 1850 763 1861 766
rect 1754 523 1765 526
rect 1770 523 1781 526
rect 1794 563 1829 566
rect 1834 613 1841 616
rect 1730 436 1733 506
rect 1746 473 1749 516
rect 1754 496 1757 523
rect 1770 516 1773 523
rect 1762 513 1773 516
rect 1754 493 1765 496
rect 1714 433 1733 436
rect 1698 423 1709 426
rect 1714 423 1733 426
rect 1698 403 1701 423
rect 1714 416 1717 423
rect 1706 413 1717 416
rect 1682 296 1685 316
rect 1678 293 1685 296
rect 1650 263 1661 266
rect 1634 233 1641 236
rect 1634 173 1637 233
rect 1658 203 1661 263
rect 1678 236 1681 293
rect 1666 196 1669 236
rect 1658 193 1669 196
rect 1674 233 1681 236
rect 1658 123 1661 193
rect 1674 106 1677 233
rect 1690 213 1693 306
rect 1698 223 1701 396
rect 1706 313 1709 413
rect 1722 336 1725 416
rect 1738 343 1757 346
rect 1714 333 1725 336
rect 1714 316 1717 333
rect 1730 323 1733 336
rect 1738 323 1741 343
rect 1746 316 1749 336
rect 1754 333 1757 343
rect 1714 313 1749 316
rect 1754 293 1757 326
rect 1762 316 1765 493
rect 1794 476 1797 563
rect 1794 473 1805 476
rect 1802 453 1805 473
rect 1786 423 1805 426
rect 1778 413 1797 416
rect 1770 323 1773 406
rect 1802 363 1805 423
rect 1810 373 1813 526
rect 1818 483 1821 536
rect 1818 403 1821 456
rect 1826 403 1829 526
rect 1834 386 1837 613
rect 1842 533 1845 596
rect 1850 576 1853 726
rect 1858 713 1861 763
rect 1866 603 1869 856
rect 1874 693 1877 836
rect 1882 833 1885 936
rect 1882 783 1885 816
rect 1890 796 1893 1016
rect 1898 943 1901 1146
rect 1906 1033 1909 1323
rect 1898 903 1901 926
rect 1906 893 1909 1026
rect 1898 813 1901 846
rect 1914 816 1917 1316
rect 1922 1013 1925 1576
rect 1946 1556 1949 1916
rect 1954 1806 1957 1996
rect 1962 1813 1965 2066
rect 1978 1993 1981 2036
rect 1986 2013 1989 2066
rect 1970 1823 1973 1946
rect 1978 1916 1981 1926
rect 1978 1913 1989 1916
rect 1994 1913 1997 2086
rect 1978 1833 1981 1906
rect 1986 1883 1989 1913
rect 1970 1806 1973 1816
rect 1954 1803 1973 1806
rect 1954 1756 1957 1776
rect 1978 1766 1981 1826
rect 1986 1803 1989 1826
rect 1994 1783 1997 1816
rect 1970 1763 1981 1766
rect 1954 1753 1961 1756
rect 1958 1666 1961 1753
rect 1970 1723 1973 1763
rect 1978 1716 1981 1756
rect 1994 1723 1997 1736
rect 1970 1713 1981 1716
rect 1954 1663 1961 1666
rect 1954 1643 1957 1663
rect 1954 1573 1957 1636
rect 1962 1603 1965 1626
rect 1946 1553 1965 1556
rect 1930 1543 1957 1546
rect 1930 1533 1933 1543
rect 1962 1536 1965 1553
rect 1930 1513 1933 1526
rect 1930 1423 1933 1456
rect 1938 1406 1941 1536
rect 1934 1403 1941 1406
rect 1946 1533 1965 1536
rect 1934 1336 1937 1403
rect 1930 1333 1937 1336
rect 1930 1263 1933 1333
rect 1930 1213 1933 1226
rect 1930 1023 1933 1206
rect 1938 1133 1941 1326
rect 1938 1056 1941 1126
rect 1946 1063 1949 1533
rect 1954 1483 1957 1526
rect 1970 1443 1973 1706
rect 1954 1313 1957 1416
rect 1978 1413 1981 1706
rect 1986 1696 1989 1716
rect 1986 1693 1993 1696
rect 1990 1626 1993 1693
rect 1986 1623 1993 1626
rect 1986 1563 1989 1623
rect 1994 1583 1997 1606
rect 2002 1563 2005 2116
rect 2010 1706 2013 2136
rect 2018 2123 2021 2136
rect 2018 2023 2021 2046
rect 2018 1943 2021 2006
rect 2018 1916 2021 1936
rect 2026 1933 2029 2173
rect 2034 2036 2037 2183
rect 2042 2083 2045 2216
rect 2050 2126 2053 2243
rect 2058 2133 2061 2156
rect 2066 2133 2069 2313
rect 2082 2303 2085 2316
rect 2050 2123 2069 2126
rect 2074 2123 2077 2256
rect 2090 2223 2101 2226
rect 2106 2213 2109 2323
rect 2122 2226 2125 2333
rect 2114 2223 2125 2226
rect 2058 2063 2061 2086
rect 2034 2033 2061 2036
rect 2034 2013 2037 2033
rect 2042 2003 2045 2026
rect 2058 2013 2061 2033
rect 2066 2006 2069 2123
rect 2050 2003 2069 2006
rect 2042 1936 2045 1996
rect 2034 1933 2045 1936
rect 2018 1913 2025 1916
rect 2022 1826 2025 1913
rect 2018 1823 2025 1826
rect 2018 1773 2021 1823
rect 2026 1776 2029 1806
rect 2034 1783 2037 1933
rect 2050 1926 2053 2003
rect 2058 1943 2069 1946
rect 2074 1943 2077 2076
rect 2042 1923 2053 1926
rect 2058 1923 2061 1936
rect 2066 1933 2069 1943
rect 2082 1936 2085 2206
rect 2114 2156 2117 2223
rect 2090 2133 2093 2156
rect 2106 2153 2117 2156
rect 2122 2166 2125 2216
rect 2138 2213 2141 2236
rect 2154 2226 2157 2316
rect 2150 2223 2157 2226
rect 2130 2193 2133 2206
rect 2122 2163 2133 2166
rect 2090 2033 2093 2116
rect 2090 1986 2093 2016
rect 2098 1996 2101 2146
rect 2106 2113 2109 2153
rect 2114 2113 2117 2146
rect 2122 2063 2125 2163
rect 2130 2133 2133 2163
rect 2130 2113 2133 2126
rect 2138 2073 2141 2176
rect 2150 2146 2153 2223
rect 2150 2143 2157 2146
rect 2146 2103 2149 2126
rect 2130 2063 2149 2066
rect 2130 2056 2133 2063
rect 2114 2053 2133 2056
rect 2106 2003 2109 2046
rect 2114 2013 2117 2053
rect 2122 2013 2133 2016
rect 2138 2013 2141 2056
rect 2146 2016 2149 2063
rect 2154 2026 2157 2143
rect 2162 2066 2165 2216
rect 2170 2203 2173 2216
rect 2178 2186 2181 2336
rect 2242 2333 2245 2356
rect 2186 2323 2245 2326
rect 2226 2273 2229 2316
rect 2234 2283 2237 2316
rect 2174 2183 2181 2186
rect 2186 2213 2205 2216
rect 2218 2213 2221 2236
rect 2174 2096 2177 2183
rect 2186 2106 2189 2213
rect 2194 2196 2197 2206
rect 2202 2203 2205 2213
rect 2226 2196 2229 2206
rect 2194 2193 2229 2196
rect 2194 2123 2197 2193
rect 2234 2183 2237 2216
rect 2242 2213 2245 2323
rect 2250 2223 2253 2363
rect 2258 2273 2261 2366
rect 2266 2333 2269 2373
rect 2298 2333 2301 2356
rect 2250 2203 2261 2206
rect 2202 2133 2229 2136
rect 2202 2123 2221 2126
rect 2186 2103 2197 2106
rect 2174 2093 2181 2096
rect 2162 2063 2173 2066
rect 2154 2023 2165 2026
rect 2146 2013 2157 2016
rect 2138 1996 2141 2006
rect 2098 1993 2141 1996
rect 2090 1983 2109 1986
rect 2090 1943 2093 1976
rect 2082 1933 2093 1936
rect 2042 1823 2045 1896
rect 2026 1773 2037 1776
rect 2018 1733 2021 1766
rect 2026 1723 2029 1756
rect 2034 1733 2037 1746
rect 2010 1703 2021 1706
rect 2018 1636 2021 1703
rect 2042 1663 2045 1816
rect 2018 1633 2029 1636
rect 2018 1613 2021 1626
rect 2026 1616 2029 1633
rect 2026 1613 2037 1616
rect 1986 1466 1989 1526
rect 1994 1483 1997 1536
rect 2010 1533 2013 1606
rect 2002 1523 2013 1526
rect 2018 1523 2021 1546
rect 1986 1463 1993 1466
rect 1990 1406 1993 1463
rect 1962 1283 1965 1406
rect 1986 1403 1993 1406
rect 1986 1346 1989 1403
rect 1970 1333 1973 1346
rect 1986 1343 1993 1346
rect 1970 1276 1973 1326
rect 1962 1273 1973 1276
rect 1938 1053 1949 1056
rect 1946 1023 1949 1053
rect 1954 1016 1957 1216
rect 1930 1013 1957 1016
rect 1962 1013 1965 1273
rect 1978 1223 1981 1336
rect 1990 1256 1993 1343
rect 1986 1253 1993 1256
rect 1986 1216 1989 1253
rect 1986 1213 1997 1216
rect 1970 1153 1973 1186
rect 1978 1146 1981 1206
rect 1970 1143 1981 1146
rect 1970 1113 1973 1143
rect 1970 1036 1973 1106
rect 1978 1053 1981 1126
rect 1970 1033 1977 1036
rect 1930 1006 1933 1013
rect 1922 1003 1933 1006
rect 1938 1003 1949 1006
rect 1922 923 1925 946
rect 1930 936 1933 1003
rect 1930 933 1949 936
rect 1910 813 1917 816
rect 1890 793 1897 796
rect 1894 736 1897 793
rect 1910 746 1913 813
rect 1922 783 1925 806
rect 1930 776 1933 816
rect 1938 786 1941 846
rect 1946 803 1949 916
rect 1954 903 1957 996
rect 1962 933 1965 1006
rect 1974 946 1977 1033
rect 1970 943 1977 946
rect 1970 923 1973 943
rect 1986 836 1989 1206
rect 1994 1153 1997 1213
rect 2002 1123 2005 1476
rect 2010 1403 2013 1523
rect 2018 1346 2021 1506
rect 2010 1343 2021 1346
rect 2010 1143 2013 1343
rect 2018 1323 2021 1336
rect 2026 1333 2029 1613
rect 2034 1596 2037 1606
rect 2042 1603 2045 1626
rect 2050 1596 2053 1806
rect 2034 1593 2053 1596
rect 2034 1323 2037 1536
rect 2042 1473 2045 1566
rect 2050 1523 2053 1576
rect 2058 1506 2061 1916
rect 2066 1863 2069 1926
rect 2066 1696 2069 1856
rect 2074 1733 2077 1816
rect 2082 1803 2085 1926
rect 2090 1923 2093 1933
rect 2106 1916 2109 1983
rect 2106 1913 2113 1916
rect 2090 1736 2093 1816
rect 2098 1803 2101 1906
rect 2110 1836 2113 1913
rect 2122 1883 2125 1936
rect 2106 1833 2113 1836
rect 2106 1803 2109 1833
rect 2082 1733 2093 1736
rect 2066 1693 2077 1696
rect 2054 1503 2061 1506
rect 2042 1393 2045 1446
rect 2054 1436 2057 1503
rect 2054 1433 2061 1436
rect 2050 1346 2053 1416
rect 2058 1386 2061 1433
rect 2066 1403 2069 1686
rect 2074 1486 2077 1693
rect 2082 1603 2085 1636
rect 2090 1596 2093 1616
rect 2098 1613 2101 1666
rect 2082 1593 2093 1596
rect 2082 1533 2085 1593
rect 2106 1543 2109 1726
rect 2114 1723 2117 1766
rect 2122 1746 2125 1816
rect 2130 1803 2133 1993
rect 2162 1976 2165 2023
rect 2170 2013 2173 2063
rect 2154 1973 2165 1976
rect 2138 1923 2141 1966
rect 2146 1883 2149 1936
rect 2154 1876 2157 1973
rect 2178 1966 2181 2093
rect 2162 1963 2181 1966
rect 2162 1923 2165 1936
rect 2170 1923 2173 1946
rect 2186 1936 2189 2026
rect 2202 1986 2205 2123
rect 2226 2116 2229 2133
rect 2234 2123 2237 2136
rect 2242 2123 2253 2126
rect 2258 2123 2261 2203
rect 2210 2016 2213 2086
rect 2218 2023 2221 2116
rect 2226 2113 2249 2116
rect 2210 2013 2221 2016
rect 2202 1983 2221 1986
rect 2178 1933 2189 1936
rect 2194 1973 2213 1976
rect 2162 1903 2165 1916
rect 2138 1873 2157 1876
rect 2122 1743 2133 1746
rect 2114 1663 2117 1716
rect 2090 1523 2093 1536
rect 2074 1483 2085 1486
rect 2074 1423 2077 1476
rect 2058 1383 2065 1386
rect 2042 1343 2053 1346
rect 2042 1323 2045 1343
rect 2042 1296 2045 1316
rect 2022 1293 2045 1296
rect 2022 1236 2025 1293
rect 2018 1233 2025 1236
rect 2018 1196 2021 1233
rect 2026 1203 2029 1216
rect 2018 1193 2029 1196
rect 2010 1116 2013 1136
rect 1994 1113 2013 1116
rect 1994 903 1997 1106
rect 2002 1013 2005 1106
rect 2010 1053 2013 1106
rect 2018 1003 2021 1136
rect 2026 1056 2029 1193
rect 2034 1076 2037 1286
rect 2050 1283 2053 1336
rect 2062 1316 2065 1383
rect 2062 1313 2069 1316
rect 2042 1123 2045 1266
rect 2050 1183 2053 1226
rect 2058 1223 2061 1306
rect 2066 1266 2069 1313
rect 2074 1303 2077 1416
rect 2082 1343 2085 1483
rect 2090 1413 2093 1436
rect 2082 1323 2085 1336
rect 2074 1283 2085 1286
rect 2066 1263 2073 1266
rect 2058 1173 2061 1206
rect 2070 1156 2073 1263
rect 2082 1223 2085 1283
rect 2082 1183 2085 1206
rect 2090 1166 2093 1406
rect 2098 1333 2101 1536
rect 2114 1533 2117 1546
rect 2106 1426 2109 1436
rect 2114 1433 2117 1446
rect 2122 1436 2125 1736
rect 2130 1443 2133 1743
rect 2138 1616 2141 1873
rect 2162 1813 2165 1886
rect 2178 1883 2181 1933
rect 2186 1903 2189 1926
rect 2194 1923 2197 1973
rect 2178 1813 2181 1856
rect 2146 1723 2149 1806
rect 2170 1763 2173 1806
rect 2146 1683 2149 1716
rect 2154 1633 2157 1736
rect 2162 1733 2173 1736
rect 2170 1683 2173 1716
rect 2162 1623 2165 1656
rect 2178 1623 2181 1806
rect 2186 1793 2189 1816
rect 2194 1803 2197 1866
rect 2186 1643 2189 1786
rect 2138 1613 2157 1616
rect 2138 1453 2141 1606
rect 2122 1433 2141 1436
rect 2106 1423 2125 1426
rect 2106 1406 2109 1416
rect 2130 1413 2133 1426
rect 2106 1403 2133 1406
rect 2106 1393 2109 1403
rect 2138 1396 2141 1433
rect 2122 1393 2141 1396
rect 2106 1283 2109 1346
rect 2114 1323 2117 1336
rect 2066 1153 2073 1156
rect 2086 1163 2093 1166
rect 2066 1103 2069 1153
rect 2034 1073 2061 1076
rect 2026 1053 2033 1056
rect 2030 996 2033 1053
rect 2026 993 2033 996
rect 2002 913 2005 986
rect 2026 943 2029 993
rect 2018 876 2021 936
rect 2026 916 2029 936
rect 2034 923 2037 966
rect 2042 933 2045 1066
rect 2050 1003 2053 1026
rect 2058 1013 2061 1073
rect 2050 923 2053 996
rect 2026 913 2053 916
rect 2018 873 2029 876
rect 1986 833 1997 836
rect 1954 823 1989 826
rect 1994 806 1997 833
rect 2002 813 2005 826
rect 1990 803 1997 806
rect 1938 783 1949 786
rect 1922 773 1933 776
rect 1910 743 1917 746
rect 1882 723 1885 736
rect 1890 733 1897 736
rect 1890 716 1893 733
rect 1882 713 1893 716
rect 1882 696 1885 713
rect 1906 706 1909 726
rect 1890 703 1909 706
rect 1882 693 1889 696
rect 1886 626 1889 693
rect 1886 623 1893 626
rect 1858 583 1861 596
rect 1850 573 1861 576
rect 1842 503 1845 526
rect 1850 493 1853 506
rect 1826 383 1837 386
rect 1802 333 1805 356
rect 1762 313 1773 316
rect 1770 256 1773 313
rect 1786 313 1805 316
rect 1770 253 1781 256
rect 1722 216 1725 236
rect 1778 223 1781 253
rect 1786 216 1789 313
rect 1810 306 1813 336
rect 1802 303 1813 306
rect 1682 203 1701 206
rect 1706 163 1709 216
rect 1722 213 1729 216
rect 1714 123 1717 186
rect 1726 136 1729 213
rect 1770 203 1773 216
rect 1778 213 1789 216
rect 1722 133 1729 136
rect 1738 133 1741 166
rect 1722 116 1725 133
rect 1666 103 1685 106
rect 1698 103 1701 116
rect 1714 113 1725 116
rect 1738 73 1741 126
rect 1778 123 1781 213
rect 1794 203 1797 236
rect 1802 213 1805 303
rect 1786 183 1789 196
rect 1786 116 1789 176
rect 1754 113 1789 116
rect 1794 83 1797 126
rect 1802 103 1805 206
rect 1826 186 1829 383
rect 1842 233 1845 406
rect 1850 303 1853 406
rect 1858 333 1861 573
rect 1874 556 1877 616
rect 1882 593 1885 606
rect 1890 603 1893 623
rect 1898 613 1901 646
rect 1866 553 1877 556
rect 1866 513 1869 553
rect 1906 546 1909 696
rect 1874 543 1909 546
rect 1874 513 1877 543
rect 1914 536 1917 743
rect 1922 613 1925 773
rect 1946 736 1949 783
rect 1938 733 1949 736
rect 1938 636 1941 733
rect 1970 723 1973 766
rect 1978 716 1981 736
rect 1962 713 1981 716
rect 1962 646 1965 713
rect 1962 643 1973 646
rect 1930 633 1941 636
rect 1882 533 1917 536
rect 1882 453 1885 533
rect 1866 386 1869 426
rect 1882 406 1885 416
rect 1890 406 1893 526
rect 1882 403 1893 406
rect 1898 403 1901 516
rect 1914 506 1917 526
rect 1910 503 1917 506
rect 1910 436 1913 503
rect 1906 433 1913 436
rect 1866 383 1877 386
rect 1874 326 1877 383
rect 1866 323 1877 326
rect 1850 213 1853 256
rect 1866 213 1869 323
rect 1882 213 1885 226
rect 1826 183 1837 186
rect 1826 143 1829 166
rect 1834 133 1837 183
rect 1850 133 1853 176
rect 1858 166 1861 206
rect 1866 203 1877 206
rect 1890 203 1893 403
rect 1898 303 1901 316
rect 1906 283 1909 433
rect 1914 406 1917 426
rect 1922 413 1925 516
rect 1930 423 1933 633
rect 1938 623 1949 626
rect 1946 523 1949 606
rect 1954 603 1957 616
rect 1970 606 1973 643
rect 1978 616 1981 706
rect 1990 686 1993 803
rect 1990 683 1997 686
rect 1986 623 1989 666
rect 1978 613 1989 616
rect 1970 603 1981 606
rect 1986 603 1989 613
rect 1954 533 1957 596
rect 1962 543 1973 546
rect 1962 516 1965 526
rect 1978 523 1981 603
rect 1938 513 1965 516
rect 1938 496 1941 513
rect 1938 493 1945 496
rect 1942 426 1945 493
rect 1938 423 1945 426
rect 1914 403 1925 406
rect 1914 316 1917 336
rect 1922 323 1925 403
rect 1930 323 1933 336
rect 1938 323 1941 423
rect 1954 413 1957 476
rect 1946 336 1949 406
rect 1946 333 1957 336
rect 1962 333 1965 436
rect 1970 413 1973 486
rect 1986 396 1989 416
rect 1978 393 1989 396
rect 1978 346 1981 393
rect 1978 343 1989 346
rect 1994 343 1997 683
rect 2002 653 2005 796
rect 2010 696 2013 806
rect 2018 713 2021 806
rect 2026 723 2029 873
rect 2042 826 2045 866
rect 2050 833 2053 913
rect 2058 843 2061 1006
rect 2034 803 2037 826
rect 2042 823 2061 826
rect 2058 813 2061 823
rect 2050 803 2061 806
rect 2066 803 2069 1026
rect 2074 963 2077 1136
rect 2086 1106 2089 1163
rect 2098 1113 2101 1186
rect 2106 1123 2109 1206
rect 2086 1103 2093 1106
rect 2074 823 2077 936
rect 2082 933 2085 1016
rect 2090 926 2093 1103
rect 2114 1096 2117 1316
rect 2106 1093 2117 1096
rect 2106 1026 2109 1093
rect 2106 1023 2117 1026
rect 2082 923 2093 926
rect 2098 1003 2109 1006
rect 2098 923 2101 1003
rect 2106 933 2109 946
rect 2082 883 2085 923
rect 2090 886 2093 906
rect 2090 883 2101 886
rect 2082 783 2085 846
rect 2098 826 2101 883
rect 2094 823 2101 826
rect 2074 733 2085 736
rect 2074 713 2077 733
rect 2094 726 2097 823
rect 2090 723 2097 726
rect 2010 693 2017 696
rect 2002 613 2005 646
rect 2014 596 2017 693
rect 2026 636 2029 706
rect 2034 643 2037 706
rect 2026 633 2045 636
rect 2042 623 2045 633
rect 2050 616 2053 706
rect 2082 703 2085 716
rect 2026 613 2053 616
rect 2014 593 2021 596
rect 2010 523 2013 536
rect 2018 506 2021 593
rect 2026 533 2029 613
rect 2026 513 2029 526
rect 2010 503 2021 506
rect 2002 386 2005 406
rect 2010 403 2013 503
rect 2026 403 2029 466
rect 2002 383 2009 386
rect 1946 316 1949 326
rect 1914 313 1949 316
rect 1898 183 1901 216
rect 1858 163 1901 166
rect 1858 123 1861 146
rect 1898 133 1901 163
rect 1898 116 1901 126
rect 1906 123 1909 176
rect 1946 133 1949 146
rect 1914 116 1917 126
rect 1898 113 1917 116
rect 1954 73 1957 333
rect 1986 313 1989 343
rect 2006 336 2009 383
rect 2034 373 2037 606
rect 2050 593 2053 613
rect 2058 586 2061 696
rect 2054 583 2061 586
rect 2042 493 2045 536
rect 2054 486 2057 583
rect 2050 483 2057 486
rect 2050 426 2053 483
rect 2046 423 2053 426
rect 2046 356 2049 423
rect 2002 333 2009 336
rect 1978 213 1981 306
rect 2002 213 2005 333
rect 2018 323 2021 356
rect 2046 353 2053 356
rect 2026 326 2029 336
rect 2034 333 2037 346
rect 2050 336 2053 353
rect 2058 346 2061 416
rect 2066 376 2069 606
rect 2074 506 2077 656
rect 2090 616 2093 723
rect 2106 706 2109 806
rect 2114 723 2117 1023
rect 2098 703 2109 706
rect 2098 623 2101 703
rect 2090 613 2101 616
rect 2082 543 2085 606
rect 2106 583 2109 606
rect 2082 513 2085 526
rect 2074 503 2085 506
rect 2074 403 2077 426
rect 2082 413 2085 503
rect 2090 433 2093 576
rect 2114 546 2117 646
rect 2106 543 2117 546
rect 2106 386 2109 543
rect 2114 523 2117 536
rect 2122 506 2125 1393
rect 2146 1346 2149 1556
rect 2130 1343 2149 1346
rect 2130 1323 2133 1343
rect 2138 1323 2141 1336
rect 2146 1303 2149 1326
rect 2154 1313 2157 1613
rect 2162 1573 2165 1616
rect 2162 1443 2165 1556
rect 2130 1203 2133 1226
rect 2130 1123 2133 1146
rect 2130 1103 2133 1116
rect 2138 1036 2141 1296
rect 2146 1213 2149 1226
rect 2162 1213 2165 1426
rect 2170 1236 2173 1536
rect 2178 1503 2181 1526
rect 2186 1523 2189 1636
rect 2194 1506 2197 1716
rect 2190 1503 2197 1506
rect 2178 1303 2181 1446
rect 2190 1406 2193 1503
rect 2186 1403 2193 1406
rect 2186 1393 2189 1403
rect 2178 1243 2181 1286
rect 2186 1243 2189 1336
rect 2194 1323 2197 1396
rect 2202 1346 2205 1966
rect 2210 1923 2213 1973
rect 2218 1903 2221 1983
rect 2226 1886 2229 2036
rect 2234 2023 2237 2106
rect 2246 2046 2249 2113
rect 2266 2106 2269 2316
rect 2274 2223 2277 2236
rect 2274 2203 2277 2216
rect 2274 2123 2277 2146
rect 2266 2103 2273 2106
rect 2246 2043 2253 2046
rect 2242 2013 2245 2026
rect 2242 1976 2245 2006
rect 2234 1973 2245 1976
rect 2234 1923 2237 1973
rect 2250 1966 2253 2043
rect 2242 1963 2253 1966
rect 2242 1933 2245 1963
rect 2258 1916 2261 2086
rect 2270 2036 2273 2103
rect 2282 2073 2285 2326
rect 2306 2323 2309 2393
rect 2322 2333 2325 2416
rect 2370 2413 2373 2453
rect 2418 2436 2421 2493
rect 2386 2403 2389 2436
rect 2418 2433 2429 2436
rect 2354 2313 2357 2386
rect 2362 2333 2381 2336
rect 2250 1913 2261 1916
rect 2266 2033 2273 2036
rect 2214 1883 2229 1886
rect 2214 1786 2217 1883
rect 2210 1783 2217 1786
rect 2210 1683 2213 1783
rect 2218 1653 2221 1766
rect 2226 1743 2229 1856
rect 2226 1703 2229 1726
rect 2234 1646 2237 1886
rect 2242 1813 2245 1826
rect 2242 1733 2245 1756
rect 2250 1713 2253 1913
rect 2258 1706 2261 1906
rect 2210 1623 2213 1636
rect 2210 1603 2213 1616
rect 2210 1583 2213 1596
rect 2210 1503 2213 1536
rect 2218 1533 2221 1646
rect 2226 1643 2237 1646
rect 2226 1616 2229 1643
rect 2242 1633 2245 1706
rect 2250 1703 2261 1706
rect 2234 1623 2245 1626
rect 2250 1623 2253 1703
rect 2226 1613 2237 1616
rect 2258 1613 2261 1686
rect 2234 1586 2237 1613
rect 2226 1523 2229 1586
rect 2234 1583 2245 1586
rect 2234 1533 2237 1583
rect 2250 1536 2253 1606
rect 2258 1543 2261 1606
rect 2250 1533 2261 1536
rect 2242 1523 2253 1526
rect 2242 1516 2245 1523
rect 2226 1513 2245 1516
rect 2258 1496 2261 1533
rect 2250 1493 2261 1496
rect 2210 1373 2213 1416
rect 2218 1396 2221 1476
rect 2226 1403 2229 1456
rect 2250 1426 2253 1493
rect 2218 1393 2229 1396
rect 2202 1343 2221 1346
rect 2202 1323 2213 1326
rect 2170 1233 2181 1236
rect 2154 1156 2157 1206
rect 2170 1203 2173 1226
rect 2146 1153 2157 1156
rect 2130 1033 2141 1036
rect 2130 903 2133 1033
rect 2138 963 2141 1026
rect 2146 923 2149 1056
rect 2154 926 2157 1146
rect 2162 933 2165 1136
rect 2170 1033 2173 1186
rect 2178 1123 2181 1233
rect 2186 1153 2189 1216
rect 2178 1103 2181 1116
rect 2170 996 2173 1026
rect 2186 1023 2189 1126
rect 2194 1016 2197 1316
rect 2202 1116 2205 1296
rect 2218 1283 2221 1343
rect 2226 1323 2229 1393
rect 2234 1313 2237 1426
rect 2250 1423 2261 1426
rect 2242 1373 2245 1406
rect 2242 1323 2245 1336
rect 2210 1143 2213 1226
rect 2202 1113 2209 1116
rect 2206 1046 2209 1113
rect 2218 1053 2221 1246
rect 2226 1203 2229 1226
rect 2234 1203 2237 1226
rect 2226 1113 2229 1146
rect 2202 1043 2209 1046
rect 2202 1023 2205 1043
rect 2178 1006 2181 1016
rect 2194 1013 2205 1016
rect 2178 1003 2189 1006
rect 2170 993 2181 996
rect 2154 923 2165 926
rect 2178 923 2181 993
rect 2186 976 2189 1003
rect 2194 986 2197 1006
rect 2202 993 2205 1013
rect 2210 1013 2221 1016
rect 2226 1013 2229 1026
rect 2210 986 2213 1013
rect 2194 983 2213 986
rect 2218 976 2221 1006
rect 2186 973 2221 976
rect 2138 823 2141 836
rect 2130 803 2141 806
rect 2146 733 2149 816
rect 2162 756 2165 923
rect 2178 826 2181 896
rect 2194 873 2197 926
rect 2202 916 2205 936
rect 2226 923 2229 936
rect 2202 913 2213 916
rect 2186 833 2197 836
rect 2178 823 2189 826
rect 2162 753 2173 756
rect 2146 723 2157 726
rect 2130 683 2133 716
rect 2146 706 2149 723
rect 2142 703 2149 706
rect 2142 636 2145 703
rect 2130 633 2145 636
rect 2130 623 2133 633
rect 2146 603 2149 626
rect 2130 543 2149 546
rect 2154 543 2157 696
rect 2162 613 2165 736
rect 2170 693 2173 753
rect 2170 623 2173 646
rect 2118 503 2125 506
rect 2118 406 2121 503
rect 2130 416 2133 526
rect 2146 523 2149 543
rect 2162 533 2173 536
rect 2154 503 2157 526
rect 2162 523 2173 526
rect 2138 423 2141 476
rect 2130 413 2141 416
rect 2146 413 2149 426
rect 2118 403 2125 406
rect 2138 403 2141 413
rect 2106 383 2113 386
rect 2066 373 2085 376
rect 2058 343 2069 346
rect 2050 333 2061 336
rect 2066 333 2069 343
rect 2026 323 2037 326
rect 2042 323 2061 326
rect 1970 173 1973 206
rect 1978 203 1989 206
rect 2002 186 2005 206
rect 2034 193 2037 323
rect 2074 313 2077 366
rect 2082 306 2085 373
rect 2098 333 2101 356
rect 2110 326 2113 383
rect 2058 303 2085 306
rect 2106 323 2113 326
rect 2058 226 2061 303
rect 2058 223 2069 226
rect 2042 186 2045 206
rect 1970 133 1973 166
rect 1978 133 1981 146
rect 1986 123 1989 186
rect 2002 183 2045 186
rect 2002 133 2005 183
rect 2026 123 2029 136
rect 2066 133 2069 223
rect 2082 213 2085 286
rect 2090 213 2093 256
rect 2082 126 2085 176
rect 2106 146 2109 323
rect 2122 203 2125 403
rect 2138 213 2141 306
rect 2146 213 2149 376
rect 2154 316 2157 416
rect 2162 403 2165 516
rect 2170 373 2173 523
rect 2178 483 2181 816
rect 2186 803 2189 823
rect 2186 733 2189 786
rect 2186 523 2189 726
rect 2194 603 2197 626
rect 2202 623 2205 746
rect 2202 533 2205 616
rect 2194 493 2197 516
rect 2202 476 2205 526
rect 2210 503 2213 913
rect 2218 816 2221 886
rect 2226 833 2229 906
rect 2218 813 2225 816
rect 2222 746 2225 813
rect 2218 743 2225 746
rect 2218 533 2221 743
rect 2226 663 2229 726
rect 2234 696 2237 1156
rect 2242 1143 2245 1216
rect 2242 853 2245 1136
rect 2250 896 2253 1396
rect 2258 1323 2261 1423
rect 2266 1243 2269 2033
rect 2274 1953 2277 2016
rect 2274 1923 2277 1946
rect 2274 1883 2277 1916
rect 2282 1903 2285 1976
rect 2274 1823 2277 1856
rect 2274 1753 2277 1816
rect 2282 1803 2285 1826
rect 2290 1763 2293 2226
rect 2330 2213 2333 2236
rect 2298 1973 2301 2126
rect 2306 2103 2309 2206
rect 2314 2133 2317 2166
rect 2330 2146 2333 2206
rect 2338 2193 2341 2206
rect 2346 2183 2349 2216
rect 2362 2213 2365 2326
rect 2378 2296 2381 2333
rect 2386 2303 2389 2366
rect 2378 2293 2385 2296
rect 2382 2236 2385 2293
rect 2370 2223 2373 2236
rect 2382 2233 2389 2236
rect 2354 2186 2357 2206
rect 2378 2193 2381 2216
rect 2354 2183 2365 2186
rect 2330 2143 2357 2146
rect 2306 2003 2309 2016
rect 2298 1933 2301 1956
rect 2298 1913 2301 1926
rect 2306 1923 2309 1966
rect 2306 1813 2309 1886
rect 2274 1703 2277 1736
rect 2298 1723 2301 1806
rect 2282 1713 2293 1716
rect 2298 1683 2301 1716
rect 2282 1606 2285 1656
rect 2274 1603 2285 1606
rect 2274 1553 2277 1603
rect 2282 1543 2285 1566
rect 2258 1186 2261 1206
rect 2266 1203 2269 1216
rect 2274 1186 2277 1536
rect 2282 1483 2285 1536
rect 2298 1523 2301 1616
rect 2282 1413 2285 1426
rect 2290 1403 2293 1426
rect 2298 1423 2301 1436
rect 2282 1313 2285 1396
rect 2298 1393 2301 1416
rect 2290 1306 2293 1336
rect 2298 1323 2301 1336
rect 2290 1303 2297 1306
rect 2282 1216 2285 1286
rect 2294 1226 2297 1303
rect 2294 1223 2301 1226
rect 2306 1223 2309 1746
rect 2314 1243 2317 2126
rect 2322 2083 2325 2136
rect 2330 2133 2341 2136
rect 2322 2013 2325 2066
rect 2322 1946 2325 1976
rect 2330 1963 2333 2133
rect 2338 2113 2341 2126
rect 2338 1986 2341 2076
rect 2354 2073 2357 2143
rect 2362 2123 2365 2183
rect 2370 2066 2373 2166
rect 2378 2113 2381 2146
rect 2370 2063 2377 2066
rect 2346 2053 2365 2056
rect 2346 1993 2349 2053
rect 2354 2013 2357 2046
rect 2362 2013 2365 2053
rect 2374 2006 2377 2063
rect 2338 1983 2345 1986
rect 2354 1983 2357 2006
rect 2370 2003 2377 2006
rect 2322 1943 2333 1946
rect 2322 1813 2325 1866
rect 2330 1853 2333 1943
rect 2342 1886 2345 1983
rect 2342 1883 2349 1886
rect 2330 1803 2333 1826
rect 2338 1803 2341 1866
rect 2322 1306 2325 1736
rect 2338 1733 2341 1766
rect 2330 1663 2333 1726
rect 2330 1526 2333 1646
rect 2338 1603 2341 1716
rect 2338 1533 2341 1556
rect 2346 1546 2349 1883
rect 2354 1766 2357 1956
rect 2362 1883 2365 1936
rect 2362 1773 2365 1806
rect 2354 1763 2365 1766
rect 2354 1723 2357 1756
rect 2362 1713 2365 1763
rect 2370 1666 2373 2003
rect 2378 1836 2381 1946
rect 2386 1923 2389 2233
rect 2394 2123 2397 2326
rect 2410 2303 2413 2336
rect 2418 2333 2421 2356
rect 2426 2323 2429 2433
rect 2434 2376 2437 2416
rect 2434 2373 2445 2376
rect 2442 2333 2445 2373
rect 2450 2323 2453 2503
rect 2562 2503 2573 2506
rect 2594 2503 2597 2543
rect 2458 2333 2461 2426
rect 2466 2413 2469 2496
rect 2482 2403 2485 2436
rect 2506 2333 2509 2416
rect 2562 2413 2565 2503
rect 2602 2443 2605 2616
rect 2618 2546 2621 2703
rect 2626 2603 2629 2616
rect 2634 2613 2637 2726
rect 2682 2723 2685 2806
rect 2698 2793 2701 2823
rect 2714 2813 2725 2816
rect 2730 2813 2733 2823
rect 2714 2766 2717 2806
rect 2722 2793 2725 2806
rect 2746 2803 2749 2823
rect 2714 2763 2721 2766
rect 2690 2603 2693 2756
rect 2718 2686 2721 2763
rect 2754 2756 2757 2943
rect 2762 2803 2765 3006
rect 2834 3003 2837 3023
rect 2794 2923 2797 2946
rect 2818 2933 2821 2956
rect 2834 2866 2837 2886
rect 2810 2863 2837 2866
rect 2794 2826 2797 2846
rect 2786 2823 2797 2826
rect 2786 2776 2789 2823
rect 2786 2773 2797 2776
rect 2746 2753 2757 2756
rect 2714 2683 2721 2686
rect 2714 2613 2717 2683
rect 2730 2633 2733 2726
rect 2746 2706 2749 2753
rect 2770 2733 2773 2756
rect 2746 2703 2757 2706
rect 2610 2543 2621 2546
rect 2610 2486 2613 2543
rect 2618 2503 2621 2536
rect 2626 2513 2629 2526
rect 2642 2523 2645 2536
rect 2690 2513 2693 2526
rect 2610 2483 2617 2486
rect 2578 2403 2581 2436
rect 2538 2333 2549 2336
rect 2442 2283 2445 2316
rect 2490 2296 2493 2326
rect 2506 2303 2509 2316
rect 2490 2293 2501 2296
rect 2402 2116 2405 2226
rect 2418 2146 2421 2206
rect 2434 2203 2437 2226
rect 2442 2213 2445 2226
rect 2442 2193 2445 2206
rect 2410 2133 2413 2146
rect 2418 2143 2437 2146
rect 2398 2113 2405 2116
rect 2398 2046 2401 2113
rect 2394 2043 2401 2046
rect 2386 1903 2389 1916
rect 2378 1833 2389 1836
rect 2378 1703 2381 1826
rect 2386 1696 2389 1833
rect 2394 1743 2397 2043
rect 2410 2033 2413 2046
rect 2402 1973 2405 2026
rect 2410 1943 2413 2016
rect 2402 1763 2405 1936
rect 2410 1903 2413 1926
rect 2410 1803 2413 1826
rect 2394 1733 2405 1736
rect 2410 1733 2413 1756
rect 2402 1713 2405 1726
rect 2386 1693 2397 1696
rect 2354 1663 2373 1666
rect 2354 1563 2357 1663
rect 2362 1653 2381 1656
rect 2362 1633 2365 1653
rect 2362 1603 2365 1616
rect 2370 1566 2373 1636
rect 2378 1623 2381 1653
rect 2362 1563 2373 1566
rect 2346 1543 2353 1546
rect 2330 1523 2341 1526
rect 2330 1393 2333 1516
rect 2338 1423 2341 1523
rect 2350 1426 2353 1543
rect 2362 1493 2365 1563
rect 2370 1533 2373 1546
rect 2378 1533 2381 1596
rect 2394 1586 2397 1693
rect 2410 1633 2413 1646
rect 2386 1583 2397 1586
rect 2386 1526 2389 1583
rect 2410 1566 2413 1626
rect 2370 1523 2389 1526
rect 2394 1563 2413 1566
rect 2370 1436 2373 1523
rect 2346 1423 2353 1426
rect 2366 1433 2373 1436
rect 2346 1386 2349 1423
rect 2330 1383 2349 1386
rect 2330 1323 2333 1383
rect 2354 1333 2357 1406
rect 2366 1356 2369 1433
rect 2366 1353 2373 1356
rect 2322 1303 2329 1306
rect 2326 1236 2329 1303
rect 2322 1233 2329 1236
rect 2298 1216 2301 1223
rect 2282 1213 2293 1216
rect 2298 1213 2309 1216
rect 2258 1183 2277 1186
rect 2258 1123 2261 1176
rect 2266 1123 2269 1183
rect 2282 1103 2285 1206
rect 2258 1013 2261 1076
rect 2274 1003 2277 1056
rect 2290 1036 2293 1213
rect 2298 1156 2301 1206
rect 2306 1183 2309 1213
rect 2298 1153 2309 1156
rect 2298 1133 2301 1146
rect 2286 1033 2293 1036
rect 2258 913 2261 926
rect 2266 923 2269 946
rect 2250 893 2257 896
rect 2242 813 2245 836
rect 2254 826 2257 893
rect 2250 823 2257 826
rect 2266 823 2269 906
rect 2242 733 2245 806
rect 2250 796 2253 823
rect 2258 803 2269 806
rect 2250 793 2261 796
rect 2250 713 2253 786
rect 2234 693 2245 696
rect 2242 636 2245 693
rect 2242 633 2253 636
rect 2234 593 2237 616
rect 2242 573 2245 606
rect 2250 566 2253 633
rect 2258 583 2261 793
rect 2266 753 2269 786
rect 2274 753 2277 936
rect 2286 876 2289 1033
rect 2286 873 2293 876
rect 2266 733 2269 746
rect 2266 576 2269 726
rect 2274 696 2277 726
rect 2282 713 2285 856
rect 2274 693 2281 696
rect 2278 626 2281 693
rect 2290 663 2293 873
rect 2298 826 2301 1026
rect 2306 956 2309 1153
rect 2314 1113 2317 1146
rect 2314 1003 2317 1056
rect 2306 953 2317 956
rect 2306 933 2309 946
rect 2306 883 2309 916
rect 2314 833 2317 953
rect 2298 823 2317 826
rect 2298 736 2301 786
rect 2306 743 2309 816
rect 2314 736 2317 823
rect 2322 743 2325 1233
rect 2338 1213 2341 1226
rect 2330 1203 2341 1206
rect 2346 1196 2349 1316
rect 2362 1276 2365 1336
rect 2354 1273 2365 1276
rect 2354 1223 2357 1273
rect 2330 1193 2349 1196
rect 2330 1106 2333 1193
rect 2338 1183 2349 1186
rect 2338 1123 2341 1156
rect 2330 1103 2337 1106
rect 2334 1026 2337 1103
rect 2330 1023 2337 1026
rect 2330 906 2333 1023
rect 2338 916 2341 1006
rect 2346 983 2349 1183
rect 2354 1143 2357 1206
rect 2354 1013 2357 1116
rect 2354 963 2357 1006
rect 2354 923 2357 946
rect 2362 943 2365 1246
rect 2362 923 2365 936
rect 2370 933 2373 1353
rect 2378 1343 2381 1426
rect 2378 1323 2381 1336
rect 2378 1213 2381 1316
rect 2386 1296 2389 1476
rect 2394 1403 2397 1563
rect 2402 1503 2405 1516
rect 2410 1496 2413 1556
rect 2418 1516 2421 2136
rect 2426 2023 2429 2106
rect 2426 1933 2429 2016
rect 2426 1863 2429 1926
rect 2426 1803 2429 1826
rect 2434 1823 2437 2143
rect 2442 2133 2445 2166
rect 2442 2103 2445 2116
rect 2434 1773 2437 1816
rect 2426 1713 2429 1736
rect 2434 1683 2437 1726
rect 2426 1543 2429 1636
rect 2418 1513 2429 1516
rect 2410 1493 2417 1496
rect 2414 1436 2417 1493
rect 2426 1463 2429 1513
rect 2414 1433 2421 1436
rect 2418 1413 2421 1433
rect 2434 1413 2437 1646
rect 2442 1613 2445 2046
rect 2450 1976 2453 2206
rect 2474 2196 2477 2246
rect 2498 2226 2501 2293
rect 2482 2203 2485 2226
rect 2498 2223 2505 2226
rect 2474 2193 2485 2196
rect 2458 2133 2469 2136
rect 2458 2113 2461 2126
rect 2450 1973 2461 1976
rect 2450 1903 2453 1966
rect 2450 1763 2453 1826
rect 2458 1816 2461 1973
rect 2466 1943 2469 2046
rect 2466 1923 2469 1936
rect 2474 1916 2477 2136
rect 2482 2103 2485 2193
rect 2482 2013 2485 2026
rect 2482 1933 2485 1946
rect 2490 1933 2493 2216
rect 2502 2146 2505 2223
rect 2498 2143 2505 2146
rect 2498 2123 2501 2143
rect 2498 2013 2501 2066
rect 2506 2003 2509 2016
rect 2490 1923 2501 1926
rect 2506 1923 2509 1976
rect 2498 1916 2501 1923
rect 2514 1916 2517 2236
rect 2530 2213 2533 2326
rect 2562 2313 2565 2366
rect 2586 2303 2589 2336
rect 2594 2286 2597 2376
rect 2602 2333 2605 2426
rect 2614 2346 2617 2483
rect 2610 2343 2617 2346
rect 2586 2283 2597 2286
rect 2610 2286 2613 2343
rect 2626 2333 2629 2416
rect 2658 2413 2661 2446
rect 2674 2403 2677 2436
rect 2634 2323 2637 2346
rect 2626 2303 2629 2316
rect 2610 2283 2621 2286
rect 2538 2223 2541 2236
rect 2538 2206 2541 2216
rect 2562 2213 2565 2226
rect 2522 2203 2541 2206
rect 2546 2203 2565 2206
rect 2522 2126 2525 2146
rect 2522 2123 2529 2126
rect 2526 2026 2529 2123
rect 2526 2023 2533 2026
rect 2522 1993 2525 2006
rect 2474 1913 2489 1916
rect 2498 1913 2517 1916
rect 2522 1913 2525 1936
rect 2474 1823 2477 1906
rect 2486 1836 2489 1913
rect 2530 1906 2533 2023
rect 2538 2003 2541 2136
rect 2546 2113 2549 2166
rect 2562 2136 2565 2203
rect 2586 2166 2589 2283
rect 2602 2176 2605 2256
rect 2618 2226 2621 2283
rect 2642 2236 2645 2396
rect 2650 2333 2653 2376
rect 2690 2366 2693 2386
rect 2682 2363 2693 2366
rect 2682 2296 2685 2363
rect 2698 2333 2701 2426
rect 2706 2303 2709 2596
rect 2754 2593 2757 2703
rect 2770 2566 2773 2616
rect 2778 2573 2781 2606
rect 2714 2533 2717 2546
rect 2730 2533 2733 2566
rect 2762 2563 2773 2566
rect 2762 2523 2765 2563
rect 2714 2336 2717 2416
rect 2754 2413 2757 2516
rect 2778 2513 2781 2526
rect 2770 2403 2773 2436
rect 2738 2343 2773 2346
rect 2714 2333 2725 2336
rect 2682 2293 2693 2296
rect 2690 2236 2693 2293
rect 2730 2236 2733 2326
rect 2738 2313 2741 2343
rect 2746 2326 2749 2336
rect 2770 2333 2773 2343
rect 2746 2323 2765 2326
rect 2642 2233 2653 2236
rect 2690 2233 2717 2236
rect 2730 2233 2741 2236
rect 2618 2223 2637 2226
rect 2610 2193 2613 2206
rect 2618 2183 2621 2206
rect 2602 2173 2609 2176
rect 2626 2173 2629 2216
rect 2634 2213 2637 2223
rect 2586 2163 2597 2166
rect 2562 2133 2573 2136
rect 2586 2133 2589 2146
rect 2594 2133 2597 2163
rect 2562 2123 2573 2126
rect 2578 2123 2597 2126
rect 2546 2013 2549 2056
rect 2554 2016 2557 2026
rect 2554 2013 2565 2016
rect 2554 1926 2557 2006
rect 2562 1933 2565 2013
rect 2538 1923 2565 1926
rect 2506 1903 2533 1906
rect 2538 1903 2541 1916
rect 2546 1913 2557 1916
rect 2486 1833 2493 1836
rect 2458 1813 2469 1816
rect 2474 1813 2485 1816
rect 2458 1743 2461 1806
rect 2466 1743 2469 1813
rect 2450 1733 2461 1736
rect 2450 1693 2453 1733
rect 2458 1723 2477 1726
rect 2474 1633 2477 1716
rect 2482 1626 2485 1776
rect 2450 1623 2461 1626
rect 2466 1623 2485 1626
rect 2458 1593 2461 1606
rect 2466 1576 2469 1623
rect 2442 1513 2445 1566
rect 2450 1523 2453 1576
rect 2462 1573 2469 1576
rect 2462 1516 2465 1573
rect 2474 1533 2477 1606
rect 2450 1513 2465 1516
rect 2450 1456 2453 1513
rect 2458 1483 2461 1506
rect 2474 1503 2477 1516
rect 2450 1453 2457 1456
rect 2418 1386 2421 1396
rect 2402 1383 2421 1386
rect 2402 1333 2405 1383
rect 2394 1313 2397 1326
rect 2410 1303 2413 1326
rect 2386 1293 2397 1296
rect 2418 1293 2421 1336
rect 2394 1246 2397 1293
rect 2386 1243 2397 1246
rect 2386 1223 2389 1243
rect 2386 1193 2389 1206
rect 2410 1203 2413 1286
rect 2418 1206 2421 1266
rect 2426 1216 2429 1406
rect 2434 1283 2437 1346
rect 2442 1333 2445 1446
rect 2454 1406 2457 1453
rect 2450 1403 2457 1406
rect 2474 1403 2477 1486
rect 2426 1213 2437 1216
rect 2418 1203 2429 1206
rect 2434 1203 2437 1213
rect 2442 1203 2445 1246
rect 2410 1156 2413 1196
rect 2378 1153 2413 1156
rect 2378 1106 2381 1153
rect 2386 1126 2389 1136
rect 2394 1133 2397 1146
rect 2402 1126 2405 1136
rect 2410 1133 2413 1153
rect 2426 1134 2429 1203
rect 2434 1153 2445 1156
rect 2386 1123 2413 1126
rect 2378 1103 2389 1106
rect 2386 1036 2389 1103
rect 2378 1033 2389 1036
rect 2378 956 2381 1033
rect 2386 1003 2389 1016
rect 2394 983 2397 1006
rect 2402 956 2405 1106
rect 2410 1016 2413 1123
rect 2418 1103 2421 1126
rect 2410 1013 2429 1016
rect 2410 963 2413 986
rect 2378 953 2397 956
rect 2402 953 2413 956
rect 2338 913 2349 916
rect 2330 903 2341 906
rect 2330 813 2333 896
rect 2338 786 2341 903
rect 2346 883 2349 913
rect 2378 876 2381 946
rect 2386 893 2389 926
rect 2354 873 2381 876
rect 2354 806 2357 873
rect 2394 853 2397 953
rect 2410 933 2413 953
rect 2402 806 2405 926
rect 2418 906 2421 936
rect 2410 903 2421 906
rect 2426 886 2429 966
rect 2422 883 2429 886
rect 2330 783 2341 786
rect 2346 803 2357 806
rect 2298 733 2309 736
rect 2314 733 2325 736
rect 2298 713 2301 726
rect 2314 706 2317 726
rect 2298 703 2317 706
rect 2298 653 2301 703
rect 2322 696 2325 733
rect 2306 693 2325 696
rect 2306 646 2309 693
rect 2306 643 2317 646
rect 2274 623 2281 626
rect 2274 603 2277 623
rect 2298 613 2309 616
rect 2290 603 2301 606
rect 2282 593 2293 596
rect 2234 563 2253 566
rect 2258 573 2269 576
rect 2218 493 2221 526
rect 2194 473 2205 476
rect 2162 353 2181 356
rect 2162 323 2165 353
rect 2170 316 2173 336
rect 2178 333 2181 353
rect 2154 313 2173 316
rect 2178 313 2181 326
rect 2186 323 2189 346
rect 2162 286 2165 306
rect 2162 283 2173 286
rect 2154 213 2157 226
rect 2106 143 2117 146
rect 2130 143 2133 206
rect 2146 173 2149 206
rect 2170 186 2173 283
rect 2194 213 2197 473
rect 2210 453 2221 456
rect 2210 436 2213 453
rect 2206 433 2213 436
rect 2206 326 2209 433
rect 2218 333 2221 416
rect 2226 403 2229 536
rect 2206 323 2213 326
rect 2210 203 2213 323
rect 2234 313 2237 563
rect 2242 506 2245 536
rect 2258 523 2261 573
rect 2242 503 2253 506
rect 2250 456 2253 503
rect 2242 453 2253 456
rect 2242 366 2245 453
rect 2266 426 2269 546
rect 2290 533 2293 593
rect 2274 513 2277 526
rect 2298 523 2301 603
rect 2306 593 2309 613
rect 2314 576 2317 643
rect 2310 573 2317 576
rect 2310 516 2313 573
rect 2290 513 2313 516
rect 2266 423 2277 426
rect 2250 393 2253 416
rect 2258 383 2261 406
rect 2274 376 2277 423
rect 2290 386 2293 513
rect 2306 423 2309 466
rect 2314 413 2317 426
rect 2290 383 2301 386
rect 2306 383 2309 406
rect 2266 373 2277 376
rect 2242 363 2253 366
rect 2250 306 2253 363
rect 2242 303 2253 306
rect 2162 183 2173 186
rect 2090 133 2109 136
rect 1986 103 1989 116
rect 2058 113 2061 126
rect 2082 123 2101 126
rect 2106 93 2109 116
rect 2114 53 2117 143
rect 2154 113 2157 136
rect 2162 103 2165 183
rect 2178 123 2181 166
rect 2194 123 2197 136
rect 2170 93 2173 116
rect 2210 113 2213 146
rect 2226 126 2229 216
rect 2242 213 2245 303
rect 2266 286 2269 373
rect 2298 363 2301 383
rect 2274 296 2277 316
rect 2290 313 2301 316
rect 2274 293 2285 296
rect 2258 283 2269 286
rect 2258 236 2261 283
rect 2258 233 2269 236
rect 2234 163 2237 206
rect 2226 123 2237 126
rect 2258 123 2261 206
rect 2266 126 2269 233
rect 2282 176 2285 293
rect 2298 286 2301 313
rect 2306 306 2309 326
rect 2314 316 2317 366
rect 2322 323 2325 686
rect 2330 633 2333 783
rect 2338 716 2341 756
rect 2346 723 2349 803
rect 2370 796 2373 806
rect 2378 803 2405 806
rect 2370 793 2389 796
rect 2338 713 2349 716
rect 2338 633 2341 646
rect 2330 623 2341 626
rect 2330 573 2333 616
rect 2338 583 2341 623
rect 2346 613 2349 713
rect 2354 683 2357 736
rect 2370 733 2373 766
rect 2378 726 2381 746
rect 2386 733 2389 793
rect 2394 773 2397 796
rect 2362 703 2365 726
rect 2370 723 2381 726
rect 2354 606 2357 666
rect 2370 623 2373 723
rect 2346 603 2357 606
rect 2330 413 2333 546
rect 2338 503 2341 516
rect 2314 313 2325 316
rect 2330 306 2333 316
rect 2306 303 2333 306
rect 2298 283 2309 286
rect 2298 203 2301 276
rect 2306 213 2309 283
rect 2330 223 2333 236
rect 2338 233 2341 476
rect 2282 173 2333 176
rect 2282 133 2285 166
rect 2266 123 2285 126
rect 2330 123 2333 173
rect 2202 103 2221 106
rect 2226 93 2229 116
rect 2234 43 2237 123
rect 2266 63 2269 123
rect 2338 116 2341 146
rect 2306 113 2341 116
rect 2346 83 2349 603
rect 2354 486 2357 586
rect 2362 523 2365 536
rect 2370 523 2373 546
rect 2354 483 2369 486
rect 2366 426 2369 483
rect 2378 446 2381 716
rect 2386 653 2389 726
rect 2394 673 2397 756
rect 2410 746 2413 806
rect 2422 766 2425 883
rect 2422 763 2429 766
rect 2410 743 2421 746
rect 2426 726 2429 763
rect 2434 756 2437 1126
rect 2442 1123 2445 1153
rect 2450 1106 2453 1403
rect 2466 1386 2469 1396
rect 2458 1383 2469 1386
rect 2458 1323 2461 1383
rect 2466 1356 2469 1376
rect 2466 1353 2473 1356
rect 2446 1103 2453 1106
rect 2446 1026 2449 1103
rect 2458 1053 2461 1296
rect 2470 1286 2473 1353
rect 2466 1283 2473 1286
rect 2446 1023 2453 1026
rect 2442 923 2445 1006
rect 2450 963 2453 1023
rect 2458 936 2461 1016
rect 2454 933 2461 936
rect 2442 766 2445 916
rect 2454 846 2457 933
rect 2450 843 2457 846
rect 2450 823 2453 843
rect 2458 813 2461 826
rect 2458 783 2461 806
rect 2442 763 2453 766
rect 2434 753 2445 756
rect 2402 683 2405 726
rect 2418 723 2429 726
rect 2434 723 2437 746
rect 2386 633 2389 646
rect 2418 636 2421 723
rect 2442 716 2445 753
rect 2450 743 2453 763
rect 2450 723 2453 736
rect 2434 713 2445 716
rect 2434 653 2437 713
rect 2418 633 2429 636
rect 2394 576 2397 626
rect 2402 613 2405 626
rect 2410 603 2413 616
rect 2426 583 2429 633
rect 2434 593 2437 616
rect 2442 603 2445 706
rect 2458 703 2461 766
rect 2450 613 2453 626
rect 2394 573 2413 576
rect 2386 453 2389 536
rect 2410 533 2413 573
rect 2402 503 2405 526
rect 2418 513 2421 526
rect 2378 443 2385 446
rect 2366 423 2373 426
rect 2354 303 2357 416
rect 2362 356 2365 406
rect 2370 393 2373 423
rect 2382 386 2385 443
rect 2394 423 2397 486
rect 2426 456 2429 526
rect 2458 503 2461 566
rect 2406 453 2429 456
rect 2394 393 2397 406
rect 2406 386 2409 453
rect 2382 383 2389 386
rect 2362 353 2369 356
rect 2366 296 2369 353
rect 2378 333 2381 366
rect 2386 333 2389 383
rect 2402 383 2409 386
rect 2402 336 2405 383
rect 2418 343 2421 416
rect 2394 333 2405 336
rect 2362 293 2369 296
rect 2362 233 2365 293
rect 2378 213 2381 326
rect 2394 266 2397 333
rect 2402 273 2405 326
rect 2410 313 2421 316
rect 2426 306 2429 416
rect 2434 313 2437 486
rect 2466 423 2469 1283
rect 2474 1083 2477 1266
rect 2474 983 2477 1016
rect 2474 923 2477 966
rect 2474 783 2477 866
rect 2474 713 2477 736
rect 2474 603 2477 616
rect 2474 496 2477 546
rect 2482 513 2485 1616
rect 2490 1413 2493 1833
rect 2498 1523 2501 1896
rect 2506 1573 2509 1903
rect 2514 1713 2517 1876
rect 2522 1756 2525 1896
rect 2562 1893 2565 1923
rect 2538 1823 2541 1886
rect 2546 1813 2549 1826
rect 2570 1816 2573 2006
rect 2578 1933 2581 2123
rect 2606 2116 2609 2173
rect 2634 2146 2637 2206
rect 2650 2166 2653 2233
rect 2602 2113 2609 2116
rect 2618 2143 2637 2146
rect 2642 2163 2653 2166
rect 2602 2036 2605 2113
rect 2618 2043 2621 2143
rect 2626 2103 2629 2136
rect 2634 2066 2637 2136
rect 2642 2073 2645 2163
rect 2674 2146 2677 2206
rect 2682 2193 2685 2216
rect 2690 2193 2693 2226
rect 2650 2143 2677 2146
rect 2650 2103 2653 2143
rect 2658 2113 2661 2136
rect 2666 2086 2669 2136
rect 2682 2126 2685 2176
rect 2674 2123 2685 2126
rect 2682 2113 2693 2116
rect 2698 2106 2701 2216
rect 2714 2146 2717 2233
rect 2730 2193 2733 2226
rect 2738 2203 2741 2233
rect 2762 2216 2765 2323
rect 2778 2313 2781 2366
rect 2794 2323 2797 2773
rect 2802 2723 2805 2806
rect 2810 2793 2813 2863
rect 2818 2766 2821 2836
rect 2826 2813 2829 2856
rect 2834 2813 2837 2863
rect 2842 2806 2845 3016
rect 2850 3013 2853 3023
rect 2850 2936 2853 3006
rect 2858 3003 2869 3006
rect 2874 2966 2877 3133
rect 2890 3123 2893 3136
rect 2898 3123 2901 3136
rect 2906 3113 2909 3143
rect 2890 3023 2893 3076
rect 2914 3003 2917 3136
rect 2930 3076 2933 3146
rect 2970 3133 2973 3146
rect 2926 3073 2933 3076
rect 2962 3123 2973 3126
rect 2926 3016 2929 3073
rect 2962 3066 2965 3123
rect 2922 3013 2929 3016
rect 2938 3063 2965 3066
rect 2866 2963 2877 2966
rect 2850 2933 2861 2936
rect 2826 2803 2845 2806
rect 2850 2803 2853 2926
rect 2858 2873 2861 2933
rect 2858 2813 2861 2846
rect 2866 2833 2869 2963
rect 2922 2956 2925 3013
rect 2938 3006 2941 3063
rect 2970 3016 2973 3116
rect 2978 3096 2981 3136
rect 2994 3113 2997 3153
rect 3018 3133 3021 3233
rect 3066 3213 3069 3233
rect 3090 3193 3093 3206
rect 3106 3193 3109 3206
rect 3058 3133 3061 3146
rect 3090 3126 3093 3136
rect 2978 3093 2989 3096
rect 2954 3013 2973 3016
rect 2986 3006 2989 3093
rect 2930 2996 2933 3006
rect 2938 3003 2949 3006
rect 2930 2993 2949 2996
rect 2954 2993 2957 3006
rect 2970 3003 2989 3006
rect 2906 2953 2925 2956
rect 2898 2906 2901 2926
rect 2890 2903 2901 2906
rect 2866 2803 2869 2816
rect 2874 2813 2877 2886
rect 2890 2826 2893 2903
rect 2890 2823 2901 2826
rect 2898 2806 2901 2823
rect 2874 2803 2901 2806
rect 2826 2793 2829 2803
rect 2906 2796 2909 2953
rect 2922 2933 2925 2946
rect 2946 2923 2949 2993
rect 2970 2966 2973 3003
rect 3018 2996 3021 3086
rect 3042 3023 3045 3126
rect 3058 3113 3061 3126
rect 3074 3123 3093 3126
rect 3090 3113 3093 3123
rect 3122 3116 3125 3126
rect 3130 3123 3133 3216
rect 3146 3146 3149 3206
rect 3146 3143 3157 3146
rect 3122 3113 3149 3116
rect 3066 3023 3069 3086
rect 3026 3013 3045 3016
rect 2962 2963 2973 2966
rect 2962 2886 2965 2963
rect 2962 2883 2973 2886
rect 2930 2803 2933 2846
rect 2866 2793 2909 2796
rect 2938 2793 2941 2816
rect 2818 2763 2837 2766
rect 2834 2746 2837 2763
rect 2834 2743 2841 2746
rect 2838 2686 2841 2743
rect 2866 2736 2869 2793
rect 2954 2766 2957 2816
rect 2962 2803 2965 2856
rect 2970 2806 2973 2883
rect 3002 2843 3005 2926
rect 3010 2913 3013 2996
rect 3018 2993 3025 2996
rect 3042 2993 3045 3006
rect 3022 2926 3025 2993
rect 3050 2936 3053 3006
rect 3114 2953 3117 3006
rect 3138 2993 3141 3016
rect 3154 2953 3157 3143
rect 3170 3133 3173 3216
rect 3226 3193 3229 3216
rect 3258 3153 3261 3206
rect 3234 3143 3285 3146
rect 3234 3133 3237 3143
rect 3258 3126 3261 3136
rect 3282 3133 3285 3143
rect 3194 3123 3221 3126
rect 3226 3123 3261 3126
rect 3018 2923 3025 2926
rect 3034 2923 3037 2936
rect 3050 2933 3069 2936
rect 3074 2933 3077 2946
rect 3018 2893 3021 2923
rect 3050 2913 3053 2926
rect 3058 2913 3061 2926
rect 2978 2813 3005 2816
rect 2970 2803 2981 2806
rect 2938 2763 2957 2766
rect 2862 2733 2869 2736
rect 2834 2683 2841 2686
rect 2802 2533 2805 2556
rect 2810 2503 2813 2536
rect 2818 2523 2821 2616
rect 2834 2456 2837 2683
rect 2842 2603 2845 2616
rect 2850 2523 2853 2726
rect 2862 2626 2865 2733
rect 2862 2623 2869 2626
rect 2866 2606 2869 2623
rect 2874 2613 2877 2726
rect 2890 2686 2893 2756
rect 2938 2723 2941 2763
rect 2978 2743 2981 2803
rect 2994 2793 2997 2806
rect 3002 2803 3005 2813
rect 2962 2723 2973 2726
rect 2890 2683 2901 2686
rect 2866 2603 2873 2606
rect 2898 2603 2901 2683
rect 2978 2676 2981 2736
rect 3010 2723 3013 2826
rect 3042 2813 3061 2816
rect 3042 2793 3045 2813
rect 3066 2806 3069 2933
rect 3082 2906 3085 2946
rect 3090 2933 3093 2946
rect 3146 2926 3149 2936
rect 3170 2926 3173 2946
rect 3178 2933 3181 3006
rect 3106 2913 3109 2926
rect 3138 2923 3149 2926
rect 3154 2923 3181 2926
rect 3186 2923 3189 3056
rect 3194 2983 3197 3016
rect 3194 2923 3197 2936
rect 3082 2903 3117 2906
rect 3114 2866 3117 2903
rect 3114 2863 3125 2866
rect 3050 2803 3069 2806
rect 2946 2673 2981 2676
rect 2938 2606 2941 2656
rect 2946 2613 2949 2673
rect 3018 2623 3021 2636
rect 3026 2623 3029 2636
rect 2870 2546 2873 2603
rect 2870 2543 2877 2546
rect 2834 2453 2841 2456
rect 2802 2333 2805 2426
rect 2818 2353 2821 2416
rect 2838 2376 2841 2453
rect 2850 2413 2853 2516
rect 2858 2503 2861 2526
rect 2874 2456 2877 2543
rect 2882 2533 2885 2556
rect 2930 2523 2933 2606
rect 2938 2603 2949 2606
rect 2978 2603 2981 2616
rect 2946 2533 2949 2603
rect 3034 2543 3037 2736
rect 3050 2653 3053 2736
rect 3074 2723 3077 2816
rect 3090 2813 3109 2816
rect 3082 2766 3085 2806
rect 3114 2803 3117 2856
rect 3122 2796 3125 2863
rect 3138 2806 3141 2923
rect 3154 2916 3157 2923
rect 3146 2913 3157 2916
rect 3162 2893 3165 2916
rect 3178 2846 3181 2923
rect 3178 2843 3213 2846
rect 3170 2833 3189 2836
rect 3170 2806 3173 2833
rect 3138 2803 3157 2806
rect 3098 2793 3125 2796
rect 3082 2763 3089 2766
rect 3086 2716 3089 2763
rect 3082 2713 3089 2716
rect 3058 2646 3061 2686
rect 3042 2643 3061 2646
rect 3042 2633 3045 2643
rect 3050 2543 3053 2626
rect 3058 2623 3061 2636
rect 3082 2613 3085 2713
rect 3098 2613 3101 2793
rect 3138 2706 3141 2726
rect 3130 2703 3141 2706
rect 3074 2533 3077 2546
rect 3082 2533 3101 2536
rect 3082 2526 3085 2533
rect 2874 2453 2909 2456
rect 2866 2403 2869 2436
rect 2834 2373 2841 2376
rect 2834 2326 2837 2373
rect 2842 2333 2845 2356
rect 2850 2333 2853 2376
rect 2890 2333 2893 2416
rect 2906 2396 2909 2453
rect 2946 2413 2949 2526
rect 2962 2403 2965 2426
rect 2898 2393 2909 2396
rect 2898 2373 2901 2393
rect 2826 2306 2829 2326
rect 2834 2323 2845 2326
rect 2786 2223 2789 2236
rect 2746 2156 2749 2216
rect 2762 2213 2789 2216
rect 2794 2213 2797 2266
rect 2754 2173 2757 2206
rect 2730 2153 2749 2156
rect 2714 2143 2721 2146
rect 2658 2083 2669 2086
rect 2634 2063 2645 2066
rect 2642 2046 2645 2063
rect 2642 2043 2649 2046
rect 2602 2033 2629 2036
rect 2586 2013 2589 2026
rect 2594 2003 2597 2016
rect 2602 2013 2605 2026
rect 2578 1873 2581 1926
rect 2586 1826 2589 1926
rect 2602 1916 2605 1986
rect 2610 1923 2613 1936
rect 2602 1913 2613 1916
rect 2610 1896 2613 1913
rect 2606 1893 2613 1896
rect 2578 1823 2589 1826
rect 2594 1823 2597 1846
rect 2606 1836 2609 1893
rect 2606 1833 2613 1836
rect 2570 1813 2601 1816
rect 2554 1803 2589 1806
rect 2562 1793 2573 1796
rect 2522 1753 2533 1756
rect 2514 1693 2517 1706
rect 2514 1613 2517 1626
rect 2522 1613 2525 1746
rect 2522 1536 2525 1606
rect 2506 1533 2525 1536
rect 2498 1406 2501 1466
rect 2490 1403 2501 1406
rect 2490 1323 2493 1403
rect 2498 1373 2501 1396
rect 2506 1346 2509 1533
rect 2498 1343 2509 1346
rect 2490 1213 2493 1246
rect 2498 1186 2501 1343
rect 2514 1336 2517 1526
rect 2522 1433 2525 1516
rect 2530 1506 2533 1753
rect 2538 1596 2541 1746
rect 2546 1606 2549 1776
rect 2554 1693 2557 1716
rect 2554 1623 2557 1666
rect 2562 1653 2565 1793
rect 2586 1733 2589 1803
rect 2598 1746 2601 1813
rect 2598 1743 2605 1746
rect 2570 1723 2597 1726
rect 2570 1713 2589 1716
rect 2570 1693 2573 1713
rect 2594 1706 2597 1723
rect 2546 1603 2557 1606
rect 2538 1593 2549 1596
rect 2538 1523 2541 1586
rect 2530 1503 2537 1506
rect 2534 1436 2537 1503
rect 2530 1433 2537 1436
rect 2522 1413 2525 1426
rect 2506 1333 2517 1336
rect 2522 1333 2525 1376
rect 2530 1346 2533 1433
rect 2538 1356 2541 1416
rect 2546 1403 2549 1593
rect 2554 1543 2557 1603
rect 2538 1353 2549 1356
rect 2530 1343 2549 1346
rect 2530 1333 2541 1336
rect 2506 1316 2509 1333
rect 2514 1323 2525 1326
rect 2506 1313 2517 1316
rect 2522 1313 2525 1323
rect 2506 1193 2509 1256
rect 2514 1193 2517 1313
rect 2530 1303 2533 1326
rect 2546 1276 2549 1343
rect 2530 1273 2549 1276
rect 2522 1213 2525 1246
rect 2522 1186 2525 1206
rect 2498 1183 2525 1186
rect 2490 1103 2493 1136
rect 2498 1133 2509 1136
rect 2498 1123 2501 1133
rect 2490 906 2493 1056
rect 2498 1013 2501 1076
rect 2498 983 2501 1006
rect 2506 996 2509 1126
rect 2514 1073 2517 1183
rect 2522 1113 2525 1126
rect 2530 1096 2533 1273
rect 2526 1093 2533 1096
rect 2526 1026 2529 1093
rect 2526 1023 2533 1026
rect 2514 1003 2525 1006
rect 2506 993 2517 996
rect 2498 933 2501 946
rect 2506 923 2509 936
rect 2514 933 2517 993
rect 2530 986 2533 1023
rect 2538 1013 2541 1256
rect 2546 1113 2549 1186
rect 2526 983 2533 986
rect 2526 916 2529 983
rect 2538 973 2541 1006
rect 2546 963 2549 1026
rect 2546 933 2549 946
rect 2538 923 2549 926
rect 2526 913 2533 916
rect 2490 903 2497 906
rect 2494 846 2497 903
rect 2494 843 2501 846
rect 2490 733 2493 836
rect 2490 653 2493 726
rect 2498 693 2501 843
rect 2506 753 2509 856
rect 2530 816 2533 913
rect 2546 856 2549 923
rect 2538 853 2549 856
rect 2538 823 2541 853
rect 2530 813 2541 816
rect 2506 646 2509 746
rect 2514 703 2517 716
rect 2522 663 2525 806
rect 2490 643 2509 646
rect 2490 616 2493 643
rect 2498 623 2525 626
rect 2490 613 2501 616
rect 2522 613 2525 623
rect 2490 536 2493 606
rect 2498 543 2501 613
rect 2490 533 2525 536
rect 2474 493 2481 496
rect 2490 493 2493 526
rect 2498 513 2509 516
rect 2478 426 2481 493
rect 2478 423 2485 426
rect 2442 403 2469 406
rect 2442 383 2445 403
rect 2474 373 2477 416
rect 2418 303 2429 306
rect 2394 263 2413 266
rect 2386 233 2405 236
rect 2394 206 2397 226
rect 2362 203 2397 206
rect 2410 203 2413 263
rect 2362 123 2365 203
rect 2402 76 2405 136
rect 2410 113 2413 126
rect 2418 83 2421 303
rect 2442 253 2445 326
rect 2466 316 2469 336
rect 2458 313 2469 316
rect 2458 236 2461 313
rect 2426 223 2429 236
rect 2458 233 2469 236
rect 2442 203 2445 216
rect 2466 213 2469 233
rect 2474 196 2477 336
rect 2482 323 2485 423
rect 2490 316 2493 486
rect 2498 333 2501 426
rect 2506 333 2509 346
rect 2486 313 2493 316
rect 2498 313 2501 326
rect 2486 246 2489 313
rect 2466 193 2477 196
rect 2482 243 2489 246
rect 2466 146 2469 193
rect 2426 76 2429 136
rect 2434 123 2437 146
rect 2466 143 2477 146
rect 2474 123 2477 143
rect 2482 133 2485 243
rect 2490 203 2493 226
rect 2506 213 2509 306
rect 2514 233 2517 326
rect 2522 323 2525 533
rect 2530 513 2533 736
rect 2538 733 2541 813
rect 2546 733 2549 816
rect 2538 633 2541 726
rect 2554 716 2557 1536
rect 2562 1413 2565 1606
rect 2570 1533 2573 1686
rect 2570 1513 2573 1526
rect 2570 1493 2573 1506
rect 2562 1373 2565 1396
rect 2570 1393 2573 1416
rect 2578 1386 2581 1706
rect 2590 1703 2597 1706
rect 2602 1703 2605 1743
rect 2590 1636 2593 1703
rect 2586 1633 2593 1636
rect 2586 1616 2589 1633
rect 2586 1613 2605 1616
rect 2602 1593 2605 1606
rect 2586 1513 2589 1546
rect 2602 1533 2605 1546
rect 2570 1383 2581 1386
rect 2586 1383 2589 1416
rect 2562 1213 2565 1336
rect 2570 1213 2573 1383
rect 2578 1353 2581 1376
rect 2578 1313 2581 1326
rect 2578 1166 2581 1226
rect 2586 1203 2589 1326
rect 2594 1323 2597 1526
rect 2602 1343 2605 1516
rect 2602 1273 2605 1336
rect 2610 1256 2613 1833
rect 2618 1803 2621 2006
rect 2626 1843 2629 2033
rect 2626 1736 2629 1826
rect 2618 1733 2629 1736
rect 2618 1693 2621 1733
rect 2626 1683 2629 1726
rect 2634 1676 2637 2016
rect 2646 1966 2649 2043
rect 2642 1963 2649 1966
rect 2642 1773 2645 1963
rect 2650 1776 2653 1946
rect 2658 1823 2661 2083
rect 2674 2016 2677 2106
rect 2666 2013 2677 2016
rect 2682 2103 2701 2106
rect 2682 2013 2685 2103
rect 2698 2013 2701 2066
rect 2666 1896 2669 2013
rect 2674 1983 2677 2006
rect 2706 1973 2709 2126
rect 2718 2056 2721 2143
rect 2730 2066 2733 2153
rect 2738 2143 2773 2146
rect 2738 2133 2741 2143
rect 2746 2066 2749 2136
rect 2754 2113 2757 2126
rect 2762 2123 2765 2136
rect 2770 2123 2773 2143
rect 2794 2136 2797 2146
rect 2778 2133 2797 2136
rect 2778 2093 2781 2126
rect 2802 2113 2805 2236
rect 2810 2096 2813 2306
rect 2826 2303 2837 2306
rect 2834 2206 2837 2303
rect 2858 2223 2861 2316
rect 2866 2213 2869 2236
rect 2818 2183 2821 2206
rect 2826 2203 2837 2206
rect 2802 2093 2813 2096
rect 2730 2063 2741 2066
rect 2746 2063 2765 2066
rect 2718 2053 2725 2056
rect 2674 1923 2701 1926
rect 2690 1903 2693 1916
rect 2666 1893 2677 1896
rect 2674 1846 2677 1893
rect 2666 1843 2677 1846
rect 2666 1826 2669 1843
rect 2666 1823 2709 1826
rect 2714 1816 2717 2006
rect 2722 1996 2725 2053
rect 2738 2013 2741 2063
rect 2746 1996 2749 2046
rect 2762 2016 2765 2063
rect 2802 2036 2805 2093
rect 2770 2023 2773 2036
rect 2802 2033 2813 2036
rect 2722 1993 2733 1996
rect 2650 1773 2661 1776
rect 2650 1713 2653 1746
rect 2650 1683 2653 1706
rect 2658 1703 2661 1726
rect 2634 1673 2645 1676
rect 2618 1403 2621 1646
rect 2626 1613 2629 1626
rect 2626 1573 2629 1606
rect 2626 1523 2629 1566
rect 2634 1533 2637 1666
rect 2642 1516 2645 1673
rect 2650 1623 2653 1646
rect 2658 1643 2661 1656
rect 2666 1636 2669 1816
rect 2658 1633 2669 1636
rect 2674 1813 2717 1816
rect 2650 1533 2653 1546
rect 2658 1536 2661 1633
rect 2666 1563 2669 1626
rect 2674 1623 2677 1813
rect 2682 1796 2685 1806
rect 2722 1803 2725 1886
rect 2730 1813 2733 1993
rect 2742 1993 2749 1996
rect 2742 1926 2745 1993
rect 2754 1936 2757 2016
rect 2762 2013 2773 2016
rect 2810 2013 2813 2033
rect 2770 2003 2773 2013
rect 2818 2006 2821 2126
rect 2826 2013 2829 2203
rect 2754 1933 2789 1936
rect 2742 1923 2749 1926
rect 2682 1793 2733 1796
rect 2682 1713 2685 1766
rect 2690 1673 2693 1776
rect 2674 1573 2677 1616
rect 2682 1606 2685 1636
rect 2690 1613 2693 1626
rect 2682 1603 2701 1606
rect 2658 1533 2689 1536
rect 2626 1413 2629 1516
rect 2638 1513 2645 1516
rect 2638 1436 2641 1513
rect 2638 1433 2645 1436
rect 2618 1373 2621 1396
rect 2634 1383 2637 1416
rect 2618 1333 2621 1366
rect 2606 1253 2613 1256
rect 2594 1173 2597 1216
rect 2606 1206 2609 1253
rect 2618 1213 2621 1306
rect 2626 1296 2629 1356
rect 2634 1333 2637 1346
rect 2634 1313 2637 1326
rect 2626 1293 2633 1296
rect 2630 1206 2633 1293
rect 2606 1203 2613 1206
rect 2562 1163 2581 1166
rect 2562 793 2565 1163
rect 2570 1023 2573 1156
rect 2610 1133 2613 1203
rect 2626 1203 2633 1206
rect 2626 1136 2629 1203
rect 2570 993 2573 1016
rect 2570 893 2573 986
rect 2578 953 2581 1036
rect 2578 933 2581 946
rect 2578 896 2581 926
rect 2586 923 2589 1126
rect 2594 1083 2597 1126
rect 2602 1123 2613 1126
rect 2618 1103 2621 1136
rect 2626 1133 2637 1136
rect 2594 916 2597 1076
rect 2610 1016 2613 1076
rect 2626 1053 2629 1126
rect 2606 1013 2613 1016
rect 2606 946 2609 1013
rect 2618 993 2621 1036
rect 2626 1006 2629 1026
rect 2634 1013 2637 1133
rect 2626 1003 2637 1006
rect 2642 986 2645 1433
rect 2650 1396 2653 1526
rect 2658 1483 2661 1526
rect 2666 1513 2677 1516
rect 2658 1406 2661 1456
rect 2666 1413 2669 1513
rect 2658 1403 2669 1406
rect 2674 1403 2677 1436
rect 2686 1406 2689 1533
rect 2682 1403 2689 1406
rect 2650 1393 2661 1396
rect 2650 1173 2653 1386
rect 2658 1253 2661 1393
rect 2666 1246 2669 1403
rect 2674 1333 2677 1346
rect 2682 1326 2685 1403
rect 2690 1343 2693 1396
rect 2674 1323 2685 1326
rect 2690 1313 2693 1326
rect 2658 1243 2669 1246
rect 2650 1073 2653 1136
rect 2602 943 2609 946
rect 2602 923 2605 943
rect 2618 933 2621 986
rect 2638 983 2645 986
rect 2610 923 2621 926
rect 2594 913 2601 916
rect 2578 893 2589 896
rect 2562 733 2565 746
rect 2554 713 2561 716
rect 2538 533 2541 576
rect 2530 216 2533 456
rect 2538 413 2541 436
rect 2538 306 2541 406
rect 2546 333 2549 696
rect 2558 646 2561 713
rect 2554 643 2561 646
rect 2554 413 2557 643
rect 2562 523 2565 626
rect 2570 546 2573 876
rect 2586 826 2589 893
rect 2578 823 2589 826
rect 2598 826 2601 913
rect 2618 893 2621 923
rect 2626 903 2629 926
rect 2638 886 2641 983
rect 2650 943 2653 1016
rect 2658 936 2661 1243
rect 2666 1203 2669 1216
rect 2666 1123 2669 1136
rect 2674 1106 2677 1286
rect 2682 1126 2685 1176
rect 2690 1133 2693 1216
rect 2682 1123 2693 1126
rect 2674 1103 2693 1106
rect 2610 883 2641 886
rect 2650 933 2661 936
rect 2598 823 2605 826
rect 2578 573 2581 823
rect 2586 673 2589 786
rect 2586 593 2589 626
rect 2594 623 2597 806
rect 2602 673 2605 823
rect 2610 813 2613 883
rect 2618 803 2621 816
rect 2610 616 2613 796
rect 2598 613 2613 616
rect 2570 543 2581 546
rect 2570 383 2573 536
rect 2578 533 2581 543
rect 2586 413 2589 586
rect 2598 556 2601 613
rect 2618 586 2621 726
rect 2610 583 2621 586
rect 2594 553 2601 556
rect 2594 496 2597 553
rect 2626 546 2629 826
rect 2634 723 2637 846
rect 2650 806 2653 933
rect 2658 813 2661 926
rect 2666 883 2669 1086
rect 2674 886 2677 1076
rect 2682 933 2685 1096
rect 2690 946 2693 1103
rect 2698 1003 2701 1596
rect 2706 1533 2709 1736
rect 2714 1716 2717 1726
rect 2730 1723 2733 1793
rect 2738 1736 2741 1846
rect 2746 1806 2749 1923
rect 2762 1913 2765 1926
rect 2770 1883 2773 1933
rect 2778 1826 2781 1926
rect 2754 1823 2781 1826
rect 2754 1813 2757 1823
rect 2746 1803 2757 1806
rect 2738 1733 2749 1736
rect 2738 1716 2741 1726
rect 2714 1713 2741 1716
rect 2714 1703 2717 1713
rect 2746 1706 2749 1733
rect 2730 1703 2749 1706
rect 2730 1626 2733 1703
rect 2754 1686 2757 1803
rect 2746 1683 2757 1686
rect 2746 1636 2749 1683
rect 2762 1653 2765 1806
rect 2770 1796 2773 1816
rect 2786 1813 2789 1926
rect 2794 1796 2797 1906
rect 2770 1793 2797 1796
rect 2746 1633 2757 1636
rect 2714 1533 2717 1626
rect 2722 1623 2733 1626
rect 2722 1556 2725 1623
rect 2754 1606 2757 1633
rect 2770 1613 2773 1786
rect 2746 1603 2757 1606
rect 2746 1596 2749 1603
rect 2738 1593 2749 1596
rect 2722 1553 2733 1556
rect 2722 1516 2725 1546
rect 2730 1523 2733 1553
rect 2738 1533 2741 1593
rect 2754 1553 2757 1596
rect 2762 1593 2765 1606
rect 2746 1536 2749 1546
rect 2746 1533 2765 1536
rect 2718 1513 2725 1516
rect 2706 1323 2709 1466
rect 2718 1446 2721 1513
rect 2718 1443 2725 1446
rect 2706 1203 2709 1226
rect 2714 1213 2717 1426
rect 2714 1133 2717 1176
rect 2706 973 2709 1126
rect 2722 1113 2725 1443
rect 2730 1203 2733 1486
rect 2738 1316 2741 1446
rect 2746 1436 2749 1533
rect 2762 1443 2765 1526
rect 2770 1473 2773 1526
rect 2746 1433 2757 1436
rect 2746 1403 2749 1426
rect 2746 1333 2749 1386
rect 2738 1313 2745 1316
rect 2742 1246 2745 1313
rect 2754 1253 2757 1433
rect 2770 1336 2773 1416
rect 2778 1413 2781 1746
rect 2786 1723 2789 1756
rect 2794 1713 2797 1736
rect 2802 1696 2805 2006
rect 2818 2003 2829 2006
rect 2818 1996 2821 2003
rect 2810 1993 2821 1996
rect 2810 1913 2813 1993
rect 2834 1986 2837 2136
rect 2842 2113 2845 2186
rect 2858 2183 2861 2206
rect 2842 2023 2845 2036
rect 2830 1983 2837 1986
rect 2830 1926 2833 1983
rect 2818 1883 2821 1926
rect 2826 1923 2833 1926
rect 2842 1923 2845 2006
rect 2850 1993 2853 2136
rect 2858 2096 2861 2126
rect 2866 2113 2869 2126
rect 2858 2093 2865 2096
rect 2862 1986 2865 2093
rect 2858 1983 2865 1986
rect 2826 1836 2829 1923
rect 2810 1833 2829 1836
rect 2810 1713 2813 1833
rect 2834 1826 2837 1916
rect 2850 1893 2853 1926
rect 2826 1823 2837 1826
rect 2802 1693 2809 1696
rect 2786 1393 2789 1636
rect 2762 1333 2773 1336
rect 2738 1243 2745 1246
rect 2738 1163 2741 1243
rect 2746 1213 2749 1226
rect 2746 1133 2749 1196
rect 2730 1113 2733 1126
rect 2690 943 2701 946
rect 2682 893 2685 916
rect 2674 883 2685 886
rect 2682 813 2685 883
rect 2642 803 2661 806
rect 2634 613 2637 666
rect 2642 603 2645 736
rect 2658 723 2661 796
rect 2666 783 2669 796
rect 2690 783 2693 936
rect 2698 863 2701 943
rect 2706 923 2709 966
rect 2714 803 2717 1036
rect 2722 873 2725 1086
rect 2730 813 2733 1066
rect 2738 913 2741 1036
rect 2746 1003 2749 1106
rect 2754 986 2757 1246
rect 2762 1176 2765 1333
rect 2770 1243 2773 1326
rect 2770 1183 2773 1216
rect 2762 1173 2773 1176
rect 2762 1036 2765 1166
rect 2770 1043 2773 1173
rect 2778 1133 2781 1346
rect 2794 1336 2797 1676
rect 2806 1616 2809 1693
rect 2818 1663 2821 1806
rect 2826 1743 2829 1823
rect 2834 1783 2837 1816
rect 2842 1793 2845 1806
rect 2802 1613 2809 1616
rect 2802 1596 2805 1613
rect 2826 1606 2829 1636
rect 2834 1613 2837 1736
rect 2842 1723 2845 1746
rect 2850 1716 2853 1816
rect 2858 1773 2861 1983
rect 2866 1913 2869 1936
rect 2874 1883 2877 2326
rect 2890 2203 2893 2316
rect 2898 2293 2901 2336
rect 2906 2226 2909 2366
rect 2962 2333 2965 2346
rect 2970 2316 2973 2326
rect 2978 2323 2981 2376
rect 2986 2316 2989 2526
rect 3058 2523 3085 2526
rect 2994 2333 2997 2416
rect 3042 2413 3045 2506
rect 3090 2413 3093 2526
rect 3098 2503 3101 2533
rect 3058 2393 3061 2406
rect 3018 2316 3021 2376
rect 3050 2343 3085 2346
rect 2970 2313 2989 2316
rect 3010 2313 3021 2316
rect 3010 2246 3013 2313
rect 3026 2246 3029 2336
rect 3050 2323 3053 2343
rect 3066 2326 3069 2336
rect 3058 2323 3069 2326
rect 3074 2323 3077 2336
rect 3058 2316 3061 2323
rect 3034 2313 3061 2316
rect 3066 2303 3069 2316
rect 3010 2243 3021 2246
rect 3026 2243 3053 2246
rect 2898 2223 2925 2226
rect 2898 2213 2901 2223
rect 2882 2133 2885 2196
rect 2882 2103 2885 2116
rect 2882 1923 2885 2026
rect 2866 1803 2869 1816
rect 2882 1803 2885 1916
rect 2890 1796 2893 2186
rect 2898 2103 2901 2206
rect 2906 2193 2909 2216
rect 2922 2196 2925 2206
rect 2930 2203 2933 2226
rect 2994 2216 2997 2226
rect 2978 2213 2997 2216
rect 2922 2193 2933 2196
rect 2906 2013 2909 2136
rect 2914 2123 2917 2166
rect 2922 2113 2925 2136
rect 2898 1933 2901 1996
rect 2898 1903 2901 1916
rect 2882 1793 2893 1796
rect 2850 1713 2861 1716
rect 2866 1706 2869 1756
rect 2874 1723 2877 1746
rect 2882 1733 2885 1793
rect 2862 1703 2869 1706
rect 2842 1623 2845 1646
rect 2826 1603 2845 1606
rect 2802 1593 2845 1596
rect 2802 1506 2805 1593
rect 2810 1526 2813 1536
rect 2834 1526 2837 1536
rect 2842 1533 2845 1556
rect 2810 1523 2837 1526
rect 2842 1513 2845 1526
rect 2850 1506 2853 1696
rect 2862 1546 2865 1703
rect 2874 1623 2877 1646
rect 2874 1573 2877 1616
rect 2882 1583 2885 1716
rect 2890 1566 2893 1736
rect 2886 1563 2893 1566
rect 2862 1543 2869 1546
rect 2802 1503 2813 1506
rect 2810 1446 2813 1503
rect 2826 1503 2853 1506
rect 2826 1456 2829 1503
rect 2802 1443 2813 1446
rect 2822 1453 2829 1456
rect 2802 1376 2805 1443
rect 2810 1403 2813 1426
rect 2822 1376 2825 1453
rect 2802 1373 2813 1376
rect 2822 1373 2829 1376
rect 2786 1333 2797 1336
rect 2786 1206 2789 1333
rect 2794 1223 2797 1326
rect 2802 1303 2805 1326
rect 2810 1313 2813 1336
rect 2818 1333 2821 1356
rect 2826 1283 2829 1373
rect 2786 1203 2793 1206
rect 2802 1203 2805 1246
rect 2790 1136 2793 1203
rect 2810 1196 2813 1256
rect 2818 1203 2821 1276
rect 2802 1193 2821 1196
rect 2818 1183 2821 1193
rect 2826 1166 2829 1216
rect 2834 1196 2837 1446
rect 2850 1413 2853 1426
rect 2858 1356 2861 1526
rect 2866 1403 2869 1543
rect 2874 1513 2877 1526
rect 2886 1476 2889 1563
rect 2886 1473 2893 1476
rect 2890 1453 2893 1473
rect 2874 1383 2877 1426
rect 2842 1353 2861 1356
rect 2842 1293 2845 1353
rect 2858 1336 2861 1346
rect 2850 1333 2861 1336
rect 2858 1306 2861 1326
rect 2854 1303 2861 1306
rect 2854 1236 2857 1303
rect 2842 1213 2845 1236
rect 2850 1233 2857 1236
rect 2850 1203 2853 1233
rect 2866 1203 2869 1376
rect 2874 1333 2877 1356
rect 2874 1213 2877 1326
rect 2882 1213 2885 1416
rect 2890 1403 2893 1416
rect 2890 1273 2893 1336
rect 2898 1326 2901 1816
rect 2906 1803 2909 2006
rect 2914 1933 2917 2066
rect 2922 2006 2925 2106
rect 2930 2063 2933 2193
rect 2938 2153 2941 2206
rect 2938 2133 2957 2136
rect 2946 2073 2949 2126
rect 2930 2013 2933 2056
rect 2946 2013 2949 2026
rect 2922 2003 2933 2006
rect 2938 2003 2949 2006
rect 2954 2003 2957 2133
rect 2962 2073 2965 2206
rect 2994 2193 2997 2206
rect 3002 2166 3005 2226
rect 2986 2163 3005 2166
rect 3010 2163 3013 2206
rect 2970 2136 2973 2156
rect 2970 2133 2977 2136
rect 2974 2046 2977 2133
rect 2986 2053 2989 2163
rect 3002 2143 3013 2146
rect 3002 2116 3005 2136
rect 3010 2133 3013 2143
rect 2998 2113 3005 2116
rect 3010 2113 3013 2126
rect 2970 2043 2977 2046
rect 2930 1916 2933 2003
rect 2946 1993 2949 2003
rect 2922 1913 2933 1916
rect 2922 1826 2925 1913
rect 2954 1866 2957 1926
rect 2962 1873 2965 2036
rect 2970 2023 2973 2043
rect 2998 2026 3001 2113
rect 3018 2106 3021 2243
rect 3026 2206 3029 2236
rect 3034 2213 3037 2226
rect 3026 2203 3037 2206
rect 3042 2196 3045 2226
rect 3026 2193 3045 2196
rect 3026 2136 3029 2193
rect 3026 2133 3037 2136
rect 3010 2103 3021 2106
rect 3026 2123 3037 2126
rect 2998 2023 3005 2026
rect 2970 1993 2973 2016
rect 2986 1936 2989 1956
rect 2994 1943 2997 2006
rect 2970 1933 2997 1936
rect 3002 1933 3005 2023
rect 3010 1996 3013 2103
rect 3026 2063 3029 2123
rect 3018 2003 3021 2056
rect 3034 2023 3037 2116
rect 3042 2003 3045 2136
rect 3010 1993 3029 1996
rect 2994 1923 2997 1933
rect 3010 1923 3021 1926
rect 2970 1913 2997 1916
rect 2970 1896 2973 1913
rect 2970 1893 2981 1896
rect 2954 1863 2965 1866
rect 2914 1823 2925 1826
rect 2906 1726 2909 1786
rect 2914 1733 2917 1823
rect 2922 1793 2925 1806
rect 2930 1733 2933 1806
rect 2946 1803 2949 1816
rect 2946 1766 2949 1786
rect 2942 1763 2949 1766
rect 2906 1723 2913 1726
rect 2910 1656 2913 1723
rect 2910 1653 2917 1656
rect 2906 1553 2909 1636
rect 2914 1623 2917 1653
rect 2922 1643 2925 1726
rect 2930 1673 2933 1716
rect 2942 1656 2945 1763
rect 2954 1753 2957 1816
rect 2962 1796 2965 1863
rect 2978 1836 2981 1893
rect 2970 1833 2981 1836
rect 2970 1813 2973 1833
rect 2970 1803 2981 1806
rect 2986 1796 2989 1816
rect 2962 1793 2989 1796
rect 2954 1713 2957 1736
rect 2970 1733 2973 1776
rect 2962 1706 2965 1726
rect 2978 1723 2981 1736
rect 2954 1703 2965 1706
rect 2954 1673 2957 1703
rect 2942 1653 2949 1656
rect 2946 1633 2949 1653
rect 2922 1563 2925 1616
rect 2930 1593 2933 1606
rect 2970 1603 2973 1716
rect 2986 1703 2989 1793
rect 2914 1513 2917 1536
rect 2922 1533 2933 1536
rect 2922 1496 2925 1526
rect 2946 1513 2949 1526
rect 2970 1523 2973 1586
rect 2970 1496 2973 1516
rect 2922 1493 2941 1496
rect 2906 1433 2917 1436
rect 2906 1413 2909 1426
rect 2914 1403 2917 1426
rect 2938 1396 2941 1493
rect 2962 1493 2973 1496
rect 2962 1446 2965 1493
rect 2978 1483 2981 1616
rect 2986 1513 2989 1646
rect 2994 1613 2997 1816
rect 3002 1603 3005 1806
rect 3010 1753 3013 1923
rect 3026 1916 3029 1993
rect 3034 1933 3037 1946
rect 3042 1933 3045 1956
rect 3022 1913 3029 1916
rect 3022 1826 3025 1913
rect 3018 1823 3025 1826
rect 3010 1586 3013 1736
rect 3018 1723 3021 1823
rect 3034 1813 3037 1916
rect 3042 1813 3045 1886
rect 3018 1613 3021 1636
rect 3010 1583 3021 1586
rect 2962 1443 2973 1446
rect 2994 1443 2997 1546
rect 2970 1426 2973 1443
rect 2978 1433 2997 1436
rect 2970 1423 2989 1426
rect 2994 1413 2997 1433
rect 3002 1406 3005 1566
rect 2986 1403 3005 1406
rect 2906 1343 2909 1396
rect 2922 1393 2941 1396
rect 2898 1323 2909 1326
rect 2906 1266 2909 1323
rect 2898 1263 2909 1266
rect 2834 1193 2853 1196
rect 2874 1193 2877 1206
rect 2818 1163 2829 1166
rect 2790 1133 2797 1136
rect 2786 1103 2789 1126
rect 2794 1083 2797 1133
rect 2818 1066 2821 1163
rect 2834 1123 2837 1186
rect 2842 1123 2845 1146
rect 2818 1063 2825 1066
rect 2778 1043 2805 1046
rect 2762 1033 2773 1036
rect 2778 1033 2781 1043
rect 2770 1026 2773 1033
rect 2746 983 2757 986
rect 2746 953 2749 983
rect 2762 976 2765 1026
rect 2770 1023 2789 1026
rect 2794 1016 2797 1036
rect 2770 1013 2797 1016
rect 2802 1006 2805 1043
rect 2822 1006 2825 1063
rect 2834 1026 2837 1096
rect 2850 1073 2853 1193
rect 2858 1133 2861 1176
rect 2890 1126 2893 1176
rect 2898 1143 2901 1263
rect 2890 1123 2897 1126
rect 2842 1043 2869 1046
rect 2842 1033 2845 1043
rect 2834 1023 2853 1026
rect 2858 1016 2861 1036
rect 2834 1013 2861 1016
rect 2802 1003 2813 1006
rect 2822 1003 2829 1006
rect 2754 973 2765 976
rect 2754 923 2757 973
rect 2770 913 2773 956
rect 2810 923 2813 1003
rect 2826 916 2829 1003
rect 2866 936 2869 1043
rect 2842 933 2869 936
rect 2874 933 2877 1036
rect 2882 943 2885 1116
rect 2894 1046 2897 1123
rect 2894 1043 2901 1046
rect 2890 936 2893 1026
rect 2882 933 2893 936
rect 2762 903 2781 906
rect 2810 866 2813 916
rect 2818 913 2829 916
rect 2818 876 2821 906
rect 2834 876 2837 926
rect 2818 873 2837 876
rect 2842 866 2845 933
rect 2882 926 2885 933
rect 2858 923 2885 926
rect 2882 903 2885 923
rect 2810 863 2845 866
rect 2714 766 2717 786
rect 2714 763 2721 766
rect 2690 733 2693 746
rect 2718 696 2721 763
rect 2730 743 2733 806
rect 2738 723 2741 736
rect 2770 723 2773 806
rect 2778 733 2781 816
rect 2802 813 2813 816
rect 2842 803 2845 846
rect 2890 813 2893 866
rect 2898 853 2901 1043
rect 2906 1023 2909 1236
rect 2922 1226 2925 1393
rect 2930 1333 2949 1336
rect 2938 1296 2941 1326
rect 2938 1293 2949 1296
rect 2922 1223 2933 1226
rect 2914 1203 2917 1216
rect 2914 1066 2917 1156
rect 2922 1123 2925 1216
rect 2930 1076 2933 1223
rect 2938 1143 2941 1286
rect 2946 1203 2949 1293
rect 2954 1283 2957 1356
rect 2946 1123 2949 1186
rect 2954 1176 2957 1266
rect 2962 1203 2965 1346
rect 2970 1333 2973 1396
rect 2986 1386 2989 1403
rect 2982 1383 2989 1386
rect 2982 1326 2985 1383
rect 2994 1353 2997 1396
rect 2994 1333 2997 1346
rect 3002 1333 3005 1366
rect 2970 1293 2973 1326
rect 2982 1323 2989 1326
rect 3010 1323 3013 1576
rect 3018 1373 3021 1583
rect 3026 1343 3029 1806
rect 3050 1803 3053 2243
rect 3058 2193 3061 2246
rect 3074 2186 3077 2236
rect 3082 2206 3085 2343
rect 3090 2333 3093 2346
rect 3106 2233 3109 2676
rect 3130 2646 3133 2703
rect 3130 2643 3141 2646
rect 3114 2513 3117 2596
rect 3098 2223 3117 2226
rect 3090 2213 3101 2216
rect 3082 2203 3101 2206
rect 3074 2183 3085 2186
rect 3058 2113 3061 2136
rect 3066 2123 3069 2166
rect 3074 2103 3077 2136
rect 3082 2096 3085 2183
rect 3074 2093 3085 2096
rect 3034 1713 3037 1756
rect 3042 1643 3045 1726
rect 3050 1653 3053 1736
rect 3034 1543 3037 1606
rect 3058 1603 3061 2026
rect 3066 1823 3069 2016
rect 3074 1976 3077 2093
rect 3090 2016 3093 2196
rect 3098 2073 3101 2156
rect 3114 2133 3117 2223
rect 3114 2113 3117 2126
rect 3122 2096 3125 2486
rect 3130 2423 3133 2626
rect 3138 2603 3141 2643
rect 3146 2633 3149 2796
rect 3154 2716 3157 2803
rect 3162 2803 3173 2806
rect 3162 2726 3165 2803
rect 3178 2793 3181 2826
rect 3210 2823 3213 2843
rect 3194 2783 3197 2816
rect 3218 2803 3221 3026
rect 3226 3003 3229 3123
rect 3234 3096 3237 3116
rect 3234 3093 3245 3096
rect 3242 3046 3245 3093
rect 3234 3043 3245 3046
rect 3234 2956 3237 3043
rect 3258 3013 3261 3026
rect 3250 2993 3253 3006
rect 3230 2953 3237 2956
rect 3230 2906 3233 2953
rect 3266 2943 3269 3126
rect 3230 2903 3237 2906
rect 3234 2746 3237 2903
rect 3250 2876 3253 2936
rect 3274 2923 3277 3016
rect 3282 3003 3285 3116
rect 3298 3076 3301 3216
rect 3306 3213 3309 3253
rect 3330 3106 3333 3126
rect 3338 3113 3341 3216
rect 3346 3213 3349 3253
rect 3370 3223 3413 3226
rect 3370 3203 3373 3223
rect 3378 3213 3389 3216
rect 3378 3203 3389 3206
rect 3410 3203 3413 3223
rect 3346 3143 3381 3146
rect 3330 3103 3337 3106
rect 3298 3073 3325 3076
rect 3290 3013 3293 3026
rect 3314 2973 3317 3016
rect 3322 2986 3325 3073
rect 3334 3046 3337 3103
rect 3346 3053 3349 3143
rect 3334 3043 3341 3046
rect 3322 2983 3333 2986
rect 3250 2873 3261 2876
rect 3314 2873 3317 2956
rect 3258 2776 3261 2873
rect 3250 2773 3261 2776
rect 3250 2753 3253 2773
rect 3282 2746 3285 2826
rect 3306 2796 3309 2816
rect 3314 2803 3317 2826
rect 3322 2796 3325 2946
rect 3330 2886 3333 2983
rect 3338 2953 3341 3043
rect 3362 3013 3365 3136
rect 3370 3096 3373 3143
rect 3378 3133 3381 3143
rect 3386 3126 3389 3203
rect 3418 3133 3421 3226
rect 3378 3116 3381 3126
rect 3386 3123 3413 3126
rect 3378 3113 3405 3116
rect 3370 3093 3381 3096
rect 3378 3006 3381 3093
rect 3370 3003 3381 3006
rect 3346 2923 3349 2936
rect 3370 2916 3373 3003
rect 3378 2923 3381 2976
rect 3410 2926 3413 3123
rect 3418 2993 3421 3016
rect 3410 2923 3429 2926
rect 3370 2913 3389 2916
rect 3330 2883 3373 2886
rect 3338 2803 3341 2876
rect 3362 2813 3365 2826
rect 3302 2793 3309 2796
rect 3314 2793 3325 2796
rect 3234 2743 3241 2746
rect 3282 2743 3293 2746
rect 3178 2733 3189 2736
rect 3162 2723 3189 2726
rect 3154 2713 3189 2716
rect 3194 2686 3197 2736
rect 3194 2683 3221 2686
rect 3154 2523 3157 2616
rect 3218 2606 3221 2683
rect 3226 2613 3229 2736
rect 3238 2666 3241 2743
rect 3274 2726 3277 2736
rect 3234 2663 3241 2666
rect 3234 2643 3237 2663
rect 3234 2606 3237 2616
rect 3250 2613 3253 2726
rect 3266 2723 3277 2726
rect 3266 2626 3269 2723
rect 3282 2716 3285 2726
rect 3290 2723 3293 2743
rect 3302 2716 3305 2793
rect 3274 2683 3277 2716
rect 3282 2713 3305 2716
rect 3282 2636 3285 2666
rect 3282 2633 3293 2636
rect 3162 2513 3165 2606
rect 3170 2603 3181 2606
rect 3218 2603 3237 2606
rect 3170 2466 3173 2603
rect 3194 2533 3197 2546
rect 3170 2463 3197 2466
rect 3138 2453 3181 2456
rect 3138 2413 3141 2453
rect 3178 2413 3181 2453
rect 3194 2406 3197 2463
rect 3154 2393 3157 2406
rect 3186 2403 3197 2406
rect 3186 2346 3189 2403
rect 3130 2343 3189 2346
rect 3130 2203 3133 2226
rect 3138 2153 3141 2336
rect 3154 2323 3157 2336
rect 3170 2333 3173 2343
rect 3162 2306 3165 2326
rect 3162 2303 3173 2306
rect 3138 2133 3141 2146
rect 3146 2143 3149 2186
rect 3154 2133 3157 2276
rect 3170 2226 3173 2303
rect 3162 2223 3173 2226
rect 3162 2166 3165 2223
rect 3178 2173 3181 2196
rect 3162 2163 3189 2166
rect 3162 2133 3165 2146
rect 3170 2143 3181 2146
rect 3118 2093 3125 2096
rect 3130 2123 3165 2126
rect 3118 2026 3121 2093
rect 3118 2023 3125 2026
rect 3090 2013 3101 2016
rect 3082 2003 3093 2006
rect 3090 1993 3093 2003
rect 3074 1973 3085 1976
rect 3082 1836 3085 1973
rect 3098 1926 3101 2013
rect 3106 1993 3109 2016
rect 3106 1973 3109 1986
rect 3114 1933 3117 2006
rect 3074 1833 3085 1836
rect 3094 1923 3101 1926
rect 3066 1793 3069 1806
rect 3066 1733 3069 1786
rect 3066 1603 3069 1656
rect 3074 1596 3077 1833
rect 3082 1803 3085 1816
rect 3094 1806 3097 1923
rect 3106 1816 3109 1916
rect 3106 1813 3113 1816
rect 3094 1803 3101 1806
rect 3098 1783 3101 1803
rect 3090 1733 3093 1776
rect 3110 1766 3113 1813
rect 3082 1723 3093 1726
rect 3098 1723 3101 1766
rect 3106 1763 3113 1766
rect 3090 1663 3093 1723
rect 3106 1676 3109 1763
rect 3114 1723 3117 1746
rect 3122 1683 3125 2023
rect 3130 1933 3133 2123
rect 3138 1943 3141 1986
rect 3138 1813 3141 1826
rect 3130 1793 3133 1806
rect 3146 1786 3149 2116
rect 3154 1933 3157 1986
rect 3154 1813 3157 1836
rect 3130 1783 3149 1786
rect 3098 1673 3109 1676
rect 3042 1593 3077 1596
rect 3042 1536 3045 1593
rect 3034 1533 3045 1536
rect 3034 1336 3037 1533
rect 3050 1523 3053 1556
rect 3066 1523 3069 1586
rect 3082 1576 3085 1616
rect 3078 1573 3085 1576
rect 3078 1516 3081 1573
rect 3050 1506 3053 1516
rect 3050 1503 3061 1506
rect 3042 1466 3045 1486
rect 3042 1463 3049 1466
rect 3046 1336 3049 1463
rect 3066 1443 3069 1516
rect 3078 1513 3085 1516
rect 3090 1513 3093 1646
rect 3098 1613 3101 1673
rect 3098 1586 3101 1606
rect 3106 1603 3109 1626
rect 3098 1583 3105 1586
rect 3026 1333 3037 1336
rect 3042 1333 3049 1336
rect 3058 1333 3061 1436
rect 3066 1393 3069 1426
rect 3066 1333 3069 1366
rect 2986 1306 2989 1323
rect 2986 1303 2997 1306
rect 2970 1273 2981 1276
rect 2970 1183 2973 1216
rect 2978 1203 2981 1273
rect 2954 1173 2977 1176
rect 2974 1126 2977 1173
rect 2994 1156 2997 1303
rect 3018 1213 3021 1236
rect 3026 1216 3029 1333
rect 3034 1223 3037 1246
rect 3026 1213 3037 1216
rect 2986 1153 2997 1156
rect 2986 1133 2989 1153
rect 3018 1136 3021 1166
rect 3010 1133 3021 1136
rect 2974 1123 2981 1126
rect 2930 1073 2937 1076
rect 2914 1063 2925 1066
rect 2914 1023 2917 1036
rect 2922 973 2925 1063
rect 2934 966 2937 1073
rect 2930 963 2937 966
rect 2906 913 2909 936
rect 2914 906 2917 926
rect 2914 903 2925 906
rect 2906 823 2909 876
rect 2922 823 2925 846
rect 2890 776 2893 806
rect 2906 803 2909 816
rect 2882 773 2893 776
rect 2842 733 2845 746
rect 2842 716 2845 726
rect 2858 723 2861 746
rect 2866 716 2869 726
rect 2842 713 2869 716
rect 2714 693 2721 696
rect 2602 523 2605 536
rect 2610 523 2613 546
rect 2618 543 2629 546
rect 2594 493 2605 496
rect 2602 436 2605 493
rect 2594 433 2605 436
rect 2570 323 2573 336
rect 2570 313 2589 316
rect 2570 306 2573 313
rect 2594 306 2597 433
rect 2602 403 2605 416
rect 2618 413 2621 543
rect 2634 513 2645 516
rect 2634 413 2637 513
rect 2650 483 2653 636
rect 2658 586 2661 606
rect 2666 603 2669 676
rect 2658 583 2665 586
rect 2662 476 2665 583
rect 2658 473 2665 476
rect 2658 416 2661 473
rect 2674 453 2677 606
rect 2698 603 2701 616
rect 2714 613 2717 693
rect 2722 603 2725 676
rect 2882 646 2885 773
rect 2882 643 2893 646
rect 2842 623 2877 626
rect 2722 586 2725 596
rect 2698 583 2725 586
rect 2682 523 2693 526
rect 2658 413 2665 416
rect 2602 313 2605 336
rect 2618 323 2621 406
rect 2642 403 2653 406
rect 2650 313 2653 403
rect 2662 366 2665 413
rect 2674 406 2677 436
rect 2682 423 2685 523
rect 2698 516 2701 583
rect 2746 576 2749 596
rect 2690 513 2701 516
rect 2706 513 2709 576
rect 2722 573 2749 576
rect 2722 543 2725 573
rect 2754 556 2757 616
rect 2778 613 2797 616
rect 2842 613 2845 623
rect 2858 613 2869 616
rect 2874 613 2877 623
rect 2762 586 2765 606
rect 2762 583 2769 586
rect 2738 553 2757 556
rect 2714 523 2717 536
rect 2738 506 2741 553
rect 2698 503 2741 506
rect 2746 503 2749 536
rect 2766 506 2769 583
rect 2778 543 2781 613
rect 2794 596 2797 613
rect 2794 593 2805 596
rect 2834 593 2837 606
rect 2778 533 2797 536
rect 2778 523 2781 533
rect 2794 513 2797 526
rect 2802 523 2805 593
rect 2818 523 2821 576
rect 2766 503 2773 506
rect 2738 466 2741 503
rect 2738 463 2757 466
rect 2706 406 2709 426
rect 2674 403 2685 406
rect 2658 363 2665 366
rect 2658 343 2661 363
rect 2682 356 2685 403
rect 2674 353 2685 356
rect 2698 403 2709 406
rect 2658 313 2661 336
rect 2674 316 2677 353
rect 2698 346 2701 403
rect 2698 343 2709 346
rect 2674 313 2685 316
rect 2538 303 2573 306
rect 2554 266 2557 296
rect 2578 286 2581 306
rect 2574 283 2581 286
rect 2586 303 2597 306
rect 2554 263 2565 266
rect 2522 213 2533 216
rect 2522 153 2525 213
rect 2530 193 2533 206
rect 2546 203 2549 216
rect 2562 186 2565 263
rect 2574 196 2577 283
rect 2586 213 2589 303
rect 2602 246 2605 306
rect 2634 303 2645 306
rect 2634 246 2637 303
rect 2602 243 2621 246
rect 2634 243 2641 246
rect 2602 213 2605 243
rect 2618 236 2621 243
rect 2610 206 2613 236
rect 2618 233 2629 236
rect 2618 213 2621 226
rect 2626 206 2629 226
rect 2602 203 2629 206
rect 2574 193 2581 196
rect 2554 183 2565 186
rect 2482 123 2493 126
rect 2498 83 2501 136
rect 2506 123 2509 136
rect 2554 126 2557 183
rect 2554 123 2565 126
rect 2562 103 2565 123
rect 2578 113 2581 193
rect 2602 186 2605 203
rect 2594 183 2605 186
rect 2594 126 2597 183
rect 2594 123 2605 126
rect 2594 96 2597 106
rect 2602 103 2605 123
rect 2610 113 2613 196
rect 2638 176 2641 243
rect 2674 236 2677 313
rect 2698 306 2701 326
rect 2634 173 2641 176
rect 2650 233 2677 236
rect 2694 303 2701 306
rect 2694 236 2697 303
rect 2694 233 2701 236
rect 2634 156 2637 173
rect 2626 153 2637 156
rect 2626 126 2629 153
rect 2650 133 2653 233
rect 2674 223 2685 226
rect 2698 216 2701 233
rect 2666 213 2701 216
rect 2706 206 2709 343
rect 2714 333 2717 416
rect 2730 413 2733 426
rect 2738 413 2741 456
rect 2714 313 2717 326
rect 2738 323 2741 406
rect 2754 376 2757 463
rect 2750 373 2757 376
rect 2750 316 2753 373
rect 2770 356 2773 503
rect 2826 446 2829 536
rect 2826 443 2837 446
rect 2810 393 2813 406
rect 2834 356 2837 443
rect 2850 413 2853 606
rect 2866 553 2869 606
rect 2890 603 2893 643
rect 2874 533 2893 536
rect 2882 513 2885 526
rect 2690 203 2709 206
rect 2722 203 2725 316
rect 2746 313 2753 316
rect 2762 353 2773 356
rect 2730 293 2733 306
rect 2746 236 2749 313
rect 2762 243 2765 353
rect 2770 303 2773 316
rect 2778 313 2781 326
rect 2786 303 2789 336
rect 2794 323 2797 356
rect 2826 353 2837 356
rect 2826 306 2829 353
rect 2858 333 2861 346
rect 2826 303 2837 306
rect 2738 216 2741 236
rect 2746 233 2773 236
rect 2734 213 2741 216
rect 2690 173 2693 203
rect 2734 146 2737 213
rect 2734 143 2741 146
rect 2618 123 2629 126
rect 2618 96 2621 123
rect 2722 113 2725 136
rect 2738 123 2741 143
rect 2746 113 2749 206
rect 2754 196 2757 216
rect 2770 203 2773 233
rect 2778 223 2781 236
rect 2778 196 2781 216
rect 2754 193 2781 196
rect 2786 156 2789 266
rect 2826 203 2829 256
rect 2834 233 2837 303
rect 2890 253 2893 533
rect 2898 506 2901 786
rect 2914 733 2917 766
rect 2922 626 2925 726
rect 2930 683 2933 963
rect 2938 923 2941 936
rect 2946 933 2949 1036
rect 2954 983 2957 1116
rect 2962 996 2965 1026
rect 2978 1023 2981 1123
rect 3010 1056 3013 1133
rect 3010 1053 3021 1056
rect 3010 1016 3013 1036
rect 2978 1013 2989 1016
rect 3002 1013 3013 1016
rect 2962 993 2973 996
rect 2986 993 2989 1006
rect 2954 913 2957 976
rect 2970 916 2973 993
rect 3002 956 3005 1013
rect 3018 966 3021 1053
rect 3034 1003 3037 1213
rect 3042 1203 3045 1333
rect 3050 1313 3061 1316
rect 3066 1296 3069 1326
rect 3050 1213 3053 1296
rect 3062 1293 3069 1296
rect 3062 1226 3065 1293
rect 3062 1223 3069 1226
rect 3066 1203 3069 1223
rect 3058 996 3061 1186
rect 3074 1173 3077 1496
rect 3082 1433 3085 1513
rect 3102 1506 3105 1583
rect 3114 1553 3117 1616
rect 3122 1606 3125 1636
rect 3130 1613 3133 1783
rect 3154 1746 3157 1806
rect 3162 1756 3165 2076
rect 3170 2003 3173 2136
rect 3178 2123 3181 2143
rect 3178 1986 3181 2046
rect 3186 1993 3189 2163
rect 3194 2083 3197 2126
rect 3202 2023 3205 2206
rect 3210 2096 3213 2326
rect 3218 2313 3221 2603
rect 3242 2593 3245 2606
rect 3258 2603 3261 2626
rect 3266 2623 3277 2626
rect 3266 2603 3269 2616
rect 3226 2333 3229 2586
rect 3274 2583 3277 2623
rect 3290 2576 3293 2633
rect 3282 2573 3293 2576
rect 3282 2556 3285 2573
rect 3278 2553 3285 2556
rect 3266 2526 3269 2536
rect 3258 2523 3269 2526
rect 3258 2516 3261 2523
rect 3234 2513 3261 2516
rect 3266 2506 3269 2516
rect 3242 2503 3269 2506
rect 3242 2446 3245 2503
rect 3278 2496 3281 2553
rect 3306 2533 3309 2616
rect 3314 2586 3317 2793
rect 3338 2663 3341 2756
rect 3362 2696 3365 2796
rect 3354 2693 3365 2696
rect 3330 2616 3333 2626
rect 3322 2613 3333 2616
rect 3338 2593 3341 2616
rect 3354 2603 3357 2693
rect 3370 2606 3373 2883
rect 3386 2866 3389 2913
rect 3382 2863 3389 2866
rect 3382 2786 3385 2863
rect 3426 2826 3429 2923
rect 3426 2823 3433 2826
rect 3378 2783 3385 2786
rect 3378 2716 3381 2783
rect 3418 2766 3421 2816
rect 3386 2763 3421 2766
rect 3386 2723 3389 2763
rect 3378 2713 3389 2716
rect 3418 2713 3421 2726
rect 3370 2603 3377 2606
rect 3314 2583 3341 2586
rect 3234 2443 3245 2446
rect 3266 2493 3281 2496
rect 3234 2333 3237 2443
rect 3250 2413 3253 2426
rect 3266 2393 3269 2493
rect 3290 2396 3293 2526
rect 3314 2506 3317 2583
rect 3338 2533 3341 2583
rect 3362 2523 3365 2596
rect 3374 2516 3377 2603
rect 3306 2503 3317 2506
rect 3370 2513 3377 2516
rect 3306 2486 3309 2503
rect 3302 2483 3309 2486
rect 3302 2406 3305 2483
rect 3314 2413 3317 2496
rect 3346 2426 3349 2436
rect 3370 2433 3373 2513
rect 3330 2423 3357 2426
rect 3362 2423 3373 2426
rect 3302 2403 3309 2406
rect 3282 2393 3293 2396
rect 3258 2333 3261 2346
rect 3218 2213 3221 2256
rect 3242 2213 3253 2216
rect 3274 2206 3277 2356
rect 3282 2323 3285 2393
rect 3306 2306 3309 2403
rect 3330 2336 3333 2423
rect 3378 2416 3381 2426
rect 3346 2403 3349 2416
rect 3362 2413 3381 2416
rect 3314 2333 3333 2336
rect 3298 2303 3309 2306
rect 3298 2226 3301 2303
rect 3298 2223 3317 2226
rect 3226 2153 3229 2196
rect 3234 2146 3237 2206
rect 3266 2203 3277 2206
rect 3226 2143 3237 2146
rect 3226 2116 3229 2143
rect 3234 2126 3237 2136
rect 3250 2133 3253 2186
rect 3266 2156 3269 2203
rect 3282 2183 3285 2196
rect 3290 2166 3293 2206
rect 3306 2203 3309 2216
rect 3314 2186 3317 2223
rect 3322 2213 3325 2326
rect 3338 2266 3341 2336
rect 3346 2333 3349 2356
rect 3362 2346 3365 2413
rect 3386 2396 3389 2713
rect 3430 2706 3433 2823
rect 3426 2703 3433 2706
rect 3402 2613 3405 2626
rect 3426 2596 3429 2703
rect 3418 2593 3429 2596
rect 3418 2536 3421 2593
rect 3406 2533 3421 2536
rect 3406 2486 3409 2533
rect 3418 2493 3421 2526
rect 3402 2483 3409 2486
rect 3394 2423 3397 2436
rect 3402 2433 3405 2483
rect 3402 2416 3405 2426
rect 3394 2413 3405 2416
rect 3354 2343 3365 2346
rect 3378 2393 3389 2396
rect 3354 2313 3357 2343
rect 3362 2303 3365 2326
rect 3378 2316 3381 2393
rect 3426 2376 3429 2426
rect 3394 2373 3429 2376
rect 3394 2323 3397 2373
rect 3378 2313 3389 2316
rect 3330 2263 3341 2266
rect 3330 2203 3333 2263
rect 3386 2256 3389 2313
rect 3402 2303 3405 2326
rect 3418 2286 3421 2316
rect 3410 2283 3421 2286
rect 3386 2253 3397 2256
rect 3346 2243 3373 2246
rect 3346 2193 3349 2243
rect 3362 2213 3365 2236
rect 3314 2183 3349 2186
rect 3290 2163 3317 2166
rect 3266 2153 3277 2156
rect 3266 2126 3269 2136
rect 3234 2123 3269 2126
rect 3226 2113 3245 2116
rect 3210 2093 3221 2096
rect 3218 2036 3221 2093
rect 3242 2056 3245 2113
rect 3242 2053 3253 2056
rect 3210 2033 3221 2036
rect 3210 2016 3213 2033
rect 3202 2013 3213 2016
rect 3178 1983 3189 1986
rect 3170 1803 3173 1916
rect 3178 1766 3181 1946
rect 3186 1823 3189 1983
rect 3202 1956 3205 2013
rect 3210 1993 3213 2006
rect 3226 1956 3229 2016
rect 3234 2013 3237 2036
rect 3250 2013 3253 2053
rect 3202 1953 3213 1956
rect 3194 1906 3197 1926
rect 3202 1923 3205 1946
rect 3194 1903 3201 1906
rect 3198 1836 3201 1903
rect 3194 1833 3201 1836
rect 3194 1793 3197 1833
rect 3178 1763 3197 1766
rect 3162 1753 3181 1756
rect 3154 1743 3165 1746
rect 3138 1716 3141 1736
rect 3162 1733 3165 1743
rect 3138 1713 3145 1716
rect 3142 1626 3145 1713
rect 3154 1713 3165 1716
rect 3154 1663 3157 1713
rect 3170 1703 3173 1726
rect 3178 1696 3181 1753
rect 3186 1733 3189 1746
rect 3194 1733 3197 1763
rect 3162 1693 3181 1696
rect 3162 1636 3165 1693
rect 3138 1623 3145 1626
rect 3158 1633 3165 1636
rect 3122 1603 3133 1606
rect 3098 1503 3105 1506
rect 3090 1423 3093 1436
rect 3082 1323 3085 1416
rect 3098 1406 3101 1503
rect 3106 1433 3109 1446
rect 3094 1403 3101 1406
rect 3106 1403 3109 1426
rect 3094 1256 3097 1403
rect 3106 1343 3109 1396
rect 3094 1253 3101 1256
rect 3090 1223 3093 1236
rect 3090 1193 3093 1216
rect 3074 1026 3077 1146
rect 3098 1056 3101 1253
rect 3106 1203 3109 1326
rect 3114 1296 3117 1416
rect 3114 1293 3121 1296
rect 3118 1196 3121 1293
rect 3114 1193 3121 1196
rect 3114 1116 3117 1193
rect 3130 1183 3133 1603
rect 3138 1563 3141 1623
rect 3146 1546 3149 1606
rect 3158 1586 3161 1633
rect 3158 1583 3165 1586
rect 3146 1543 3157 1546
rect 3154 1413 3157 1543
rect 3162 1396 3165 1583
rect 3178 1573 3181 1686
rect 3178 1513 3181 1526
rect 3158 1393 3165 1396
rect 3158 1226 3161 1393
rect 3158 1223 3165 1226
rect 3138 1203 3141 1216
rect 3130 1143 3133 1156
rect 3154 1136 3157 1206
rect 3138 1133 3157 1136
rect 3162 1126 3165 1223
rect 3146 1123 3165 1126
rect 3114 1113 3125 1116
rect 3098 1053 3105 1056
rect 3050 993 3061 996
rect 3070 1023 3077 1026
rect 3018 963 3029 966
rect 2986 933 2989 956
rect 3002 953 3013 956
rect 2986 916 2989 926
rect 3002 923 3005 936
rect 3010 923 3013 953
rect 3026 916 3029 963
rect 2970 913 2989 916
rect 3018 913 3029 916
rect 2938 723 2941 866
rect 2946 856 2949 876
rect 2946 853 2957 856
rect 2954 786 2957 853
rect 3018 846 3021 913
rect 3018 843 3029 846
rect 2946 783 2957 786
rect 2946 696 2949 783
rect 2986 776 2989 826
rect 3002 783 3005 806
rect 3026 776 3029 843
rect 3050 826 3053 993
rect 3070 976 3073 1023
rect 3082 983 3085 1016
rect 3102 986 3105 1053
rect 3122 1046 3125 1113
rect 3098 983 3105 986
rect 3114 1043 3125 1046
rect 3070 973 3077 976
rect 3074 946 3077 973
rect 3098 963 3101 983
rect 3074 943 3081 946
rect 3078 896 3081 943
rect 3042 823 3053 826
rect 3074 893 3081 896
rect 3042 783 3045 823
rect 3050 793 3053 816
rect 2986 773 3005 776
rect 2954 733 2957 766
rect 2962 736 2965 746
rect 2962 733 2997 736
rect 2970 703 2973 726
rect 2946 693 2973 696
rect 2922 623 2965 626
rect 2938 613 2965 616
rect 2906 523 2909 606
rect 2938 603 2941 613
rect 2962 586 2965 606
rect 2954 583 2965 586
rect 2898 503 2909 506
rect 2906 386 2909 503
rect 2930 473 2933 536
rect 2938 513 2941 526
rect 2954 516 2957 583
rect 2970 523 2973 693
rect 2978 583 2981 733
rect 2986 706 2989 726
rect 3002 723 3005 773
rect 3010 773 3029 776
rect 2986 703 2997 706
rect 2994 646 2997 703
rect 2986 643 2997 646
rect 2986 626 2989 643
rect 3010 633 3013 773
rect 3018 646 3021 736
rect 3066 733 3069 746
rect 3050 703 3053 726
rect 3018 643 3053 646
rect 2986 623 3045 626
rect 2986 533 2989 596
rect 3002 586 3005 616
rect 3026 613 3045 616
rect 2994 583 3005 586
rect 2994 523 2997 583
rect 2954 513 2965 516
rect 2930 393 2933 406
rect 2898 383 2909 386
rect 2898 343 2901 383
rect 2962 366 2965 513
rect 3002 486 3005 536
rect 3018 533 3021 576
rect 3010 513 3013 526
rect 2978 483 3005 486
rect 2978 413 2981 483
rect 2906 363 2965 366
rect 2906 323 2909 363
rect 3010 346 3013 476
rect 3026 403 3029 596
rect 3042 586 3045 606
rect 3050 603 3053 643
rect 3038 583 3045 586
rect 3038 416 3041 583
rect 3034 413 3041 416
rect 3050 413 3053 596
rect 3058 423 3061 536
rect 3066 523 3069 536
rect 3066 413 3069 516
rect 3074 506 3077 893
rect 3090 813 3093 956
rect 3090 776 3093 806
rect 3098 783 3101 936
rect 3086 773 3093 776
rect 3086 726 3089 773
rect 3106 763 3109 816
rect 3114 753 3117 1043
rect 3122 896 3125 996
rect 3130 943 3133 1016
rect 3138 1013 3141 1026
rect 3138 913 3141 926
rect 3146 923 3149 1123
rect 3170 1023 3173 1506
rect 3178 1323 3181 1406
rect 3178 1223 3181 1236
rect 3186 1233 3189 1246
rect 3186 1213 3189 1226
rect 3178 1133 3181 1206
rect 3178 1113 3181 1126
rect 3186 1123 3189 1176
rect 3194 1163 3197 1536
rect 3202 1476 3205 1746
rect 3210 1583 3213 1953
rect 3218 1953 3229 1956
rect 3218 1916 3221 1953
rect 3234 1946 3237 2006
rect 3226 1943 3237 1946
rect 3226 1933 3229 1943
rect 3218 1913 3229 1916
rect 3226 1846 3229 1913
rect 3218 1843 3229 1846
rect 3210 1493 3213 1526
rect 3218 1503 3221 1843
rect 3226 1653 3229 1826
rect 3242 1793 3245 1946
rect 3258 1913 3261 2096
rect 3266 1896 3269 2123
rect 3258 1893 3269 1896
rect 3258 1766 3261 1893
rect 3258 1763 3269 1766
rect 3266 1743 3269 1763
rect 3274 1736 3277 2153
rect 3282 2136 3285 2146
rect 3306 2143 3309 2156
rect 3282 2133 3301 2136
rect 3314 2126 3317 2163
rect 3282 2043 3285 2126
rect 3298 2123 3317 2126
rect 3322 2116 3325 2176
rect 3330 2123 3333 2146
rect 3338 2123 3341 2136
rect 3346 2116 3349 2183
rect 3354 2136 3357 2206
rect 3362 2163 3365 2206
rect 3370 2173 3373 2243
rect 3394 2186 3397 2253
rect 3410 2206 3413 2283
rect 3426 2213 3429 2326
rect 3410 2203 3421 2206
rect 3386 2183 3397 2186
rect 3370 2143 3373 2156
rect 3354 2133 3373 2136
rect 3282 1923 3285 2006
rect 3290 1913 3293 1946
rect 3298 1896 3301 2026
rect 3306 2003 3309 2116
rect 3322 2113 3333 2116
rect 3346 2113 3365 2116
rect 3306 1923 3309 1936
rect 3314 1933 3317 1986
rect 3330 1956 3333 2113
rect 3362 2026 3365 2113
rect 3326 1953 3333 1956
rect 3346 2023 3365 2026
rect 3294 1893 3301 1896
rect 3306 1896 3309 1916
rect 3326 1906 3329 1953
rect 3326 1903 3333 1906
rect 3306 1893 3317 1896
rect 3294 1836 3297 1893
rect 3314 1846 3317 1893
rect 3306 1843 3317 1846
rect 3294 1833 3301 1836
rect 3298 1816 3301 1833
rect 3282 1803 3285 1816
rect 3290 1813 3301 1816
rect 3306 1813 3309 1843
rect 3330 1826 3333 1903
rect 3346 1876 3349 2023
rect 3354 1993 3357 2006
rect 3386 1993 3389 2183
rect 3418 2166 3421 2203
rect 3402 2133 3405 2166
rect 3418 2163 3429 2166
rect 3394 2103 3397 2126
rect 3410 2123 3413 2156
rect 3426 2116 3429 2163
rect 3418 2113 3429 2116
rect 3418 2006 3421 2113
rect 3418 2003 3429 2006
rect 3394 1903 3397 1926
rect 3410 1876 3413 1996
rect 3426 1956 3429 2003
rect 3346 1873 3357 1876
rect 3314 1816 3317 1826
rect 3330 1823 3337 1826
rect 3314 1813 3325 1816
rect 3290 1793 3293 1813
rect 3298 1776 3301 1813
rect 3298 1773 3313 1776
rect 3266 1733 3277 1736
rect 3234 1723 3245 1726
rect 3226 1613 3229 1646
rect 3258 1623 3261 1726
rect 3242 1613 3261 1616
rect 3226 1556 3229 1576
rect 3226 1553 3233 1556
rect 3230 1496 3233 1553
rect 3242 1533 3245 1613
rect 3250 1526 3253 1586
rect 3226 1493 3233 1496
rect 3242 1523 3253 1526
rect 3202 1473 3213 1476
rect 3210 1356 3213 1473
rect 3226 1406 3229 1493
rect 3242 1413 3245 1523
rect 3258 1516 3261 1596
rect 3250 1513 3261 1516
rect 3202 1353 3213 1356
rect 3222 1403 3229 1406
rect 3202 1323 3205 1353
rect 3222 1336 3225 1403
rect 3234 1383 3237 1396
rect 3218 1333 3225 1336
rect 3218 1316 3221 1333
rect 3234 1326 3237 1336
rect 3242 1333 3245 1406
rect 3214 1313 3221 1316
rect 3214 1256 3217 1313
rect 3226 1266 3229 1326
rect 3234 1323 3245 1326
rect 3226 1263 3233 1266
rect 3214 1253 3221 1256
rect 3194 1133 3197 1156
rect 3202 1133 3205 1236
rect 3210 1223 3213 1236
rect 3210 1136 3213 1206
rect 3218 1143 3221 1253
rect 3230 1196 3233 1263
rect 3242 1233 3245 1323
rect 3242 1213 3245 1226
rect 3230 1193 3237 1196
rect 3210 1133 3221 1136
rect 3186 1016 3189 1106
rect 3170 1013 3189 1016
rect 3154 993 3157 1006
rect 3162 983 3165 1006
rect 3170 933 3181 936
rect 3186 933 3189 1013
rect 3202 1006 3205 1126
rect 3202 1003 3213 1006
rect 3122 893 3133 896
rect 3130 836 3133 893
rect 3170 836 3173 933
rect 3194 923 3197 956
rect 3122 833 3133 836
rect 3162 833 3173 836
rect 3114 736 3117 746
rect 3098 733 3117 736
rect 3086 723 3093 726
rect 3090 523 3093 723
rect 3114 646 3117 716
rect 3106 643 3117 646
rect 3098 533 3101 616
rect 3106 506 3109 643
rect 3122 626 3125 833
rect 3146 803 3149 826
rect 3118 623 3125 626
rect 3118 536 3121 623
rect 3118 533 3125 536
rect 3130 533 3133 756
rect 3138 603 3141 776
rect 3162 756 3165 833
rect 3162 753 3173 756
rect 3146 733 3157 736
rect 3146 696 3149 733
rect 3162 713 3165 736
rect 3146 693 3157 696
rect 3154 636 3157 693
rect 3146 633 3157 636
rect 3146 613 3149 633
rect 3170 623 3173 753
rect 3178 696 3181 826
rect 3202 816 3205 986
rect 3210 923 3213 1003
rect 3218 906 3221 1133
rect 3226 1116 3229 1126
rect 3234 1123 3237 1193
rect 3250 1126 3253 1513
rect 3266 1506 3269 1656
rect 3274 1633 3277 1733
rect 3282 1643 3285 1736
rect 3290 1706 3293 1726
rect 3290 1703 3301 1706
rect 3298 1646 3301 1703
rect 3290 1643 3301 1646
rect 3310 1646 3313 1773
rect 3322 1733 3325 1813
rect 3334 1766 3337 1823
rect 3354 1776 3357 1873
rect 3330 1763 3337 1766
rect 3346 1773 3357 1776
rect 3402 1873 3413 1876
rect 3418 1953 3429 1956
rect 3402 1776 3405 1873
rect 3418 1856 3421 1953
rect 3426 1923 3429 1936
rect 3414 1853 3421 1856
rect 3414 1796 3417 1853
rect 3414 1793 3421 1796
rect 3402 1773 3413 1776
rect 3310 1643 3317 1646
rect 3290 1626 3293 1643
rect 3274 1623 3309 1626
rect 3274 1533 3277 1623
rect 3262 1503 3269 1506
rect 3262 1426 3265 1503
rect 3258 1423 3265 1426
rect 3258 1223 3261 1423
rect 3266 1386 3269 1406
rect 3274 1403 3277 1526
rect 3282 1456 3285 1616
rect 3290 1546 3293 1616
rect 3306 1613 3309 1623
rect 3298 1603 3309 1606
rect 3314 1603 3317 1643
rect 3290 1543 3301 1546
rect 3290 1513 3293 1536
rect 3298 1466 3301 1543
rect 3298 1463 3309 1466
rect 3282 1453 3293 1456
rect 3290 1413 3293 1453
rect 3306 1396 3309 1463
rect 3322 1443 3325 1716
rect 3330 1593 3333 1763
rect 3346 1633 3349 1773
rect 3370 1713 3373 1726
rect 3370 1613 3373 1626
rect 3346 1573 3349 1606
rect 3338 1533 3341 1546
rect 3354 1533 3373 1536
rect 3338 1523 3349 1526
rect 3354 1506 3357 1533
rect 3346 1503 3357 1506
rect 3346 1426 3349 1503
rect 3346 1423 3357 1426
rect 3354 1406 3357 1423
rect 3362 1413 3365 1526
rect 3370 1493 3373 1526
rect 3378 1436 3381 1666
rect 3386 1533 3397 1536
rect 3378 1433 3385 1436
rect 3370 1413 3373 1426
rect 3274 1393 3309 1396
rect 3266 1383 3277 1386
rect 3282 1383 3285 1393
rect 3274 1336 3277 1383
rect 3258 1203 3261 1216
rect 3266 1176 3269 1336
rect 3274 1333 3293 1336
rect 3298 1333 3301 1386
rect 3274 1313 3277 1326
rect 3258 1173 3269 1176
rect 3274 1146 3277 1226
rect 3282 1213 3285 1246
rect 3290 1213 3293 1316
rect 3266 1143 3277 1146
rect 3250 1123 3257 1126
rect 3226 1113 3245 1116
rect 3226 1023 3229 1086
rect 3226 983 3229 1016
rect 3234 993 3237 1006
rect 3242 1003 3245 1113
rect 3254 1076 3257 1123
rect 3266 1083 3269 1143
rect 3274 1113 3277 1136
rect 3254 1073 3269 1076
rect 3250 1013 3261 1016
rect 3258 993 3261 1006
rect 3266 986 3269 1073
rect 3290 1026 3293 1136
rect 3298 1123 3301 1326
rect 3314 1226 3317 1326
rect 3338 1323 3341 1406
rect 3354 1403 3365 1406
rect 3362 1393 3365 1403
rect 3362 1333 3365 1346
rect 3370 1316 3373 1406
rect 3382 1346 3385 1433
rect 3394 1403 3397 1526
rect 3402 1513 3405 1536
rect 3410 1453 3413 1773
rect 3418 1706 3421 1793
rect 3426 1723 3429 1916
rect 3418 1703 3425 1706
rect 3422 1636 3425 1703
rect 3418 1633 3425 1636
rect 3418 1526 3421 1633
rect 3426 1543 3429 1616
rect 3434 1533 3437 1906
rect 3418 1523 3425 1526
rect 3366 1313 3373 1316
rect 3378 1343 3385 1346
rect 3402 1343 3405 1426
rect 3410 1403 3413 1446
rect 3314 1223 3333 1226
rect 3314 1203 3317 1223
rect 3314 1113 3317 1126
rect 3314 1086 3317 1106
rect 3306 1083 3317 1086
rect 3322 1086 3325 1186
rect 3338 1103 3341 1226
rect 3346 1213 3349 1226
rect 3354 1223 3357 1236
rect 3366 1206 3369 1313
rect 3366 1203 3373 1206
rect 3370 1183 3373 1203
rect 3378 1136 3381 1343
rect 3394 1333 3405 1336
rect 3386 1233 3389 1326
rect 3402 1233 3405 1333
rect 3410 1323 3413 1396
rect 3422 1316 3425 1523
rect 3418 1313 3425 1316
rect 3386 1196 3389 1216
rect 3394 1213 3397 1226
rect 3410 1213 3413 1226
rect 3418 1196 3421 1313
rect 3386 1193 3397 1196
rect 3322 1083 3333 1086
rect 3306 1036 3309 1083
rect 3306 1033 3317 1036
rect 3242 983 3269 986
rect 3242 943 3245 983
rect 3242 923 3245 936
rect 3266 923 3269 946
rect 3218 903 3229 906
rect 3226 826 3229 903
rect 3274 896 3277 1026
rect 3286 1023 3293 1026
rect 3286 936 3289 1023
rect 3266 893 3277 896
rect 3282 933 3289 936
rect 3226 823 3245 826
rect 3202 813 3221 816
rect 3202 806 3205 813
rect 3186 743 3189 806
rect 3194 803 3205 806
rect 3194 716 3197 803
rect 3202 736 3205 796
rect 3226 753 3229 806
rect 3242 776 3245 823
rect 3266 803 3269 893
rect 3282 876 3285 933
rect 3290 886 3293 926
rect 3298 893 3301 1016
rect 3314 1013 3317 1033
rect 3330 1026 3333 1083
rect 3322 1023 3333 1026
rect 3306 986 3309 1006
rect 3306 983 3313 986
rect 3310 906 3313 983
rect 3322 923 3325 1023
rect 3338 946 3341 996
rect 3346 983 3349 1136
rect 3374 1133 3381 1136
rect 3330 943 3341 946
rect 3338 933 3357 936
rect 3310 903 3317 906
rect 3290 883 3301 886
rect 3278 873 3285 876
rect 3238 773 3245 776
rect 3266 773 3269 796
rect 3202 733 3221 736
rect 3226 723 3229 746
rect 3194 713 3229 716
rect 3178 693 3189 696
rect 3186 636 3189 693
rect 3226 643 3229 713
rect 3238 706 3241 773
rect 3266 713 3269 766
rect 3278 756 3281 873
rect 3290 813 3293 836
rect 3290 773 3293 806
rect 3278 753 3285 756
rect 3238 703 3245 706
rect 3242 646 3245 703
rect 3234 643 3245 646
rect 3178 633 3189 636
rect 3178 616 3181 633
rect 3170 546 3173 616
rect 3178 613 3189 616
rect 3178 583 3181 606
rect 3194 603 3197 616
rect 3202 593 3205 616
rect 3234 613 3237 643
rect 3146 543 3173 546
rect 3122 513 3125 533
rect 3130 506 3133 526
rect 3074 503 3085 506
rect 3106 503 3133 506
rect 3082 426 3085 503
rect 3138 476 3141 536
rect 3146 513 3149 543
rect 3154 523 3157 536
rect 3194 516 3197 536
rect 3218 533 3221 546
rect 3242 526 3245 536
rect 3186 513 3197 516
rect 3138 473 3149 476
rect 3146 456 3149 473
rect 3186 456 3189 513
rect 3146 453 3153 456
rect 3074 423 3085 426
rect 2986 333 2989 346
rect 3010 343 3021 346
rect 2938 263 2941 326
rect 3018 296 3021 343
rect 3034 323 3037 413
rect 3058 393 3061 406
rect 3074 383 3077 423
rect 3082 353 3085 406
rect 3122 383 3125 406
rect 3150 396 3153 453
rect 3170 453 3189 456
rect 3146 393 3153 396
rect 3098 333 3101 346
rect 3010 293 3021 296
rect 3010 236 3013 293
rect 2874 193 2877 206
rect 2890 203 2893 216
rect 2906 213 2925 216
rect 2754 153 2789 156
rect 2754 133 2757 153
rect 2834 143 2869 146
rect 2834 133 2837 143
rect 2842 133 2861 136
rect 2778 113 2781 126
rect 2850 103 2853 126
rect 2858 106 2861 133
rect 2866 123 2869 143
rect 2874 113 2877 136
rect 2890 126 2893 136
rect 2882 123 2893 126
rect 2882 106 2885 123
rect 2898 113 2901 206
rect 2930 196 2933 226
rect 2938 203 2941 236
rect 2978 233 3013 236
rect 2922 193 2933 196
rect 2922 146 2925 193
rect 2922 143 2933 146
rect 2930 123 2933 143
rect 2858 103 2885 106
rect 2938 106 2941 196
rect 2962 156 2965 226
rect 2978 203 2981 233
rect 3066 223 3069 326
rect 3146 323 3149 393
rect 3162 366 3165 426
rect 3170 413 3173 453
rect 3202 436 3205 526
rect 3234 523 3245 526
rect 3234 516 3237 523
rect 3210 513 3237 516
rect 3250 513 3253 626
rect 3266 603 3277 606
rect 3258 533 3261 546
rect 3266 516 3269 603
rect 3282 583 3285 753
rect 3298 696 3301 883
rect 3314 756 3317 903
rect 3338 803 3341 933
rect 3346 913 3349 926
rect 3362 893 3365 1106
rect 3374 1046 3377 1133
rect 3394 1126 3397 1193
rect 3386 1123 3397 1126
rect 3410 1193 3421 1196
rect 3410 1126 3413 1193
rect 3410 1123 3421 1126
rect 3374 1043 3381 1046
rect 3386 1043 3389 1123
rect 3370 1013 3373 1026
rect 3346 813 3349 836
rect 3346 796 3349 806
rect 3330 793 3349 796
rect 3362 793 3365 806
rect 3306 753 3317 756
rect 3306 723 3309 753
rect 3338 733 3349 736
rect 3354 733 3357 746
rect 3314 703 3317 716
rect 3322 713 3325 726
rect 3298 693 3313 696
rect 3310 636 3313 693
rect 3298 623 3301 636
rect 3310 633 3317 636
rect 3262 513 3269 516
rect 3262 436 3265 513
rect 3274 446 3277 526
rect 3298 503 3301 606
rect 3306 533 3309 616
rect 3306 513 3309 526
rect 3274 443 3281 446
rect 3202 433 3213 436
rect 3262 433 3269 436
rect 3202 413 3205 426
rect 3162 363 3169 366
rect 3166 286 3169 363
rect 3210 356 3213 433
rect 3234 383 3237 406
rect 3258 393 3261 416
rect 3202 353 3213 356
rect 3162 283 3169 286
rect 3026 203 3029 216
rect 3074 203 3077 216
rect 3090 203 3093 236
rect 3098 193 3101 206
rect 3162 203 3165 283
rect 3178 246 3181 326
rect 3202 306 3205 353
rect 3226 333 3229 346
rect 3266 323 3269 433
rect 3278 376 3281 443
rect 3274 373 3281 376
rect 3274 313 3277 373
rect 3170 243 3181 246
rect 3170 193 3173 243
rect 3178 223 3181 236
rect 3186 186 3189 306
rect 3202 303 3221 306
rect 3194 193 3197 236
rect 3202 206 3205 226
rect 3202 203 3213 206
rect 3186 183 3197 186
rect 2962 153 2989 156
rect 2962 113 2965 126
rect 2970 106 2973 126
rect 2938 103 2973 106
rect 2986 103 2989 153
rect 3058 133 3061 146
rect 3074 133 3077 156
rect 3066 123 3085 126
rect 3090 123 3093 146
rect 3106 133 3109 176
rect 3146 133 3149 156
rect 3194 133 3197 183
rect 3218 173 3221 303
rect 3226 153 3229 216
rect 3242 136 3245 286
rect 3306 283 3309 326
rect 3314 296 3317 633
rect 3322 613 3325 646
rect 3338 633 3341 726
rect 3346 603 3349 726
rect 3354 703 3357 726
rect 3362 713 3365 726
rect 3370 626 3373 936
rect 3378 786 3381 1043
rect 3386 1013 3389 1036
rect 3386 813 3389 946
rect 3402 916 3405 1106
rect 3418 1036 3421 1123
rect 3426 1113 3429 1236
rect 3414 1033 3421 1036
rect 3414 936 3417 1033
rect 3414 933 3421 936
rect 3402 913 3413 916
rect 3402 893 3405 906
rect 3402 813 3405 836
rect 3386 803 3397 806
rect 3378 783 3389 786
rect 3386 636 3389 783
rect 3410 733 3413 856
rect 3418 836 3421 933
rect 3426 853 3429 1026
rect 3418 833 3425 836
rect 3410 706 3413 726
rect 3354 623 3373 626
rect 3322 513 3325 536
rect 3354 526 3357 623
rect 3362 606 3365 616
rect 3370 613 3373 623
rect 3378 633 3389 636
rect 3402 703 3413 706
rect 3402 636 3405 703
rect 3422 696 3425 833
rect 3418 693 3425 696
rect 3402 633 3413 636
rect 3362 603 3373 606
rect 3330 516 3333 526
rect 3338 523 3357 526
rect 3330 513 3357 516
rect 3362 413 3365 536
rect 3370 533 3373 603
rect 3378 586 3381 633
rect 3386 603 3389 616
rect 3378 583 3389 586
rect 3386 536 3389 583
rect 3378 533 3389 536
rect 3378 513 3381 533
rect 3402 523 3405 616
rect 3410 613 3413 633
rect 3410 583 3413 606
rect 3418 566 3421 693
rect 3414 563 3421 566
rect 3414 506 3417 563
rect 3426 513 3429 606
rect 3434 543 3437 1456
rect 3370 486 3373 506
rect 3410 503 3417 506
rect 3370 483 3381 486
rect 3378 406 3381 483
rect 3338 383 3341 406
rect 3362 403 3381 406
rect 3410 406 3413 503
rect 3426 413 3429 506
rect 3410 403 3421 406
rect 3362 346 3365 403
rect 3418 363 3421 403
rect 3338 333 3341 346
rect 3362 343 3373 346
rect 3314 293 3325 296
rect 3322 236 3325 293
rect 3338 266 3341 316
rect 3370 296 3373 343
rect 3386 323 3389 336
rect 3434 333 3437 536
rect 3362 293 3373 296
rect 3338 263 3349 266
rect 3266 233 3325 236
rect 3266 203 3269 233
rect 3322 213 3341 216
rect 3226 133 3245 136
rect 3178 123 3245 126
rect 3082 116 3085 123
rect 3250 116 3253 156
rect 3314 133 3317 206
rect 3322 193 3325 206
rect 3330 193 3333 206
rect 3322 133 3325 156
rect 3346 133 3349 263
rect 3362 203 3365 293
rect 3418 236 3421 326
rect 3370 233 3421 236
rect 3370 136 3373 233
rect 3354 133 3373 136
rect 3330 123 3373 126
rect 3082 113 3109 116
rect 3242 113 3253 116
rect 3378 113 3381 156
rect 3426 133 3429 206
rect 3434 203 3437 216
rect 2594 93 2621 96
rect 2402 73 2429 76
rect 3446 37 3466 3303
rect 3470 13 3490 3327
<< metal3 >>
rect 649 3272 1326 3277
rect 1361 3262 1854 3267
rect 2793 3262 2918 3267
rect 1041 3252 1286 3257
rect 609 3242 686 3247
rect 825 3242 950 3247
rect 825 3237 830 3242
rect 617 3232 662 3237
rect 801 3232 830 3237
rect 945 3237 950 3242
rect 1041 3237 1046 3252
rect 1281 3247 1286 3252
rect 2201 3252 2310 3257
rect 2201 3247 2206 3252
rect 1281 3242 1358 3247
rect 1857 3242 2094 3247
rect 2177 3242 2206 3247
rect 2305 3247 2310 3252
rect 2449 3252 2718 3257
rect 2305 3242 2334 3247
rect 1129 3237 1230 3242
rect 2449 3237 2454 3252
rect 2713 3237 2718 3252
rect 945 3232 1046 3237
rect 1065 3232 1134 3237
rect 1225 3232 1366 3237
rect 1417 3232 1502 3237
rect 2081 3232 2262 3237
rect 2425 3232 2454 3237
rect 2489 3232 2694 3237
rect 2713 3232 2742 3237
rect 2857 3232 2998 3237
rect 3073 3232 3278 3237
rect 2489 3227 2494 3232
rect 841 3222 990 3227
rect 1145 3222 1542 3227
rect 1561 3222 1662 3227
rect 1681 3222 1774 3227
rect 1817 3222 1926 3227
rect 2041 3222 2110 3227
rect 2321 3222 2438 3227
rect 2465 3222 2494 3227
rect 2689 3227 2694 3232
rect 2689 3222 2870 3227
rect 1561 3217 1566 3222
rect 553 3212 630 3217
rect 721 3212 1214 3217
rect 1225 3212 1318 3217
rect 1345 3212 1566 3217
rect 1657 3217 1662 3222
rect 2433 3217 2438 3222
rect 1657 3212 1878 3217
rect 2033 3212 2174 3217
rect 2265 3212 2342 3217
rect 2433 3212 2806 3217
rect 1897 3207 2014 3212
rect 3073 3207 3078 3232
rect 3273 3217 3278 3232
rect 3273 3212 3382 3217
rect 329 3202 390 3207
rect 737 3202 910 3207
rect 1121 3202 1342 3207
rect 1473 3202 1902 3207
rect 2009 3202 2142 3207
rect 2201 3202 2518 3207
rect 2793 3202 3078 3207
rect 3089 3202 3262 3207
rect 985 3197 1102 3202
rect 1361 3197 1478 3202
rect 3089 3197 3094 3202
rect 3257 3197 3262 3202
rect 3353 3202 3382 3207
rect 3353 3197 3358 3202
rect 305 3192 422 3197
rect 529 3192 742 3197
rect 761 3192 990 3197
rect 1097 3192 1206 3197
rect 1297 3192 1366 3197
rect 1489 3192 1590 3197
rect 1601 3192 1702 3197
rect 1761 3192 1998 3197
rect 2041 3192 2134 3197
rect 2177 3192 2286 3197
rect 2321 3192 2438 3197
rect 2633 3192 2710 3197
rect 2761 3192 2782 3197
rect 2977 3192 3006 3197
rect 417 3182 502 3187
rect 737 3177 742 3192
rect 3001 3187 3006 3192
rect 3065 3192 3094 3197
rect 3105 3192 3134 3197
rect 3065 3187 3070 3192
rect 785 3182 910 3187
rect 985 3182 1142 3187
rect 1337 3182 1582 3187
rect 1729 3182 1966 3187
rect 1993 3182 2126 3187
rect 2497 3182 2814 3187
rect 3001 3182 3070 3187
rect 3129 3187 3134 3192
rect 3201 3192 3230 3197
rect 3257 3192 3358 3197
rect 3201 3187 3206 3192
rect 3129 3182 3206 3187
rect 1169 3177 1318 3182
rect 1601 3177 1734 3182
rect 217 3172 310 3177
rect 529 3172 622 3177
rect 737 3172 766 3177
rect 857 3172 902 3177
rect 913 3172 1102 3177
rect 1145 3172 1174 3177
rect 1313 3172 1430 3177
rect 1505 3172 1606 3177
rect 1753 3172 1862 3177
rect 1929 3172 2222 3177
rect 2337 3172 2422 3177
rect 2577 3172 2646 3177
rect 529 3167 534 3172
rect 361 3162 486 3167
rect 505 3162 534 3167
rect 617 3167 622 3172
rect 761 3167 862 3172
rect 897 3167 902 3172
rect 2641 3167 2646 3172
rect 2825 3172 2902 3177
rect 2825 3167 2830 3172
rect 617 3162 646 3167
rect 897 3162 1134 3167
rect 1185 3162 1406 3167
rect 1521 3162 1622 3167
rect 1673 3162 1790 3167
rect 1969 3162 2006 3167
rect 2025 3162 2334 3167
rect 2569 3162 2622 3167
rect 2641 3162 2830 3167
rect 361 3157 366 3162
rect 89 3152 302 3157
rect 337 3152 366 3157
rect 481 3157 486 3162
rect 481 3152 774 3157
rect 793 3152 894 3157
rect 921 3152 1158 3157
rect 1185 3147 1190 3162
rect 1617 3157 1622 3162
rect 1233 3152 1438 3157
rect 1617 3152 1782 3157
rect 1953 3152 2446 3157
rect 2521 3152 2606 3157
rect 3233 3152 3262 3157
rect 65 3142 270 3147
rect 377 3142 510 3147
rect 545 3142 598 3147
rect 609 3142 670 3147
rect 745 3142 1014 3147
rect 1089 3142 1190 3147
rect 1209 3142 1254 3147
rect 265 3137 382 3142
rect 593 3137 598 3142
rect 1265 3137 1270 3147
rect 1313 3142 1406 3147
rect 1545 3142 1646 3147
rect 1793 3142 1822 3147
rect 1985 3142 2342 3147
rect 2353 3142 2462 3147
rect 2849 3142 2934 3147
rect 2969 3142 3062 3147
rect 1641 3137 1798 3142
rect 2353 3137 2358 3142
rect 137 3132 246 3137
rect 409 3132 526 3137
rect 593 3132 718 3137
rect 753 3132 1022 3137
rect 1121 3132 1374 3137
rect 1473 3132 1542 3137
rect 1921 3132 2062 3137
rect 2305 3132 2358 3137
rect 2369 3132 2534 3137
rect 2681 3132 2774 3137
rect 2865 3132 2902 3137
rect 2977 3132 3134 3137
rect 2185 3127 2286 3132
rect 2865 3127 2870 3132
rect 281 3122 470 3127
rect 617 3122 1142 3127
rect 1273 3122 1334 3127
rect 1401 3122 1606 3127
rect 1625 3122 1702 3127
rect 497 3117 598 3122
rect 1625 3117 1630 3122
rect 329 3112 358 3117
rect 353 3107 358 3112
rect 473 3112 502 3117
rect 593 3112 758 3117
rect 833 3112 926 3117
rect 1025 3112 1294 3117
rect 1521 3112 1630 3117
rect 1697 3117 1702 3122
rect 1745 3122 1846 3127
rect 1865 3122 2022 3127
rect 2161 3122 2190 3127
rect 2281 3122 2446 3127
rect 2481 3122 2638 3127
rect 2689 3122 2870 3127
rect 2889 3122 2966 3127
rect 3033 3122 3062 3127
rect 1745 3117 1750 3122
rect 1697 3112 1750 3117
rect 1841 3117 1846 3122
rect 2961 3117 3038 3122
rect 1841 3112 2070 3117
rect 2209 3112 2630 3117
rect 3233 3112 3238 3152
rect 3281 3112 3342 3117
rect 473 3107 478 3112
rect 833 3107 838 3112
rect 1025 3107 1030 3112
rect 1313 3107 1462 3112
rect 353 3102 478 3107
rect 497 3102 566 3107
rect 577 3102 638 3107
rect 649 3102 838 3107
rect 865 3102 1030 3107
rect 1113 3102 1318 3107
rect 1457 3102 1686 3107
rect 1737 3102 2150 3107
rect 2249 3102 2502 3107
rect 2593 3102 2718 3107
rect 2737 3102 2934 3107
rect 505 3092 1206 3097
rect 1217 3092 1574 3097
rect 1593 3092 1814 3097
rect 1825 3092 1966 3097
rect 2081 3092 2126 3097
rect 1201 3087 1206 3092
rect 1569 3087 1574 3092
rect 273 3082 494 3087
rect 489 3077 494 3082
rect 601 3082 630 3087
rect 649 3082 678 3087
rect 849 3082 918 3087
rect 1201 3082 1542 3087
rect 1569 3082 1686 3087
rect 1809 3082 1814 3092
rect 2145 3087 2150 3102
rect 2737 3097 2742 3102
rect 2225 3092 2358 3097
rect 2385 3092 2566 3097
rect 2713 3092 2742 3097
rect 2929 3097 2934 3102
rect 2977 3102 3086 3107
rect 2977 3097 2982 3102
rect 2929 3092 2982 3097
rect 3081 3097 3086 3102
rect 3081 3092 3270 3097
rect 2561 3087 2662 3092
rect 2145 3082 2382 3087
rect 2657 3082 2918 3087
rect 601 3077 606 3082
rect 489 3072 606 3077
rect 673 3077 678 3082
rect 745 3077 854 3082
rect 1809 3077 1894 3082
rect 2913 3077 2918 3082
rect 2993 3082 3070 3087
rect 2993 3077 2998 3082
rect 673 3072 750 3077
rect 985 3072 1414 3077
rect 1889 3072 2134 3077
rect 2249 3072 2278 3077
rect 2617 3072 2646 3077
rect 2129 3067 2254 3072
rect 2641 3067 2646 3072
rect 2865 3072 2894 3077
rect 2913 3072 2998 3077
rect 2865 3067 2870 3072
rect 769 3062 974 3067
rect 1241 3062 1462 3067
rect 1497 3062 1878 3067
rect 2361 3062 2582 3067
rect 2641 3062 2870 3067
rect 969 3057 1158 3062
rect 1241 3057 1246 3062
rect 385 3052 638 3057
rect 657 3052 806 3057
rect 1153 3052 1246 3057
rect 1265 3052 1534 3057
rect 1713 3052 1926 3057
rect 2105 3052 2190 3057
rect 3185 3052 3350 3057
rect 385 3047 390 3052
rect 233 3042 390 3047
rect 633 3047 638 3052
rect 633 3042 1022 3047
rect 1081 3042 1134 3047
rect 1377 3042 1638 3047
rect 1705 3042 1750 3047
rect 2041 3042 2110 3047
rect 2345 3042 2374 3047
rect 1265 3037 1358 3042
rect 593 3032 670 3037
rect 705 3032 838 3037
rect 1097 3032 1270 3037
rect 1353 3032 1502 3037
rect 1577 3032 1646 3037
rect 1705 3032 1758 3037
rect 1809 3032 1854 3037
rect 1993 3032 2126 3037
rect 2177 3032 2238 3037
rect 2329 3032 2374 3037
rect 2409 3032 2574 3037
rect 2657 3032 2742 3037
rect 865 3027 966 3032
rect 2369 3027 2374 3032
rect 401 3022 494 3027
rect 553 3022 590 3027
rect 649 3022 742 3027
rect 777 3022 830 3027
rect 841 3022 870 3027
rect 961 3022 990 3027
rect 1073 3022 1150 3027
rect 1281 3022 1310 3027
rect 1329 3022 1422 3027
rect 1433 3022 1606 3027
rect 1665 3022 1870 3027
rect 1953 3022 2158 3027
rect 2169 3022 2350 3027
rect 2369 3022 2430 3027
rect 2649 3022 2798 3027
rect 2969 3022 3158 3027
rect 3217 3022 3294 3027
rect 1393 3017 1398 3022
rect 353 3012 390 3017
rect 689 3012 1358 3017
rect 1393 3012 1574 3017
rect 1593 3012 2286 3017
rect 2553 3012 2758 3017
rect 385 3007 390 3012
rect 2553 3007 2558 3012
rect 2969 3007 2974 3022
rect 137 3002 214 3007
rect 385 3002 406 3007
rect 689 3002 726 3007
rect 785 3002 1022 3007
rect 1057 3002 1558 3007
rect 1625 3002 1950 3007
rect 2009 3002 2070 3007
rect 2121 3002 2246 3007
rect 2433 3002 2558 3007
rect 2641 3002 2918 3007
rect 2945 3002 2974 3007
rect 3153 3007 3158 3022
rect 3153 3002 3182 3007
rect 3313 3002 3398 3007
rect 3313 2997 3318 3002
rect 137 2992 230 2997
rect 249 2992 358 2997
rect 521 2992 598 2997
rect 673 2992 750 2997
rect 801 2992 854 2997
rect 1009 2992 1134 2997
rect 1201 2992 1494 2997
rect 1569 2992 1790 2997
rect 1841 2992 2166 2997
rect 2289 2992 2326 2997
rect 2489 2992 2710 2997
rect 1489 2987 1574 2992
rect 2161 2987 2166 2992
rect 2705 2987 2710 2992
rect 2929 2992 3014 2997
rect 3041 2992 3142 2997
rect 3249 2992 3318 2997
rect 3393 2997 3398 3002
rect 3393 2992 3422 2997
rect 2929 2987 2934 2992
rect 537 2982 726 2987
rect 817 2982 998 2987
rect 1081 2982 1254 2987
rect 1345 2982 1430 2987
rect 1721 2982 1982 2987
rect 2017 2982 2150 2987
rect 2161 2982 2630 2987
rect 2705 2982 2934 2987
rect 3049 2982 3078 2987
rect 3169 2982 3198 2987
rect 993 2977 1086 2982
rect 3073 2977 3174 2982
rect 193 2972 294 2977
rect 561 2972 798 2977
rect 1105 2972 1214 2977
rect 1305 2972 1414 2977
rect 1441 2972 1550 2977
rect 1929 2972 2046 2977
rect 2097 2972 2318 2977
rect 2521 2972 2582 2977
rect 3313 2972 3382 2977
rect 2097 2967 2102 2972
rect 2313 2967 2526 2972
rect 545 2962 622 2967
rect 681 2962 798 2967
rect 817 2962 886 2967
rect 969 2962 1158 2967
rect 1337 2962 1422 2967
rect 1657 2962 1758 2967
rect 1785 2962 1822 2967
rect 1865 2962 2102 2967
rect 2169 2962 2246 2967
rect 2545 2962 2686 2967
rect 2993 2962 3094 2967
rect 817 2957 822 2962
rect 569 2952 822 2957
rect 881 2957 886 2962
rect 881 2952 910 2957
rect 1033 2952 1878 2957
rect 1937 2952 2102 2957
rect 2217 2952 2254 2957
rect 2353 2952 2510 2957
rect 2593 2952 2822 2957
rect 257 2942 334 2947
rect 417 2942 526 2947
rect 609 2942 678 2947
rect 689 2942 918 2947
rect 929 2942 1014 2947
rect 1121 2942 1310 2947
rect 1337 2942 1422 2947
rect 1441 2942 1462 2947
rect 1601 2942 1734 2947
rect 913 2937 918 2942
rect 1441 2937 1446 2942
rect 1873 2937 1878 2952
rect 2097 2947 2102 2952
rect 2817 2947 2822 2952
rect 2993 2947 2998 2962
rect 3089 2957 3094 2962
rect 3089 2952 3158 2957
rect 3313 2952 3342 2957
rect 1897 2942 1958 2947
rect 2001 2942 2086 2947
rect 2097 2942 2166 2947
rect 2233 2942 2278 2947
rect 2537 2942 2622 2947
rect 2689 2942 2798 2947
rect 2817 2942 2998 2947
rect 3009 2942 3078 2947
rect 3089 2942 3190 2947
rect 3265 2942 3326 2947
rect 2161 2937 2166 2942
rect 265 2932 310 2937
rect 505 2932 702 2937
rect 913 2932 958 2937
rect 1105 2932 1190 2937
rect 1393 2932 1446 2937
rect 1497 2932 1614 2937
rect 1721 2932 1782 2937
rect 1873 2932 1934 2937
rect 2017 2932 2142 2937
rect 2161 2932 2230 2937
rect 2281 2932 2342 2937
rect 3033 2932 3198 2937
rect 633 2922 718 2927
rect 889 2922 1102 2927
rect 1201 2922 2358 2927
rect 2417 2922 2574 2927
rect 2857 2922 2886 2927
rect 1097 2917 1206 2922
rect 209 2912 326 2917
rect 353 2912 486 2917
rect 529 2912 646 2917
rect 785 2912 830 2917
rect 1385 2912 1510 2917
rect 1529 2912 1782 2917
rect 1969 2912 2038 2917
rect 2105 2912 2326 2917
rect 2353 2912 2358 2922
rect 2881 2917 2886 2922
rect 2993 2922 3054 2927
rect 3249 2922 3350 2927
rect 2993 2917 2998 2922
rect 2881 2912 2998 2917
rect 3057 2912 3110 2917
rect 353 2907 358 2912
rect 297 2902 358 2907
rect 481 2907 486 2912
rect 993 2907 1078 2912
rect 1505 2907 1510 2912
rect 481 2902 606 2907
rect 657 2902 782 2907
rect 777 2897 782 2902
rect 889 2902 918 2907
rect 969 2902 998 2907
rect 1073 2902 1174 2907
rect 889 2897 894 2902
rect 1169 2897 1174 2902
rect 1305 2902 1334 2907
rect 1505 2902 1550 2907
rect 1569 2902 1662 2907
rect 1305 2897 1310 2902
rect 369 2892 534 2897
rect 777 2892 894 2897
rect 961 2892 1062 2897
rect 1169 2892 1310 2897
rect 1657 2897 1662 2902
rect 1793 2902 1870 2907
rect 2177 2902 2230 2907
rect 2241 2902 2430 2907
rect 1793 2897 1798 2902
rect 2241 2897 2246 2902
rect 1657 2892 1798 2897
rect 2201 2892 2246 2897
rect 2289 2892 2406 2897
rect 2497 2892 2590 2897
rect 2609 2892 2662 2897
rect 3017 2892 3166 2897
rect 2497 2887 2502 2892
rect 913 2882 1006 2887
rect 1057 2882 1142 2887
rect 1329 2882 1374 2887
rect 1905 2882 2158 2887
rect 2321 2882 2502 2887
rect 2585 2887 2590 2892
rect 2585 2882 2638 2887
rect 2681 2882 2814 2887
rect 2833 2882 2878 2887
rect 2897 2882 2998 2887
rect 1905 2877 1910 2882
rect 1065 2872 1150 2877
rect 1441 2872 1910 2877
rect 2153 2877 2158 2882
rect 2681 2877 2686 2882
rect 2153 2872 2334 2877
rect 321 2862 1094 2867
rect 1441 2847 1446 2872
rect 2329 2867 2334 2872
rect 2425 2872 2686 2877
rect 2809 2877 2814 2882
rect 2897 2877 2902 2882
rect 2809 2872 2862 2877
rect 2881 2872 2902 2877
rect 2993 2877 2998 2882
rect 2993 2872 3342 2877
rect 2425 2867 2430 2872
rect 2881 2867 2886 2872
rect 1713 2862 1742 2867
rect 993 2842 1046 2847
rect 1193 2842 1446 2847
rect 1737 2847 1742 2862
rect 1921 2862 2190 2867
rect 2329 2862 2430 2867
rect 2657 2862 2886 2867
rect 1921 2847 1926 2862
rect 2449 2857 2662 2862
rect 2233 2852 2310 2857
rect 2449 2847 2454 2857
rect 2681 2852 3118 2857
rect 1737 2842 1926 2847
rect 1945 2842 2454 2847
rect 2465 2842 2670 2847
rect 2769 2842 2862 2847
rect 2929 2842 3006 2847
rect 641 2832 838 2837
rect 345 2822 446 2827
rect 457 2822 630 2827
rect 641 2817 646 2832
rect 833 2827 838 2832
rect 881 2832 950 2837
rect 881 2827 886 2832
rect 833 2822 886 2827
rect 945 2827 950 2832
rect 1193 2827 1198 2842
rect 2449 2837 2454 2842
rect 2665 2837 2774 2842
rect 2057 2832 2150 2837
rect 2449 2832 2478 2837
rect 2817 2832 2870 2837
rect 945 2822 1198 2827
rect 1473 2822 1598 2827
rect 1473 2817 1478 2822
rect 497 2812 646 2817
rect 665 2812 734 2817
rect 809 2812 958 2817
rect 1209 2812 1478 2817
rect 1593 2817 1598 2822
rect 1641 2822 1718 2827
rect 2073 2822 2198 2827
rect 2249 2822 2366 2827
rect 2417 2822 2558 2827
rect 2601 2822 2630 2827
rect 1641 2817 1646 2822
rect 1593 2812 1646 2817
rect 1713 2817 1718 2822
rect 2625 2817 2630 2822
rect 2737 2822 3014 2827
rect 3313 2822 3366 2827
rect 2737 2817 2742 2822
rect 1713 2812 2398 2817
rect 2393 2807 2398 2812
rect 2489 2812 2534 2817
rect 2625 2812 2742 2817
rect 2761 2812 2870 2817
rect 2489 2807 2494 2812
rect 577 2802 662 2807
rect 689 2802 942 2807
rect 1641 2802 1726 2807
rect 1849 2802 1910 2807
rect 1985 2802 2062 2807
rect 2225 2802 2310 2807
rect 2393 2802 2494 2807
rect 2529 2797 2534 2812
rect 729 2792 838 2797
rect 977 2792 1046 2797
rect 1161 2792 1254 2797
rect 1489 2792 1614 2797
rect 2529 2792 2830 2797
rect 2937 2792 3046 2797
rect 3145 2792 3366 2797
rect 449 2782 478 2787
rect 793 2782 902 2787
rect 1025 2782 1086 2787
rect 1977 2782 2030 2787
rect 2409 2782 2502 2787
rect 3081 2782 3198 2787
rect 137 2772 422 2777
rect 793 2767 886 2772
rect 609 2762 718 2767
rect 609 2757 614 2762
rect 529 2752 614 2757
rect 713 2757 718 2762
rect 769 2762 798 2767
rect 881 2762 910 2767
rect 1113 2762 1950 2767
rect 2289 2762 2390 2767
rect 769 2757 774 2762
rect 713 2752 774 2757
rect 905 2757 910 2762
rect 2289 2757 2294 2762
rect 905 2752 966 2757
rect 2265 2752 2294 2757
rect 2385 2757 2390 2762
rect 2449 2762 2518 2767
rect 2449 2757 2454 2762
rect 2385 2752 2454 2757
rect 2513 2757 2518 2762
rect 2561 2762 2630 2767
rect 2561 2757 2566 2762
rect 2513 2752 2566 2757
rect 2625 2757 2630 2762
rect 2625 2752 3342 2757
rect 1281 2747 1374 2752
rect 785 2742 894 2747
rect 1089 2742 1246 2747
rect 1257 2742 1286 2747
rect 1369 2742 1398 2747
rect 2065 2742 2214 2747
rect 2313 2742 2358 2747
rect 2465 2742 2606 2747
rect 2065 2737 2070 2742
rect 625 2732 726 2737
rect 721 2727 726 2732
rect 841 2732 894 2737
rect 841 2727 846 2732
rect 721 2722 846 2727
rect 889 2727 894 2732
rect 977 2732 1310 2737
rect 977 2727 982 2732
rect 1305 2727 1310 2732
rect 1409 2732 2070 2737
rect 2209 2737 2214 2742
rect 2209 2732 2454 2737
rect 1409 2727 1414 2732
rect 889 2722 982 2727
rect 1041 2722 1150 2727
rect 1305 2722 1414 2727
rect 2449 2727 2454 2732
rect 2577 2732 2678 2737
rect 3033 2732 3062 2737
rect 2577 2727 2582 2732
rect 3057 2727 3062 2732
rect 3153 2732 3182 2737
rect 3153 2727 3158 2732
rect 2449 2722 2582 2727
rect 2873 2722 2966 2727
rect 3057 2722 3158 2727
rect 1257 2712 1286 2717
rect 1281 2707 1286 2712
rect 1449 2712 2414 2717
rect 1449 2707 1454 2712
rect 545 2702 702 2707
rect 1281 2702 1454 2707
rect 2409 2707 2414 2712
rect 2601 2712 2630 2717
rect 3265 2712 3422 2717
rect 2601 2707 2606 2712
rect 2409 2702 2606 2707
rect 937 2692 1070 2697
rect 1681 2692 1734 2697
rect 1577 2682 1662 2687
rect 1801 2682 1894 2687
rect 1913 2682 2390 2687
rect 1577 2677 1582 2682
rect 1137 2672 1534 2677
rect 1553 2672 1582 2677
rect 1657 2677 1662 2682
rect 1913 2677 1918 2682
rect 1657 2672 1790 2677
rect 1889 2672 1918 2677
rect 2385 2677 2390 2682
rect 2921 2682 3038 2687
rect 3057 2682 3278 2687
rect 2921 2677 2926 2682
rect 2385 2672 2926 2677
rect 3033 2677 3038 2682
rect 3033 2672 3110 2677
rect 1137 2657 1142 2672
rect 401 2652 494 2657
rect 1113 2652 1142 2657
rect 1529 2657 1534 2672
rect 1785 2667 1894 2672
rect 2073 2662 2350 2667
rect 3281 2662 3342 2667
rect 2073 2657 2078 2662
rect 1529 2652 2078 2657
rect 2345 2657 2350 2662
rect 2345 2652 2374 2657
rect 2937 2652 3054 2657
rect 401 2647 406 2652
rect 241 2642 342 2647
rect 377 2642 406 2647
rect 489 2647 494 2652
rect 2113 2647 2326 2652
rect 489 2642 518 2647
rect 705 2642 1518 2647
rect 1513 2637 1518 2642
rect 2089 2642 2118 2647
rect 2321 2642 2590 2647
rect 2609 2642 2710 2647
rect 3105 2642 3238 2647
rect 2089 2637 2094 2642
rect 2609 2637 2614 2642
rect 305 2632 566 2637
rect 1513 2632 2094 2637
rect 2113 2632 2206 2637
rect 2265 2632 2350 2637
rect 2385 2632 2422 2637
rect 2561 2632 2614 2637
rect 2705 2637 2710 2642
rect 2705 2632 2734 2637
rect 3025 2632 3150 2637
rect 193 2627 286 2632
rect 169 2622 198 2627
rect 281 2622 574 2627
rect 2449 2622 2526 2627
rect 2449 2617 2454 2622
rect 137 2612 294 2617
rect 321 2612 414 2617
rect 433 2612 462 2617
rect 289 2597 294 2612
rect 457 2607 462 2612
rect 545 2612 886 2617
rect 897 2612 2118 2617
rect 2177 2612 2350 2617
rect 2369 2612 2454 2617
rect 2521 2617 2526 2622
rect 2913 2622 2998 2627
rect 3017 2622 3134 2627
rect 3225 2622 3262 2627
rect 3329 2622 3406 2627
rect 2913 2617 2918 2622
rect 2521 2612 2918 2617
rect 2993 2617 2998 2622
rect 2993 2612 3014 2617
rect 545 2607 550 2612
rect 457 2602 550 2607
rect 881 2597 886 2612
rect 2369 2607 2374 2612
rect 3009 2607 3014 2612
rect 3073 2612 3102 2617
rect 3137 2612 3270 2617
rect 3073 2607 3078 2612
rect 1073 2602 1102 2607
rect 1529 2602 1598 2607
rect 1697 2602 1742 2607
rect 1833 2602 1902 2607
rect 2297 2602 2374 2607
rect 2441 2602 2510 2607
rect 2929 2602 2982 2607
rect 3009 2602 3078 2607
rect 1073 2597 1078 2602
rect 2161 2597 2278 2602
rect 81 2592 182 2597
rect 289 2592 390 2597
rect 881 2592 1078 2597
rect 2137 2592 2166 2597
rect 2273 2592 2598 2597
rect 2705 2592 2758 2597
rect 3241 2592 3342 2597
rect 121 2582 238 2587
rect 1273 2582 2014 2587
rect 2033 2582 2302 2587
rect 2353 2582 2950 2587
rect 3225 2582 3278 2587
rect 1273 2577 1278 2582
rect 801 2572 1206 2577
rect 1249 2572 1278 2577
rect 2009 2577 2014 2582
rect 2009 2572 2062 2577
rect 2169 2572 2782 2577
rect 1313 2567 1486 2572
rect 1737 2567 1886 2572
rect 2057 2567 2174 2572
rect 241 2562 310 2567
rect 441 2562 526 2567
rect 1153 2562 1222 2567
rect 1289 2562 1318 2567
rect 1481 2562 1742 2567
rect 1881 2562 2038 2567
rect 2193 2562 2262 2567
rect 2313 2562 2382 2567
rect 2497 2562 2734 2567
rect 2257 2557 2262 2562
rect 385 2552 902 2557
rect 913 2552 2246 2557
rect 2257 2552 2310 2557
rect 2489 2552 2574 2557
rect 2593 2552 2886 2557
rect 897 2547 902 2552
rect 2241 2547 2246 2552
rect 153 2542 222 2547
rect 457 2542 710 2547
rect 897 2542 926 2547
rect 1185 2542 2142 2547
rect 2241 2542 2822 2547
rect 2897 2542 3054 2547
rect 3073 2542 3198 2547
rect 921 2537 1190 2542
rect 2817 2537 2902 2542
rect 529 2532 662 2537
rect 801 2532 878 2537
rect 1209 2532 1310 2537
rect 1401 2532 1598 2537
rect 801 2527 806 2532
rect 137 2522 806 2527
rect 873 2527 878 2532
rect 1305 2527 1406 2532
rect 1593 2527 1598 2532
rect 1841 2532 2494 2537
rect 1841 2527 1846 2532
rect 2545 2527 2622 2532
rect 873 2522 1190 2527
rect 1209 2522 1286 2527
rect 1425 2522 1574 2527
rect 1593 2522 1846 2527
rect 1865 2522 2174 2527
rect 2281 2522 2550 2527
rect 2617 2522 2646 2527
rect 2817 2522 2950 2527
rect 1185 2517 1190 2522
rect 793 2512 974 2517
rect 1185 2512 1502 2517
rect 2049 2512 2446 2517
rect 2561 2512 2630 2517
rect 2689 2512 2758 2517
rect 2777 2512 2854 2517
rect 577 2507 774 2512
rect 233 2502 262 2507
rect 257 2497 262 2502
rect 329 2502 582 2507
rect 769 2502 1254 2507
rect 1409 2502 1438 2507
rect 1529 2502 2006 2507
rect 2017 2502 2430 2507
rect 2593 2502 2646 2507
rect 329 2497 334 2502
rect 1433 2497 1534 2502
rect 2001 2497 2006 2502
rect 2641 2497 2646 2502
rect 2785 2502 2814 2507
rect 2857 2502 3046 2507
rect 2785 2497 2790 2502
rect 257 2492 334 2497
rect 593 2492 878 2497
rect 1129 2492 1270 2497
rect 2001 2492 2054 2497
rect 2065 2492 2206 2497
rect 2401 2492 2470 2497
rect 2641 2492 2790 2497
rect 3313 2492 3422 2497
rect 897 2482 1070 2487
rect 1201 2482 1878 2487
rect 609 2477 902 2482
rect 1065 2477 1070 2482
rect 1873 2477 1878 2482
rect 1937 2482 1990 2487
rect 1937 2477 1942 2482
rect 353 2472 614 2477
rect 1065 2472 1190 2477
rect 1185 2467 1190 2472
rect 1825 2472 1854 2477
rect 1873 2472 1942 2477
rect 1825 2467 1830 2472
rect 625 2462 958 2467
rect 1009 2462 1054 2467
rect 1185 2462 1830 2467
rect 1985 2467 1990 2482
rect 2289 2482 2390 2487
rect 2289 2477 2294 2482
rect 2209 2472 2294 2477
rect 2385 2477 2390 2482
rect 2481 2482 2582 2487
rect 2481 2477 2486 2482
rect 2385 2472 2486 2477
rect 2577 2477 2582 2482
rect 3057 2482 3126 2487
rect 3057 2477 3062 2482
rect 2577 2472 3062 2477
rect 2209 2467 2214 2472
rect 1985 2462 2214 2467
rect 2313 2462 2366 2467
rect 73 2452 470 2457
rect 465 2447 470 2452
rect 681 2452 774 2457
rect 873 2452 1150 2457
rect 681 2447 686 2452
rect 769 2447 878 2452
rect 401 2442 446 2447
rect 465 2442 686 2447
rect 705 2442 750 2447
rect 1169 2442 1366 2447
rect 897 2437 1062 2442
rect 1169 2437 1174 2442
rect 873 2432 902 2437
rect 1057 2432 1174 2437
rect 1361 2437 1366 2442
rect 1409 2442 1590 2447
rect 1361 2432 1390 2437
rect 1409 2427 1414 2442
rect 689 2422 790 2427
rect 809 2422 1046 2427
rect 1185 2422 1294 2427
rect 1313 2422 1414 2427
rect 1585 2427 1590 2442
rect 1729 2442 1854 2447
rect 2233 2442 2294 2447
rect 2601 2442 2662 2447
rect 1729 2437 1734 2442
rect 1705 2432 1734 2437
rect 1849 2437 1854 2442
rect 1849 2432 1878 2437
rect 2001 2432 2886 2437
rect 3345 2432 3398 2437
rect 2881 2427 2886 2432
rect 1585 2422 2030 2427
rect 2433 2422 2806 2427
rect 2881 2422 2966 2427
rect 3129 2422 3406 2427
rect 689 2417 694 2422
rect 329 2412 694 2417
rect 785 2417 790 2422
rect 2025 2417 2166 2422
rect 2313 2417 2438 2422
rect 785 2412 1094 2417
rect 1113 2412 1174 2417
rect 1249 2412 1278 2417
rect 1353 2412 1574 2417
rect 1809 2412 2006 2417
rect 2161 2412 2318 2417
rect 1089 2407 1094 2412
rect 1169 2407 1254 2412
rect 649 2402 806 2407
rect 1089 2402 1110 2407
rect 1105 2397 1110 2402
rect 1617 2402 1686 2407
rect 2049 2402 2142 2407
rect 2337 2402 2622 2407
rect 3289 2402 3350 2407
rect 1617 2397 1622 2402
rect 97 2392 222 2397
rect 705 2392 798 2397
rect 937 2392 1094 2397
rect 1105 2392 1206 2397
rect 1249 2392 1342 2397
rect 1361 2392 1470 2397
rect 1481 2392 1622 2397
rect 1681 2397 1686 2402
rect 2337 2397 2342 2402
rect 1681 2392 1710 2397
rect 1769 2392 2342 2397
rect 2617 2397 2622 2402
rect 2617 2392 2646 2397
rect 3057 2392 3110 2397
rect 3153 2392 3270 2397
rect 2377 2387 2598 2392
rect 1097 2382 1750 2387
rect 2353 2382 2382 2387
rect 2593 2382 2694 2387
rect 2713 2382 2830 2387
rect 2097 2377 2278 2382
rect 2713 2377 2718 2382
rect 753 2372 830 2377
rect 753 2367 758 2372
rect 225 2362 398 2367
rect 577 2362 710 2367
rect 729 2362 758 2367
rect 825 2367 830 2372
rect 1041 2372 1366 2377
rect 1449 2372 1566 2377
rect 1593 2372 1654 2377
rect 1753 2372 1830 2377
rect 1849 2372 2054 2377
rect 2073 2372 2102 2377
rect 2273 2372 2598 2377
rect 2649 2372 2718 2377
rect 2825 2377 2830 2382
rect 2825 2372 2854 2377
rect 2897 2372 3022 2377
rect 825 2362 854 2367
rect 873 2362 998 2367
rect 577 2357 582 2362
rect 129 2352 254 2357
rect 553 2352 582 2357
rect 705 2357 710 2362
rect 873 2357 878 2362
rect 705 2352 878 2357
rect 993 2357 998 2362
rect 1041 2357 1046 2372
rect 1361 2367 1454 2372
rect 1649 2367 1734 2372
rect 1849 2367 1854 2372
rect 1081 2362 1182 2367
rect 1313 2362 1342 2367
rect 1473 2362 1630 2367
rect 1729 2362 1854 2367
rect 2049 2367 2054 2372
rect 2049 2362 2262 2367
rect 2385 2362 2910 2367
rect 1177 2357 1318 2362
rect 993 2352 1046 2357
rect 1089 2352 1158 2357
rect 1465 2352 2654 2357
rect 2817 2352 2846 2357
rect 2985 2352 3070 2357
rect 2985 2347 2990 2352
rect 377 2342 422 2347
rect 521 2342 566 2347
rect 601 2342 726 2347
rect 825 2342 1038 2347
rect 1193 2342 1222 2347
rect 1249 2342 1374 2347
rect 1457 2342 1494 2347
rect 1537 2342 1614 2347
rect 1641 2342 1702 2347
rect 1737 2342 1806 2347
rect 2089 2342 2790 2347
rect 2801 2342 2990 2347
rect 3065 2347 3070 2352
rect 3113 2352 3278 2357
rect 3329 2352 3350 2357
rect 3113 2347 3118 2352
rect 3065 2342 3118 2347
rect 3217 2342 3286 2347
rect 1033 2337 1198 2342
rect 1801 2337 1806 2342
rect 1905 2337 2094 2342
rect 2785 2337 2790 2342
rect 241 2332 326 2337
rect 761 2332 1014 2337
rect 1329 2332 1662 2337
rect 1801 2332 1910 2337
rect 2113 2332 2550 2337
rect 2785 2332 2854 2337
rect 3001 2332 3142 2337
rect 3153 2332 3262 2337
rect 1225 2327 1310 2332
rect 2849 2327 3006 2332
rect 201 2322 1102 2327
rect 1145 2322 1230 2327
rect 1305 2322 1782 2327
rect 1953 2322 2094 2327
rect 2569 2322 2646 2327
rect 1953 2317 1958 2322
rect 689 2312 1150 2317
rect 1241 2312 1358 2317
rect 1929 2312 1958 2317
rect 2089 2317 2094 2322
rect 2209 2317 2574 2322
rect 2641 2317 2646 2322
rect 2689 2322 2766 2327
rect 2689 2317 2694 2322
rect 2761 2317 2830 2322
rect 2089 2312 2214 2317
rect 2641 2312 2694 2317
rect 2825 2312 3094 2317
rect 425 2307 638 2312
rect 1145 2307 1246 2312
rect 1689 2307 1830 2312
rect 3089 2307 3094 2312
rect 3273 2312 3422 2317
rect 3273 2307 3278 2312
rect 401 2302 430 2307
rect 633 2302 710 2307
rect 817 2302 1126 2307
rect 1265 2302 1382 2307
rect 1457 2302 1518 2307
rect 1561 2302 1694 2307
rect 1825 2302 1958 2307
rect 1977 2302 2086 2307
rect 2225 2302 2390 2307
rect 2409 2302 2510 2307
rect 2585 2302 2630 2307
rect 2705 2302 2814 2307
rect 2905 2302 2934 2307
rect 3041 2302 3070 2307
rect 3089 2302 3278 2307
rect 3361 2302 3406 2307
rect 2929 2297 3046 2302
rect 353 2292 622 2297
rect 697 2292 902 2297
rect 913 2292 1094 2297
rect 1153 2292 1246 2297
rect 1329 2292 1550 2297
rect 1705 2292 2902 2297
rect 897 2287 902 2292
rect 1153 2287 1158 2292
rect 537 2282 766 2287
rect 897 2282 1158 2287
rect 1241 2287 1246 2292
rect 1241 2282 1502 2287
rect 1889 2282 2014 2287
rect 2233 2282 2446 2287
rect 2921 2282 3102 2287
rect 417 2277 518 2282
rect 785 2277 878 2282
rect 1681 2277 1806 2282
rect 2033 2277 2206 2282
rect 2465 2277 2646 2282
rect 2729 2277 2926 2282
rect 3097 2277 3102 2282
rect 393 2272 422 2277
rect 513 2272 790 2277
rect 873 2272 1038 2277
rect 1169 2272 1566 2277
rect 1657 2272 1686 2277
rect 1801 2272 1830 2277
rect 1953 2272 2038 2277
rect 2201 2272 2230 2277
rect 2257 2272 2470 2277
rect 2641 2272 2734 2277
rect 3097 2272 3158 2277
rect 385 2262 558 2267
rect 633 2262 1046 2267
rect 1177 2262 1446 2267
rect 1633 2262 2630 2267
rect 2745 2262 3086 2267
rect 1065 2257 1158 2262
rect 1465 2257 1614 2262
rect 2625 2257 2750 2262
rect 3081 2257 3086 2262
rect 289 2252 366 2257
rect 553 2252 702 2257
rect 713 2252 742 2257
rect 833 2252 1070 2257
rect 1153 2252 1470 2257
rect 1609 2252 1678 2257
rect 1833 2252 1862 2257
rect 2001 2252 2606 2257
rect 3081 2252 3222 2257
rect 441 2247 534 2252
rect 737 2247 838 2252
rect 1673 2247 1838 2252
rect 2769 2247 3038 2252
rect 209 2242 446 2247
rect 529 2242 614 2247
rect 857 2242 886 2247
rect 1009 2242 1302 2247
rect 1313 2242 1654 2247
rect 1977 2242 2774 2247
rect 3033 2242 3062 2247
rect 881 2237 1014 2242
rect 297 2232 390 2237
rect 457 2232 718 2237
rect 737 2232 806 2237
rect 1033 2232 1190 2237
rect 1337 2232 1374 2237
rect 1417 2232 1446 2237
rect 1505 2232 1798 2237
rect 1817 2232 2142 2237
rect 2217 2232 2278 2237
rect 2329 2232 2374 2237
rect 2513 2232 2542 2237
rect 2785 2232 2806 2237
rect 2865 2232 3030 2237
rect 3073 2232 3110 2237
rect 3321 2232 3366 2237
rect 481 2222 694 2227
rect 857 2222 918 2227
rect 1137 2222 1494 2227
rect 1001 2217 1102 2222
rect 1505 2217 1510 2232
rect 1601 2222 1638 2227
rect 1793 2222 1798 2232
rect 2585 2227 2702 2232
rect 2025 2222 2094 2227
rect 2249 2222 2294 2227
rect 2401 2222 2446 2227
rect 2481 2222 2590 2227
rect 2697 2222 2726 2227
rect 2857 2222 2934 2227
rect 2993 2222 3134 2227
rect 3153 2222 3222 2227
rect 1793 2217 1870 2222
rect 2113 2217 2230 2222
rect 2721 2217 2838 2222
rect 3153 2217 3158 2222
rect 89 2212 198 2217
rect 465 2212 750 2217
rect 897 2212 950 2217
rect 977 2212 1006 2217
rect 1097 2212 1126 2217
rect 1233 2212 1350 2217
rect 1401 2212 1510 2217
rect 1865 2212 2118 2217
rect 2225 2212 2702 2217
rect 2833 2212 3158 2217
rect 3217 2217 3222 2222
rect 3217 2212 3246 2217
rect 273 2202 614 2207
rect 665 2202 694 2207
rect 689 2197 694 2202
rect 753 2202 806 2207
rect 937 2202 1046 2207
rect 1065 2202 1230 2207
rect 1345 2202 1430 2207
rect 1713 2202 1750 2207
rect 1761 2202 1854 2207
rect 2081 2202 2334 2207
rect 2433 2202 2926 2207
rect 2961 2202 3118 2207
rect 3281 2202 3310 2207
rect 753 2197 758 2202
rect 513 2192 598 2197
rect 689 2192 758 2197
rect 777 2192 822 2197
rect 1041 2187 1046 2202
rect 1345 2197 1350 2202
rect 1105 2192 1350 2197
rect 1361 2192 1446 2197
rect 1609 2192 1710 2197
rect 1745 2192 1750 2202
rect 2081 2197 2086 2202
rect 3113 2197 3286 2202
rect 1857 2192 2086 2197
rect 2129 2192 2382 2197
rect 2441 2192 2686 2197
rect 2729 2192 2886 2197
rect 2905 2192 2998 2197
rect 3057 2192 3094 2197
rect 377 2182 550 2187
rect 1041 2182 1134 2187
rect 1161 2182 1254 2187
rect 1729 2182 1926 2187
rect 2001 2182 2030 2187
rect 569 2177 662 2182
rect 2001 2177 2006 2182
rect 497 2172 574 2177
rect 657 2172 894 2177
rect 913 2172 1022 2177
rect 1041 2172 1326 2177
rect 1553 2172 1758 2177
rect 1769 2172 2006 2177
rect 2025 2177 2030 2182
rect 2113 2182 2518 2187
rect 2617 2182 2846 2187
rect 2857 2182 2894 2187
rect 3145 2182 3254 2187
rect 3281 2182 3358 2187
rect 2113 2177 2118 2182
rect 2513 2177 2598 2182
rect 2913 2177 3086 2182
rect 2025 2172 2118 2177
rect 2137 2172 2494 2177
rect 2593 2172 2630 2177
rect 2681 2172 2918 2177
rect 3081 2172 3230 2177
rect 3321 2172 3374 2177
rect 913 2167 918 2172
rect 369 2162 646 2167
rect 745 2162 774 2167
rect 889 2162 918 2167
rect 1017 2167 1022 2172
rect 1017 2162 1070 2167
rect 1121 2162 1150 2167
rect 1257 2162 1622 2167
rect 1721 2162 1830 2167
rect 1953 2162 2006 2167
rect 2313 2162 2446 2167
rect 2545 2162 3070 2167
rect 3313 2162 3406 2167
rect 769 2157 894 2162
rect 1145 2157 1262 2162
rect 2193 2157 2294 2162
rect 241 2152 270 2157
rect 305 2152 678 2157
rect 913 2152 1078 2157
rect 1409 2152 1438 2157
rect 1505 2152 1542 2157
rect 1585 2152 1750 2157
rect 2057 2152 2094 2157
rect 2113 2152 2198 2157
rect 2289 2152 2974 2157
rect 3097 2152 3142 2157
rect 3305 2152 3414 2157
rect 1281 2147 1414 2152
rect 137 2142 214 2147
rect 353 2142 566 2147
rect 585 2142 742 2147
rect 777 2142 926 2147
rect 953 2142 982 2147
rect 1009 2142 1062 2147
rect 1081 2142 1158 2147
rect 1201 2142 1286 2147
rect 1425 2142 1630 2147
rect 1673 2142 1974 2147
rect 1993 2142 2102 2147
rect 2113 2142 2118 2152
rect 2209 2142 2382 2147
rect 2409 2142 2526 2147
rect 2545 2142 2662 2147
rect 2793 2142 3142 2147
rect 3161 2142 3334 2147
rect 233 2137 326 2142
rect 561 2137 566 2142
rect 1057 2137 1062 2142
rect 1201 2137 1206 2142
rect 1969 2137 1974 2142
rect 2129 2137 2214 2142
rect 2545 2137 2550 2142
rect 2657 2137 2774 2142
rect 177 2132 238 2137
rect 321 2132 518 2137
rect 561 2132 670 2137
rect 753 2132 926 2137
rect 993 2132 1046 2137
rect 1057 2132 1206 2137
rect 1225 2132 1270 2137
rect 1281 2132 1342 2137
rect 1353 2132 1582 2137
rect 1633 2132 1782 2137
rect 1969 2132 2134 2137
rect 2233 2132 2366 2137
rect 2465 2132 2550 2137
rect 2593 2132 2638 2137
rect 2769 2132 2862 2137
rect 2985 2132 3014 2137
rect 3113 2132 3174 2137
rect 3289 2132 3342 2137
rect 1817 2127 1950 2132
rect 2361 2127 2454 2132
rect 2857 2127 2990 2132
rect 81 2122 134 2127
rect 201 2122 310 2127
rect 489 2122 750 2127
rect 841 2122 1174 2127
rect 1193 2122 1382 2127
rect 1465 2122 1574 2127
rect 1649 2122 1822 2127
rect 1945 2122 2342 2127
rect 2449 2122 2550 2127
rect 2569 2122 2686 2127
rect 2761 2122 2822 2127
rect 3041 2122 3182 2127
rect 345 2117 454 2122
rect 1649 2117 1654 2122
rect 97 2112 198 2117
rect 265 2112 350 2117
rect 449 2112 606 2117
rect 649 2112 718 2117
rect 865 2112 1022 2117
rect 1073 2112 1478 2117
rect 1497 2112 1654 2117
rect 1665 2112 1750 2117
rect 1817 2112 1942 2117
rect 2001 2112 2110 2117
rect 2129 2112 2278 2117
rect 2337 2112 2342 2122
rect 2377 2112 2462 2117
rect 2657 2112 2686 2117
rect 2753 2112 2806 2117
rect 2865 2112 2926 2117
rect 3009 2112 3062 2117
rect 3113 2112 3190 2117
rect 3209 2112 3310 2117
rect 1073 2107 1078 2112
rect 2273 2107 2278 2112
rect 3185 2107 3190 2112
rect 113 2102 262 2107
rect 361 2102 454 2107
rect 505 2102 598 2107
rect 609 2102 702 2107
rect 865 2102 894 2107
rect 953 2102 996 2107
rect 1001 2102 1078 2107
rect 1097 2102 1190 2107
rect 1329 2102 1638 2107
rect 1729 2102 1854 2107
rect 1913 2102 2150 2107
rect 2193 2102 2238 2107
rect 2273 2102 2430 2107
rect 2441 2102 2486 2107
rect 2505 2102 2606 2107
rect 2625 2102 2678 2107
rect 2697 2102 2886 2107
rect 2897 2102 2926 2107
rect 2953 2102 3142 2107
rect 3185 2102 3398 2107
rect 991 2097 996 2102
rect 2505 2097 2510 2102
rect 89 2092 142 2097
rect 217 2092 702 2097
rect 737 2092 838 2097
rect 889 2092 982 2097
rect 991 2092 1134 2097
rect 1161 2092 1318 2097
rect 1481 2092 2510 2097
rect 2601 2097 2606 2102
rect 2881 2097 2886 2102
rect 3137 2097 3142 2102
rect 2601 2092 2782 2097
rect 2881 2092 3038 2097
rect 3137 2092 3262 2097
rect 737 2087 742 2092
rect 137 2082 542 2087
rect 601 2082 742 2087
rect 833 2087 838 2092
rect 1313 2087 1486 2092
rect 833 2082 1062 2087
rect 1121 2082 1222 2087
rect 1505 2082 1654 2087
rect 1689 2082 1742 2087
rect 1993 2082 2046 2087
rect 2057 2082 2262 2087
rect 2321 2082 2990 2087
rect 3049 2082 3198 2087
rect 1761 2077 1870 2082
rect 2985 2077 3054 2082
rect 129 2072 238 2077
rect 321 2072 1142 2077
rect 1337 2072 1382 2077
rect 1393 2072 1470 2077
rect 1489 2072 1766 2077
rect 1865 2072 2142 2077
rect 2281 2072 2342 2077
rect 2353 2072 2518 2077
rect 2641 2072 2726 2077
rect 2889 2072 2966 2077
rect 3097 2072 3166 2077
rect 233 2067 326 2072
rect 1161 2067 1318 2072
rect 1393 2067 1398 2072
rect 2161 2067 2262 2072
rect 2513 2067 2622 2072
rect 2721 2067 2894 2072
rect 345 2062 630 2067
rect 657 2062 830 2067
rect 929 2062 1166 2067
rect 1313 2062 1398 2067
rect 1441 2062 1606 2067
rect 1601 2057 1606 2062
rect 1673 2062 1798 2067
rect 1809 2062 1854 2067
rect 1937 2062 1966 2067
rect 1985 2062 2062 2067
rect 2121 2062 2166 2067
rect 2257 2062 2502 2067
rect 2617 2062 2702 2067
rect 2913 2062 2934 2067
rect 3025 2062 3094 2067
rect 1673 2057 1678 2062
rect 1809 2057 1814 2062
rect 273 2052 358 2057
rect 537 2052 958 2057
rect 977 2052 1030 2057
rect 1041 2052 1582 2057
rect 1601 2052 1678 2057
rect 1713 2052 1750 2057
rect 1761 2052 1814 2057
rect 1833 2052 2550 2057
rect 2593 2052 2934 2057
rect 2985 2052 3022 2057
rect 1025 2047 1030 2052
rect 2593 2047 2598 2052
rect 233 2042 318 2047
rect 337 2042 534 2047
rect 585 2042 758 2047
rect 793 2042 918 2047
rect 937 2042 1014 2047
rect 1025 2042 1166 2047
rect 1305 2042 1558 2047
rect 1737 2042 1790 2047
rect 1801 2042 1830 2047
rect 1841 2042 2022 2047
rect 2105 2042 2358 2047
rect 2409 2042 2446 2047
rect 2465 2042 2598 2047
rect 2617 2042 2750 2047
rect 2905 2042 2998 2047
rect 3033 2042 3286 2047
rect 1185 2037 1286 2042
rect 2993 2037 2998 2042
rect 65 2032 110 2037
rect 305 2032 638 2037
rect 673 2032 1190 2037
rect 1281 2032 1366 2037
rect 1449 2032 1478 2037
rect 1545 2032 1630 2037
rect 1721 2032 1766 2037
rect 1777 2032 1862 2037
rect 1921 2032 1958 2037
rect 1977 2032 2094 2037
rect 2145 2032 2614 2037
rect 2745 2032 2774 2037
rect 2841 2032 2966 2037
rect 2993 2032 3094 2037
rect 305 2027 310 2032
rect 1777 2027 1782 2032
rect 2145 2027 2150 2032
rect 2609 2027 2750 2032
rect 3089 2027 3094 2032
rect 3177 2032 3238 2037
rect 3177 2027 3182 2032
rect 105 2022 150 2027
rect 233 2022 270 2027
rect 281 2022 310 2027
rect 321 2022 382 2027
rect 417 2022 542 2027
rect 561 2022 654 2027
rect 681 2022 798 2027
rect 849 2022 1046 2027
rect 1057 2022 1198 2027
rect 1257 2022 1534 2027
rect 217 2012 254 2017
rect 321 2007 326 2022
rect 409 2012 486 2017
rect 665 2012 702 2017
rect 801 2012 854 2017
rect 929 2012 1278 2017
rect 697 2007 806 2012
rect 1297 2007 1406 2012
rect 105 2002 214 2007
rect 225 2002 326 2007
rect 505 2002 678 2007
rect 825 2002 1302 2007
rect 1401 2002 1430 2007
rect 225 1987 230 2002
rect 289 1992 342 1997
rect 353 1992 430 1997
rect 441 1992 574 1997
rect 769 1992 1382 1997
rect 1417 1992 1470 1997
rect 1569 1992 1574 2027
rect 1601 2022 1654 2027
rect 1681 2022 1710 2027
rect 1721 2022 1782 2027
rect 1857 2022 2150 2027
rect 2169 2022 2590 2027
rect 2945 2022 3062 2027
rect 3089 2022 3182 2027
rect 3201 2022 3302 2027
rect 1593 2012 2126 2017
rect 2305 2012 2486 2017
rect 2505 2012 2934 2017
rect 3041 2012 3070 2017
rect 2145 2007 2286 2012
rect 2929 2007 3046 2012
rect 1625 2002 1670 2007
rect 1705 2002 2150 2007
rect 2281 2002 2598 2007
rect 3233 2002 3334 2007
rect 3233 1997 3238 2002
rect 1601 1992 1766 1997
rect 1785 1992 1822 1997
rect 1841 1992 1894 1997
rect 1953 1992 1982 1997
rect 2017 1992 2526 1997
rect 2849 1992 2902 1997
rect 2945 1992 2974 1997
rect 3089 1992 3110 1997
rect 3209 1992 3238 1997
rect 3329 1997 3334 2002
rect 3329 1992 3414 1997
rect 201 1982 230 1987
rect 377 1982 414 1987
rect 561 1982 750 1987
rect 809 1982 958 1987
rect 993 1982 1046 1987
rect 1121 1982 1270 1987
rect 1481 1982 1774 1987
rect 1793 1982 2606 1987
rect 2673 1982 2838 1987
rect 433 1977 542 1982
rect 1313 1977 1486 1982
rect 305 1972 438 1977
rect 537 1972 566 1977
rect 745 1972 822 1977
rect 833 1972 870 1977
rect 897 1972 1174 1977
rect 1273 1972 1318 1977
rect 1513 1972 1654 1977
rect 1665 1972 1750 1977
rect 1777 1972 2094 1977
rect 2113 1972 2182 1977
rect 2225 1972 2286 1977
rect 2297 1972 2326 1977
rect 2401 1972 2454 1977
rect 2505 1972 2534 1977
rect 1777 1967 1782 1972
rect 2113 1967 2118 1972
rect 2177 1967 2182 1972
rect 2529 1967 2534 1972
rect 2617 1972 2710 1977
rect 2617 1967 2622 1972
rect 121 1962 246 1967
rect 377 1962 582 1967
rect 601 1962 694 1967
rect 713 1962 1078 1967
rect 1105 1962 1286 1967
rect 1361 1962 1406 1967
rect 1433 1962 1606 1967
rect 1633 1962 1782 1967
rect 1801 1962 1846 1967
rect 1857 1962 1886 1967
rect 1921 1962 2118 1967
rect 2137 1962 2166 1967
rect 2177 1962 2206 1967
rect 2249 1962 2310 1967
rect 2329 1962 2454 1967
rect 2529 1962 2622 1967
rect 2833 1967 2838 1982
rect 2961 1982 3318 1987
rect 2961 1967 2966 1982
rect 3105 1972 3158 1977
rect 2833 1962 2966 1967
rect 3153 1967 3158 1972
rect 3233 1972 3262 1977
rect 3233 1967 3238 1972
rect 3153 1962 3238 1967
rect 601 1957 606 1962
rect 345 1952 366 1957
rect 433 1952 462 1957
rect 497 1952 606 1957
rect 689 1957 694 1962
rect 689 1952 798 1957
rect 865 1952 1230 1957
rect 1345 1952 1406 1957
rect 1425 1952 1478 1957
rect 1625 1952 1726 1957
rect 1769 1952 2278 1957
rect 2297 1952 2358 1957
rect 2985 1952 3134 1957
rect 1473 1947 1630 1952
rect 105 1942 134 1947
rect 241 1942 262 1947
rect 289 1942 462 1947
rect 289 1937 294 1942
rect 457 1937 462 1942
rect 577 1942 1086 1947
rect 1097 1942 1142 1947
rect 1185 1942 1238 1947
rect 1313 1942 1358 1947
rect 1649 1942 1710 1947
rect 1737 1942 1766 1947
rect 1881 1942 1910 1947
rect 1969 1942 2022 1947
rect 2033 1942 2062 1947
rect 2073 1942 2174 1947
rect 2273 1942 2414 1947
rect 2433 1942 2470 1947
rect 2481 1942 2654 1947
rect 2993 1942 3038 1947
rect 3201 1942 3230 1947
rect 3329 1942 3406 1947
rect 577 1937 582 1942
rect 1377 1937 1454 1942
rect 2033 1937 2038 1942
rect 2433 1937 2438 1942
rect 3329 1937 3334 1942
rect 97 1927 102 1937
rect 233 1932 318 1937
rect 329 1932 366 1937
rect 457 1932 582 1937
rect 609 1932 1382 1937
rect 1449 1932 1510 1937
rect 1529 1932 1998 1937
rect 2017 1932 2038 1937
rect 2121 1932 2438 1937
rect 2465 1932 2494 1937
rect 2745 1932 2822 1937
rect 3281 1932 3334 1937
rect 3401 1937 3406 1942
rect 3401 1932 3430 1937
rect 1505 1927 1510 1932
rect 2745 1927 2750 1932
rect 65 1922 102 1927
rect 145 1922 214 1927
rect 225 1922 438 1927
rect 601 1922 630 1927
rect 713 1922 742 1927
rect 809 1922 910 1927
rect 1065 1922 1222 1927
rect 1233 1922 1438 1927
rect 1505 1922 1630 1927
rect 1721 1922 2062 1927
rect 2081 1922 2198 1927
rect 2233 1922 2302 1927
rect 2585 1922 2614 1927
rect 2713 1922 2750 1927
rect 2817 1927 2822 1932
rect 2817 1922 2846 1927
rect 65 1907 70 1922
rect 625 1917 718 1922
rect 945 1917 1046 1922
rect 2369 1917 2502 1922
rect 81 1912 110 1917
rect 177 1912 270 1917
rect 321 1912 350 1917
rect 449 1912 590 1917
rect 817 1912 950 1917
rect 1041 1912 1278 1917
rect 1345 1912 1374 1917
rect 1425 1912 1470 1917
rect 1545 1912 2374 1917
rect 2497 1912 2550 1917
rect 2761 1912 2814 1917
rect 2865 1912 3174 1917
rect 3289 1912 3430 1917
rect 345 1907 454 1912
rect 2569 1907 2670 1912
rect 65 1902 86 1907
rect 233 1902 294 1907
rect 537 1902 654 1907
rect 753 1902 854 1907
rect 961 1902 1126 1907
rect 1145 1902 1262 1907
rect 1281 1902 1318 1907
rect 1497 1902 1670 1907
rect 1729 1902 1790 1907
rect 1889 1902 1950 1907
rect 2001 1902 2102 1907
rect 2161 1902 2190 1907
rect 2217 1902 2262 1907
rect 2385 1902 2414 1907
rect 2449 1902 2478 1907
rect 2537 1902 2574 1907
rect 2665 1902 2694 1907
rect 2793 1902 2902 1907
rect 3393 1902 3438 1907
rect 873 1897 966 1902
rect 2001 1897 2006 1902
rect 297 1892 830 1897
rect 841 1892 878 1897
rect 985 1892 1174 1897
rect 1281 1892 1446 1897
rect 1505 1892 1598 1897
rect 1857 1892 2006 1897
rect 2041 1892 2406 1897
rect 2497 1892 2854 1897
rect 1169 1887 1262 1892
rect 2401 1887 2406 1892
rect 2897 1887 2982 1892
rect 793 1882 1046 1887
rect 1073 1882 1158 1887
rect 1257 1882 1358 1887
rect 1385 1882 1478 1887
rect 1529 1882 1558 1887
rect 1633 1882 1702 1887
rect 1745 1882 1942 1887
rect 1985 1882 2126 1887
rect 2145 1882 2166 1887
rect 2177 1882 2278 1887
rect 2305 1882 2366 1887
rect 2401 1882 2726 1887
rect 2769 1882 2822 1887
rect 2873 1882 2902 1887
rect 2977 1882 3046 1887
rect 529 1877 734 1882
rect 225 1872 286 1877
rect 281 1867 286 1872
rect 401 1872 534 1877
rect 729 1872 1686 1877
rect 1705 1872 1742 1877
rect 401 1867 406 1872
rect 1681 1867 1686 1872
rect 1737 1867 1742 1872
rect 1889 1872 2790 1877
rect 2937 1872 2966 1877
rect 1889 1867 1894 1872
rect 2785 1867 2942 1872
rect 281 1862 406 1867
rect 545 1862 718 1867
rect 801 1862 910 1867
rect 921 1862 1142 1867
rect 1153 1862 1486 1867
rect 1601 1862 1630 1867
rect 1681 1862 1718 1867
rect 1737 1862 1894 1867
rect 1977 1862 2046 1867
rect 2065 1862 2198 1867
rect 2209 1862 2326 1867
rect 2337 1862 2430 1867
rect 2569 1862 2598 1867
rect 2977 1862 3014 1867
rect 1481 1857 1606 1862
rect 593 1852 894 1857
rect 913 1852 990 1857
rect 1017 1852 1054 1857
rect 1065 1852 1118 1857
rect 1193 1852 1390 1857
rect 1441 1852 1462 1857
rect 425 1842 494 1847
rect 521 1842 926 1847
rect 1025 1842 1558 1847
rect 193 1832 1310 1837
rect 1337 1832 1486 1837
rect 1617 1832 1638 1837
rect 1649 1832 1670 1837
rect 441 1822 670 1827
rect 745 1822 990 1827
rect 1009 1822 1102 1827
rect 1217 1822 1254 1827
rect 1329 1822 1422 1827
rect 1449 1822 1494 1827
rect 1009 1817 1014 1822
rect 1489 1817 1494 1822
rect 337 1812 422 1817
rect 601 1812 646 1817
rect 697 1812 774 1817
rect 849 1812 918 1817
rect 929 1812 1014 1817
rect 1041 1812 1494 1817
rect 1601 1812 1622 1817
rect 337 1807 342 1812
rect 417 1807 582 1812
rect 1633 1807 1638 1832
rect 1681 1827 1686 1862
rect 2209 1857 2214 1862
rect 2593 1857 2766 1862
rect 2977 1857 2982 1862
rect 1913 1852 2214 1857
rect 2225 1852 2334 1857
rect 2761 1852 2982 1857
rect 1729 1842 1774 1847
rect 1809 1842 2398 1847
rect 2449 1842 2550 1847
rect 2593 1842 2742 1847
rect 3033 1842 3134 1847
rect 2449 1837 2454 1842
rect 1697 1832 2454 1837
rect 2545 1837 2550 1842
rect 3033 1837 3038 1842
rect 2545 1832 2686 1837
rect 2753 1832 3038 1837
rect 3129 1837 3134 1842
rect 3129 1832 3158 1837
rect 2681 1827 2758 1832
rect 1649 1822 1686 1827
rect 1769 1822 1862 1827
rect 1881 1822 1958 1827
rect 1977 1822 2070 1827
rect 2169 1822 2246 1827
rect 2281 1822 2334 1827
rect 2409 1822 2550 1827
rect 2065 1817 2174 1822
rect 1841 1812 1910 1817
rect 1961 1812 2046 1817
rect 2193 1812 2478 1817
rect 1657 1807 1822 1812
rect 2577 1807 2582 1827
rect 2625 1822 2662 1827
rect 3137 1822 3230 1827
rect 3241 1822 3318 1827
rect 2801 1817 2878 1822
rect 2729 1812 2806 1817
rect 2873 1812 2902 1817
rect 3009 1812 3086 1817
rect 3177 1812 3286 1817
rect 225 1802 342 1807
rect 577 1802 1374 1807
rect 1433 1802 1478 1807
rect 1545 1802 1662 1807
rect 1817 1802 1990 1807
rect 2049 1802 2110 1807
rect 2129 1802 2182 1807
rect 2201 1802 2342 1807
rect 2385 1802 2430 1807
rect 2457 1802 2582 1807
rect 2593 1802 2734 1807
rect 2817 1802 2870 1807
rect 2905 1802 2934 1807
rect 2945 1802 2974 1807
rect 3049 1802 3158 1807
rect 225 1797 230 1802
rect 2593 1797 2598 1802
rect 2729 1797 2822 1802
rect 201 1792 230 1797
rect 337 1792 742 1797
rect 809 1792 926 1797
rect 977 1792 1046 1797
rect 1057 1792 1198 1797
rect 1209 1792 1358 1797
rect 1385 1792 1454 1797
rect 1465 1792 2598 1797
rect 2841 1792 3070 1797
rect 3129 1792 3198 1797
rect 1057 1787 1062 1792
rect 2617 1787 2710 1792
rect 225 1782 310 1787
rect 401 1782 430 1787
rect 465 1782 502 1787
rect 601 1782 1062 1787
rect 1081 1782 1230 1787
rect 1273 1782 1374 1787
rect 1457 1782 1550 1787
rect 1577 1782 1998 1787
rect 2033 1782 2622 1787
rect 2705 1782 2774 1787
rect 2833 1782 2910 1787
rect 2945 1782 3102 1787
rect 305 1777 406 1782
rect 137 1772 206 1777
rect 609 1772 854 1777
rect 865 1772 966 1777
rect 985 1772 1038 1777
rect 1049 1772 1214 1777
rect 1305 1772 1502 1777
rect 1601 1772 1734 1777
rect 1777 1772 1958 1777
rect 2001 1772 2022 1777
rect 2033 1772 2486 1777
rect 2545 1772 2646 1777
rect 2657 1772 2694 1777
rect 2857 1772 3094 1777
rect 609 1767 614 1772
rect 1497 1767 1606 1772
rect 2001 1767 2006 1772
rect 137 1762 198 1767
rect 377 1762 462 1767
rect 481 1762 534 1767
rect 545 1762 614 1767
rect 625 1762 798 1767
rect 953 1762 1038 1767
rect 1057 1762 1270 1767
rect 1313 1762 1478 1767
rect 1625 1762 1790 1767
rect 1905 1762 2006 1767
rect 2017 1762 2174 1767
rect 2217 1762 2294 1767
rect 2337 1762 2406 1767
rect 2449 1762 2686 1767
rect 2849 1762 3102 1767
rect 433 1757 438 1762
rect 817 1757 910 1762
rect 2849 1757 2854 1762
rect 273 1752 326 1757
rect 433 1752 486 1757
rect 553 1752 630 1757
rect 641 1752 822 1757
rect 905 1752 1302 1757
rect 1417 1752 1606 1757
rect 1649 1752 1918 1757
rect 1977 1752 2030 1757
rect 2241 1752 2854 1757
rect 2865 1752 2958 1757
rect 3009 1752 3038 1757
rect 129 1742 214 1747
rect 129 1737 134 1742
rect 105 1732 134 1737
rect 209 1737 214 1742
rect 321 1737 326 1752
rect 641 1747 646 1752
rect 1297 1747 1422 1752
rect 345 1742 646 1747
rect 665 1742 774 1747
rect 833 1742 886 1747
rect 913 1742 1158 1747
rect 1185 1742 1278 1747
rect 1593 1742 1702 1747
rect 1713 1742 1878 1747
rect 1889 1742 2038 1747
rect 2129 1742 2230 1747
rect 2305 1742 2398 1747
rect 2465 1742 2526 1747
rect 2537 1742 2830 1747
rect 2841 1742 3190 1747
rect 3201 1742 3270 1747
rect 1441 1737 1550 1742
rect 209 1732 310 1737
rect 321 1732 638 1737
rect 753 1732 926 1737
rect 937 1732 1086 1737
rect 1201 1732 1342 1737
rect 1417 1732 1446 1737
rect 1545 1732 1630 1737
rect 1649 1732 1726 1737
rect 1753 1732 1838 1737
rect 1857 1732 1918 1737
rect 1993 1732 3070 1737
rect 305 1727 310 1732
rect 1649 1727 1654 1732
rect 1857 1727 1862 1732
rect 113 1722 198 1727
rect 305 1722 414 1727
rect 505 1722 558 1727
rect 593 1722 630 1727
rect 649 1722 758 1727
rect 817 1722 1102 1727
rect 1145 1722 1214 1727
rect 1265 1722 1358 1727
rect 1441 1722 1534 1727
rect 1609 1722 1654 1727
rect 1729 1722 1862 1727
rect 1873 1722 1902 1727
rect 1913 1722 3014 1727
rect 81 1712 166 1717
rect 177 1712 518 1717
rect 177 1707 182 1712
rect 161 1702 182 1707
rect 545 1702 614 1707
rect 625 1702 630 1722
rect 3009 1717 3014 1722
rect 3105 1722 3238 1727
rect 3105 1717 3110 1722
rect 721 1712 1262 1717
rect 1401 1712 1534 1717
rect 1545 1712 1662 1717
rect 1681 1712 1782 1717
rect 1881 1712 2158 1717
rect 2193 1712 2254 1717
rect 2281 1712 2326 1717
rect 2337 1712 2366 1717
rect 2401 1712 2430 1717
rect 2473 1712 2518 1717
rect 2633 1712 2798 1717
rect 2809 1712 2886 1717
rect 2953 1712 2974 1717
rect 3009 1712 3110 1717
rect 3321 1712 3374 1717
rect 2321 1707 2326 1712
rect 641 1702 870 1707
rect 889 1702 1014 1707
rect 1033 1702 1222 1707
rect 1257 1702 1350 1707
rect 1497 1702 1574 1707
rect 1721 1702 2230 1707
rect 2241 1702 2278 1707
rect 2321 1702 2446 1707
rect 2577 1702 2606 1707
rect 2657 1702 2718 1707
rect 2769 1702 2990 1707
rect 3129 1702 3174 1707
rect 281 1697 526 1702
rect 609 1697 614 1702
rect 865 1697 870 1702
rect 1009 1697 1014 1702
rect 177 1692 286 1697
rect 521 1692 574 1697
rect 609 1692 678 1697
rect 865 1692 990 1697
rect 1009 1692 1310 1697
rect 1329 1692 1414 1697
rect 1433 1692 1654 1697
rect 1761 1692 1806 1697
rect 1849 1692 1902 1697
rect 1929 1692 2454 1697
rect 2513 1692 2534 1697
rect 2553 1692 2574 1697
rect 2617 1692 2678 1697
rect 2825 1692 2854 1697
rect 2529 1687 2534 1692
rect 2673 1687 2830 1692
rect 281 1682 726 1687
rect 745 1682 1302 1687
rect 1465 1682 1494 1687
rect 1601 1682 1910 1687
rect 1937 1682 2070 1687
rect 2145 1682 2262 1687
rect 2297 1682 2374 1687
rect 2433 1682 2510 1687
rect 2529 1682 2574 1687
rect 2625 1682 2654 1687
rect 3121 1682 3182 1687
rect 2369 1677 2374 1682
rect 345 1672 374 1677
rect 473 1672 950 1677
rect 1065 1672 2358 1677
rect 2369 1672 2798 1677
rect 2929 1672 2958 1677
rect 369 1667 478 1672
rect 961 1667 1070 1672
rect 2353 1667 2358 1672
rect 497 1662 614 1667
rect 705 1662 798 1667
rect 929 1662 966 1667
rect 1113 1662 1174 1667
rect 1185 1662 1358 1667
rect 1465 1662 1638 1667
rect 1657 1662 1702 1667
rect 1825 1662 1846 1667
rect 1897 1662 2102 1667
rect 2113 1662 2334 1667
rect 2353 1662 2558 1667
rect 2633 1662 2822 1667
rect 3089 1662 3158 1667
rect 3273 1662 3382 1667
rect 817 1657 910 1662
rect 177 1652 302 1657
rect 329 1652 422 1657
rect 449 1652 582 1657
rect 593 1652 822 1657
rect 905 1652 998 1657
rect 1113 1652 1302 1657
rect 1433 1652 1462 1657
rect 1513 1652 1710 1657
rect 1753 1652 2134 1657
rect 2161 1652 2262 1657
rect 2281 1652 2566 1657
rect 2657 1652 2766 1657
rect 3049 1652 3070 1657
rect 3225 1652 3270 1657
rect 577 1647 582 1652
rect 2257 1647 2262 1652
rect 65 1642 94 1647
rect 193 1642 342 1647
rect 385 1642 566 1647
rect 577 1642 662 1647
rect 681 1642 926 1647
rect 969 1642 1286 1647
rect 1321 1642 1414 1647
rect 1457 1642 1486 1647
rect 65 1607 70 1642
rect 1321 1637 1326 1642
rect 89 1632 302 1637
rect 313 1632 382 1637
rect 513 1632 630 1637
rect 641 1632 1326 1637
rect 1409 1637 1414 1642
rect 1513 1637 1518 1647
rect 1617 1642 1654 1647
rect 1729 1642 1782 1647
rect 1817 1642 1918 1647
rect 1953 1642 2222 1647
rect 2257 1642 2334 1647
rect 2409 1642 2654 1647
rect 2841 1642 2878 1647
rect 2921 1642 2990 1647
rect 3041 1642 3094 1647
rect 3225 1642 3286 1647
rect 1409 1632 1518 1637
rect 1577 1632 1694 1637
rect 1873 1632 1910 1637
rect 1937 1632 2086 1637
rect 2185 1632 2486 1637
rect 2649 1632 2862 1637
rect 401 1627 494 1632
rect 2481 1627 2654 1632
rect 2857 1627 2862 1632
rect 2921 1632 3022 1637
rect 3121 1632 3350 1637
rect 2921 1627 2926 1632
rect 113 1622 182 1627
rect 305 1622 406 1627
rect 489 1622 526 1627
rect 665 1622 702 1627
rect 769 1622 838 1627
rect 921 1622 1126 1627
rect 1185 1622 1214 1627
rect 1249 1622 1350 1627
rect 1385 1622 1934 1627
rect 2017 1622 2046 1627
rect 2121 1622 2214 1627
rect 2241 1622 2462 1627
rect 2673 1622 2718 1627
rect 2857 1622 2926 1627
rect 3001 1622 3110 1627
rect 3257 1622 3286 1627
rect 113 1612 150 1617
rect 65 1602 110 1607
rect 177 1597 182 1622
rect 569 1617 646 1622
rect 329 1612 574 1617
rect 641 1612 974 1617
rect 1001 1612 1054 1617
rect 1121 1607 1126 1622
rect 1193 1612 1214 1617
rect 1409 1612 1662 1617
rect 1913 1612 2110 1617
rect 2185 1612 2518 1617
rect 2625 1612 2694 1617
rect 1409 1607 1414 1612
rect 1657 1607 1918 1612
rect 2105 1607 2190 1612
rect 209 1602 326 1607
rect 433 1602 462 1607
rect 585 1602 870 1607
rect 1025 1602 1110 1607
rect 1121 1602 1302 1607
rect 1329 1602 1414 1607
rect 1425 1602 1582 1607
rect 1609 1602 1638 1607
rect 1937 1602 1966 1607
rect 2209 1602 2254 1607
rect 2361 1602 2414 1607
rect 2481 1597 2582 1602
rect 2833 1597 2838 1617
rect 3281 1612 3286 1622
rect 3329 1622 3374 1627
rect 3329 1607 3334 1622
rect 3057 1602 3102 1607
rect 3305 1602 3334 1607
rect 113 1592 142 1597
rect 177 1592 302 1597
rect 321 1592 406 1597
rect 417 1592 446 1597
rect 537 1592 678 1597
rect 921 1592 1374 1597
rect 1457 1592 1558 1597
rect 1657 1592 1718 1597
rect 1785 1592 1854 1597
rect 1929 1592 2038 1597
rect 2057 1592 2190 1597
rect 2297 1592 2382 1597
rect 2457 1592 2486 1597
rect 2577 1592 2606 1597
rect 2697 1592 2838 1597
rect 2849 1592 2934 1597
rect 3257 1592 3334 1597
rect 697 1587 902 1592
rect 1369 1587 1462 1592
rect 2057 1587 2062 1592
rect 225 1582 254 1587
rect 385 1582 702 1587
rect 897 1582 1094 1587
rect 1145 1582 1270 1587
rect 1305 1582 1350 1587
rect 1481 1582 1574 1587
rect 1777 1582 1830 1587
rect 1881 1582 2062 1587
rect 2185 1587 2190 1592
rect 2849 1587 2854 1592
rect 2185 1582 2230 1587
rect 2241 1582 2270 1587
rect 2393 1582 2702 1587
rect 225 1572 230 1582
rect 2265 1577 2398 1582
rect 2697 1577 2702 1582
rect 2793 1582 2854 1587
rect 2881 1582 3070 1587
rect 3209 1582 3254 1587
rect 2793 1577 2798 1582
rect 273 1572 358 1577
rect 385 1572 406 1577
rect 425 1572 774 1577
rect 785 1572 1158 1577
rect 1233 1572 1294 1577
rect 1313 1572 1478 1577
rect 1537 1572 1638 1577
rect 1697 1572 1910 1577
rect 1921 1572 1958 1577
rect 2049 1572 2190 1577
rect 2417 1572 2454 1577
rect 2505 1572 2678 1577
rect 2697 1572 2798 1577
rect 2873 1572 3150 1577
rect 3177 1572 3254 1577
rect 273 1567 278 1572
rect 89 1562 278 1567
rect 353 1567 358 1572
rect 401 1567 406 1572
rect 1153 1567 1158 1572
rect 2417 1567 2422 1572
rect 3249 1567 3254 1572
rect 3313 1572 3350 1577
rect 3313 1567 3318 1572
rect 353 1562 382 1567
rect 401 1562 422 1567
rect 457 1562 502 1567
rect 545 1562 574 1567
rect 625 1562 662 1567
rect 809 1562 918 1567
rect 1001 1562 1134 1567
rect 1153 1562 1198 1567
rect 1241 1562 1286 1567
rect 1297 1562 1334 1567
rect 1369 1562 1630 1567
rect 1657 1562 1990 1567
rect 2001 1562 2046 1567
rect 2281 1562 2422 1567
rect 2441 1562 2670 1567
rect 2817 1562 2966 1567
rect 3001 1562 3142 1567
rect 3249 1562 3318 1567
rect 681 1557 790 1562
rect 1297 1557 1302 1562
rect 2817 1557 2822 1562
rect 2961 1557 2966 1562
rect 129 1547 134 1557
rect 249 1552 686 1557
rect 785 1552 814 1557
rect 977 1552 1022 1557
rect 1065 1552 1214 1557
rect 1257 1552 1302 1557
rect 1337 1552 1430 1557
rect 1449 1552 2150 1557
rect 2161 1552 2278 1557
rect 2337 1552 2414 1557
rect 2529 1552 2822 1557
rect 2841 1552 2910 1557
rect 2961 1552 3118 1557
rect 2433 1547 2534 1552
rect 89 1542 390 1547
rect 409 1542 462 1547
rect 521 1542 582 1547
rect 593 1542 614 1547
rect 633 1542 886 1547
rect 921 1542 1190 1547
rect 1201 1542 1254 1547
rect 1265 1542 1318 1547
rect 1337 1542 1382 1547
rect 1489 1542 1598 1547
rect 1817 1542 2022 1547
rect 2033 1542 2118 1547
rect 2257 1542 2374 1547
rect 385 1537 390 1542
rect 609 1537 614 1542
rect 881 1537 886 1542
rect 1249 1537 1254 1542
rect 1409 1537 1494 1542
rect 1617 1537 1742 1542
rect 2033 1537 2038 1542
rect 2433 1537 2438 1547
rect 2553 1542 2590 1547
rect 2601 1542 2718 1547
rect 3337 1542 3430 1547
rect 97 1532 150 1537
rect 233 1532 254 1537
rect 265 1532 334 1537
rect 385 1532 598 1537
rect 609 1532 694 1537
rect 705 1532 822 1537
rect 841 1532 870 1537
rect 881 1532 1086 1537
rect 1249 1532 1278 1537
rect 1289 1532 1358 1537
rect 1385 1532 1414 1537
rect 1505 1532 1622 1537
rect 1737 1532 2038 1537
rect 2089 1532 2238 1537
rect 2281 1532 2438 1537
rect 2481 1532 2558 1537
rect 2833 1532 2934 1537
rect 2969 1532 3070 1537
rect 3193 1532 3278 1537
rect 3393 1532 3438 1537
rect 249 1527 254 1532
rect 817 1527 822 1532
rect 1105 1527 1230 1532
rect 2481 1527 2486 1532
rect 2969 1527 2974 1532
rect 65 1522 142 1527
rect 153 1522 182 1527
rect 201 1522 246 1527
rect 249 1522 286 1527
rect 417 1522 438 1527
rect 449 1522 542 1527
rect 737 1522 790 1527
rect 817 1522 998 1527
rect 1041 1522 1110 1527
rect 1225 1522 1726 1527
rect 1905 1522 2022 1527
rect 2121 1522 2486 1527
rect 2513 1522 2734 1527
rect 2841 1522 2974 1527
rect 3065 1527 3070 1532
rect 3065 1522 3206 1527
rect 3241 1522 3342 1527
rect 177 1507 182 1522
rect 241 1517 246 1522
rect 649 1517 718 1522
rect 1721 1517 1910 1522
rect 2017 1517 2126 1522
rect 241 1512 654 1517
rect 713 1512 1430 1517
rect 1665 1512 1702 1517
rect 1929 1512 1998 1517
rect 2145 1512 2574 1517
rect 2585 1512 2606 1517
rect 2913 1512 3054 1517
rect 3177 1512 3406 1517
rect 1425 1507 1670 1512
rect 105 1502 182 1507
rect 225 1502 278 1507
rect 401 1502 486 1507
rect 505 1502 590 1507
rect 665 1502 710 1507
rect 769 1502 1406 1507
rect 1689 1502 1798 1507
rect 1913 1502 2022 1507
rect 2177 1502 2214 1507
rect 2401 1502 2478 1507
rect 2641 1502 2750 1507
rect 3169 1502 3222 1507
rect 2041 1497 2158 1502
rect 2233 1497 2302 1502
rect 2641 1497 2646 1502
rect 185 1492 270 1497
rect 497 1492 990 1497
rect 1073 1492 1174 1497
rect 1201 1492 1414 1497
rect 1481 1492 1574 1497
rect 1649 1492 2046 1497
rect 2153 1492 2238 1497
rect 2297 1492 2646 1497
rect 2745 1497 2750 1502
rect 2961 1497 3054 1502
rect 2745 1492 2966 1497
rect 3049 1492 3214 1497
rect 3297 1492 3374 1497
rect 289 1487 422 1492
rect 265 1482 294 1487
rect 417 1482 838 1487
rect 857 1482 1494 1487
rect 1513 1482 1710 1487
rect 1769 1482 1958 1487
rect 1993 1482 2286 1487
rect 2457 1482 2478 1487
rect 2657 1482 2734 1487
rect 2977 1482 3046 1487
rect 313 1472 406 1477
rect 513 1472 542 1477
rect 641 1472 686 1477
rect 729 1472 870 1477
rect 881 1472 1078 1477
rect 1097 1472 1238 1477
rect 1265 1472 1318 1477
rect 1329 1472 1374 1477
rect 1601 1472 1838 1477
rect 2001 1472 2046 1477
rect 2073 1472 2222 1477
rect 2241 1472 2774 1477
rect 433 1467 518 1472
rect 1393 1467 1494 1472
rect 1857 1467 1950 1472
rect 2241 1467 2246 1472
rect 81 1462 238 1467
rect 273 1462 310 1467
rect 337 1462 438 1467
rect 537 1462 598 1467
rect 793 1462 822 1467
rect 305 1457 310 1462
rect 617 1457 710 1462
rect 817 1457 822 1462
rect 881 1462 1398 1467
rect 1489 1462 1590 1467
rect 1705 1462 1862 1467
rect 1945 1462 2246 1467
rect 2425 1462 2526 1467
rect 2633 1462 2710 1467
rect 2793 1462 2870 1467
rect 881 1457 886 1462
rect 1585 1457 1710 1462
rect 2521 1457 2638 1462
rect 2793 1457 2798 1462
rect 137 1452 158 1457
rect 193 1452 238 1457
rect 257 1452 294 1457
rect 305 1452 342 1457
rect 449 1452 622 1457
rect 705 1452 734 1457
rect 817 1452 886 1457
rect 929 1452 990 1457
rect 1025 1452 1270 1457
rect 1305 1452 1374 1457
rect 1385 1452 1486 1457
rect 1729 1452 1934 1457
rect 2025 1452 2078 1457
rect 2137 1452 2230 1457
rect 2265 1452 2406 1457
rect 2657 1452 2798 1457
rect 2865 1457 2870 1462
rect 2865 1452 2894 1457
rect 3409 1452 3438 1457
rect 2265 1447 2270 1452
rect 65 1442 174 1447
rect 193 1442 750 1447
rect 945 1442 1462 1447
rect 1561 1442 1606 1447
rect 1745 1442 1830 1447
rect 1889 1442 1974 1447
rect 2041 1442 2166 1447
rect 2177 1442 2270 1447
rect 2401 1447 2406 1452
rect 2401 1442 2446 1447
rect 2505 1442 2638 1447
rect 2737 1442 2766 1447
rect 2833 1442 2998 1447
rect 3065 1442 3110 1447
rect 3321 1442 3414 1447
rect 193 1437 198 1442
rect 1889 1437 1894 1442
rect 2289 1437 2382 1442
rect 2505 1437 2510 1442
rect 153 1432 198 1437
rect 241 1432 422 1437
rect 545 1432 582 1437
rect 737 1432 774 1437
rect 905 1432 1014 1437
rect 1049 1432 1094 1437
rect 1105 1432 1214 1437
rect 1313 1432 1382 1437
rect 1553 1432 1694 1437
rect 1777 1432 1894 1437
rect 1913 1432 2030 1437
rect 2137 1432 2294 1437
rect 2377 1432 2510 1437
rect 2633 1437 2638 1442
rect 2633 1432 2910 1437
rect 2025 1427 2142 1432
rect 81 1422 110 1427
rect 217 1422 358 1427
rect 433 1422 526 1427
rect 577 1422 790 1427
rect 809 1422 942 1427
rect 993 1422 1030 1427
rect 1081 1422 1110 1427
rect 1137 1422 1182 1427
rect 1281 1422 1302 1427
rect 1425 1422 1462 1427
rect 1537 1422 1566 1427
rect 1681 1422 1798 1427
rect 2161 1422 2262 1427
rect 2281 1422 2302 1427
rect 2321 1422 2382 1427
rect 2521 1422 2814 1427
rect 2849 1422 2910 1427
rect 3089 1422 3110 1427
rect 3289 1422 3374 1427
rect 81 1407 86 1422
rect 785 1417 790 1422
rect 2257 1417 2262 1422
rect 2321 1417 2326 1422
rect 97 1412 206 1417
rect 249 1412 278 1417
rect 385 1412 566 1417
rect 689 1412 750 1417
rect 785 1412 854 1417
rect 985 1412 1102 1417
rect 1129 1412 1302 1417
rect 1345 1412 1446 1417
rect 1457 1412 2078 1417
rect 2129 1407 2134 1417
rect 2257 1412 2326 1417
rect 2393 1412 2574 1417
rect 2777 1412 2894 1417
rect 2937 1412 3062 1417
rect 3113 1412 3246 1417
rect 2593 1407 2758 1412
rect 2937 1407 2942 1412
rect 81 1402 126 1407
rect 193 1402 318 1407
rect 377 1402 638 1407
rect 705 1402 862 1407
rect 921 1402 966 1407
rect 977 1402 1054 1407
rect 1153 1402 1582 1407
rect 1673 1402 1742 1407
rect 1777 1402 1830 1407
rect 2089 1402 2134 1407
rect 2161 1402 2598 1407
rect 2753 1402 2942 1407
rect 3057 1407 3062 1412
rect 3057 1402 3086 1407
rect 3177 1402 3278 1407
rect 3369 1402 3398 1407
rect 977 1397 982 1402
rect 1577 1397 1678 1402
rect 1777 1397 1782 1402
rect 1849 1397 2022 1402
rect 2161 1397 2166 1402
rect 97 1392 174 1397
rect 273 1392 710 1397
rect 865 1392 982 1397
rect 993 1392 1206 1397
rect 1233 1392 1558 1397
rect 1697 1392 1782 1397
rect 1801 1392 1854 1397
rect 2017 1392 2046 1397
rect 2105 1392 2166 1397
rect 2185 1392 2286 1397
rect 2297 1392 2334 1397
rect 2377 1392 2542 1397
rect 2569 1392 3070 1397
rect 3361 1392 3414 1397
rect 81 1382 102 1387
rect 273 1382 278 1392
rect 361 1382 454 1387
rect 497 1382 670 1387
rect 961 1382 990 1387
rect 1073 1382 1174 1387
rect 1217 1382 1270 1387
rect 1313 1382 1366 1387
rect 1377 1382 1470 1387
rect 1553 1382 1606 1387
rect 1665 1382 2654 1387
rect 2745 1382 2878 1387
rect 3233 1382 3286 1387
rect 1361 1377 1366 1382
rect 345 1372 430 1377
rect 641 1372 742 1377
rect 881 1372 1110 1377
rect 1121 1372 1238 1377
rect 1257 1372 1350 1377
rect 1361 1372 1414 1377
rect 1513 1372 1566 1377
rect 1585 1372 1734 1377
rect 1769 1372 1878 1377
rect 2049 1372 2246 1377
rect 2465 1372 2502 1377
rect 2521 1372 2566 1377
rect 2577 1372 2622 1377
rect 2809 1372 2870 1377
rect 2993 1372 3022 1377
rect 1105 1367 1110 1372
rect 1233 1367 1238 1372
rect 1897 1367 2030 1372
rect 2265 1367 2446 1372
rect 321 1362 350 1367
rect 441 1362 846 1367
rect 1105 1362 1214 1367
rect 1233 1362 1262 1367
rect 1273 1362 1574 1367
rect 1625 1362 1902 1367
rect 2025 1362 2270 1367
rect 2441 1362 2622 1367
rect 2833 1362 3070 1367
rect 345 1357 446 1362
rect 2833 1357 2838 1362
rect 465 1352 502 1357
rect 665 1352 694 1357
rect 977 1352 1430 1357
rect 1681 1352 2630 1357
rect 2705 1352 2838 1357
rect 2841 1352 2878 1357
rect 2953 1352 2998 1357
rect 713 1347 886 1352
rect 1465 1347 1582 1352
rect 2841 1347 2846 1352
rect 81 1342 158 1347
rect 353 1342 390 1347
rect 529 1342 598 1347
rect 649 1342 718 1347
rect 881 1342 1006 1347
rect 1089 1342 1118 1347
rect 1137 1342 1286 1347
rect 1313 1342 1430 1347
rect 1441 1342 1470 1347
rect 1577 1342 1606 1347
rect 1697 1342 2846 1347
rect 2857 1342 2910 1347
rect 2961 1342 3110 1347
rect 3361 1342 3406 1347
rect 1313 1337 1318 1342
rect 1425 1337 1430 1342
rect 257 1332 294 1337
rect 385 1332 422 1337
rect 537 1332 614 1337
rect 673 1332 942 1337
rect 953 1332 1110 1337
rect 1265 1332 1318 1337
rect 1329 1332 1406 1337
rect 1425 1332 1478 1337
rect 1537 1332 1790 1337
rect 1857 1332 1974 1337
rect 2017 1332 2102 1337
rect 2113 1332 2534 1337
rect 2633 1332 2782 1337
rect 2945 1332 2998 1337
rect 3233 1332 3302 1337
rect 209 1322 598 1327
rect 721 1322 918 1327
rect 1185 1322 1870 1327
rect 1969 1322 2038 1327
rect 2113 1322 2118 1332
rect 2137 1322 2198 1327
rect 2209 1322 2230 1327
rect 2241 1322 2246 1332
rect 2801 1327 2918 1332
rect 2297 1322 2462 1327
rect 2585 1322 2806 1327
rect 2913 1322 3110 1327
rect 3201 1322 3278 1327
rect 97 1312 158 1317
rect 281 1312 318 1317
rect 353 1312 398 1317
rect 481 1312 686 1317
rect 761 1312 870 1317
rect 913 1312 918 1322
rect 1065 1312 1238 1317
rect 1265 1312 1806 1317
rect 1833 1312 1918 1317
rect 1953 1312 2118 1317
rect 2153 1312 2350 1317
rect 2393 1312 2582 1317
rect 2633 1312 2694 1317
rect 2809 1312 2902 1317
rect 3025 1312 3054 1317
rect 2897 1307 3030 1312
rect 289 1302 470 1307
rect 465 1297 470 1302
rect 553 1302 582 1307
rect 793 1302 1062 1307
rect 1129 1302 1182 1307
rect 1201 1302 1478 1307
rect 1553 1302 1590 1307
rect 1601 1302 2062 1307
rect 2073 1302 2878 1307
rect 553 1297 558 1302
rect 249 1292 342 1297
rect 465 1292 558 1297
rect 617 1292 670 1297
rect 729 1292 758 1297
rect 953 1292 974 1297
rect 1225 1292 1662 1297
rect 1777 1292 2142 1297
rect 2201 1292 2422 1297
rect 2457 1292 2846 1297
rect 2881 1292 3054 1297
rect 801 1287 934 1292
rect 993 1287 1206 1292
rect 305 1282 430 1287
rect 593 1282 806 1287
rect 929 1282 998 1287
rect 1201 1282 1254 1287
rect 1297 1282 1446 1287
rect 1633 1282 1694 1287
rect 1785 1282 1838 1287
rect 1961 1282 2038 1287
rect 2049 1282 2078 1287
rect 2105 1282 2182 1287
rect 2217 1282 2286 1287
rect 2409 1282 2438 1287
rect 2673 1282 2702 1287
rect 2793 1282 2830 1287
rect 2937 1282 2958 1287
rect 297 1272 734 1277
rect 817 1272 886 1277
rect 905 1272 1014 1277
rect 1065 1272 1262 1277
rect 1009 1267 1014 1272
rect 1297 1267 1302 1282
rect 1465 1277 1590 1282
rect 2457 1277 2582 1282
rect 2697 1277 2798 1282
rect 329 1262 358 1267
rect 353 1257 358 1262
rect 441 1262 478 1267
rect 633 1262 750 1267
rect 865 1262 990 1267
rect 1009 1262 1302 1267
rect 1313 1272 1470 1277
rect 1585 1272 1638 1277
rect 1825 1272 2462 1277
rect 2577 1272 2606 1277
rect 2817 1272 2974 1277
rect 441 1257 446 1262
rect 545 1257 614 1262
rect 1313 1257 1318 1272
rect 1401 1262 1774 1267
rect 353 1252 446 1257
rect 465 1252 550 1257
rect 609 1252 1054 1257
rect 1169 1252 1318 1257
rect 1449 1252 1702 1257
rect 1825 1247 1830 1272
rect 1929 1262 2046 1267
rect 2081 1262 2422 1267
rect 2473 1262 2958 1267
rect 1841 1252 2510 1257
rect 2537 1252 2662 1257
rect 2753 1252 2814 1257
rect 2833 1247 2926 1252
rect 561 1242 694 1247
rect 881 1242 926 1247
rect 961 1242 1062 1247
rect 1089 1242 1142 1247
rect 1209 1242 1366 1247
rect 1585 1242 1622 1247
rect 1761 1242 1862 1247
rect 1873 1242 2190 1247
rect 2217 1242 2270 1247
rect 2313 1242 2366 1247
rect 2441 1242 2526 1247
rect 2753 1242 2774 1247
rect 2801 1242 2838 1247
rect 2921 1242 3038 1247
rect 3185 1242 3286 1247
rect 777 1232 1206 1237
rect 201 1222 342 1227
rect 377 1222 406 1227
rect 441 1222 518 1227
rect 649 1222 694 1227
rect 937 1222 1126 1227
rect 1185 1222 1294 1227
rect 1329 1217 1334 1242
rect 1641 1237 1742 1242
rect 2545 1237 2734 1242
rect 1385 1232 1646 1237
rect 1737 1232 2406 1237
rect 2505 1232 2550 1237
rect 2729 1232 2910 1237
rect 3017 1232 3094 1237
rect 3177 1232 3214 1237
rect 3297 1232 3358 1237
rect 3401 1232 3430 1237
rect 2401 1227 2486 1232
rect 1345 1222 1430 1227
rect 1569 1222 1654 1227
rect 1681 1222 1734 1227
rect 1873 1222 1934 1227
rect 2057 1222 2134 1227
rect 2145 1222 2174 1227
rect 2209 1222 2310 1227
rect 2337 1222 2390 1227
rect 2481 1222 2710 1227
rect 2745 1222 2798 1227
rect 3337 1222 3398 1227
rect 1473 1217 1550 1222
rect 209 1212 262 1217
rect 297 1212 326 1217
rect 577 1212 670 1217
rect 817 1207 822 1217
rect 985 1212 1070 1217
rect 1329 1212 1478 1217
rect 1545 1212 2166 1217
rect 2177 1212 2886 1217
rect 2913 1212 3094 1217
rect 3185 1212 3350 1217
rect 3385 1212 3414 1217
rect 857 1207 966 1212
rect 1089 1207 1206 1212
rect 2177 1207 2182 1212
rect 105 1202 422 1207
rect 457 1202 590 1207
rect 641 1202 822 1207
rect 833 1202 862 1207
rect 961 1202 1094 1207
rect 1201 1202 1398 1207
rect 1489 1202 2030 1207
rect 2129 1202 2182 1207
rect 2233 1202 2270 1207
rect 2337 1202 2446 1207
rect 2465 1202 2950 1207
rect 3137 1202 3262 1207
rect 1393 1197 1494 1202
rect 2465 1197 2470 1202
rect 313 1192 1142 1197
rect 1161 1192 1190 1197
rect 1289 1192 1374 1197
rect 1513 1192 2198 1197
rect 2281 1192 2470 1197
rect 2513 1192 2878 1197
rect 169 1187 270 1192
rect 2193 1187 2286 1192
rect 145 1182 174 1187
rect 265 1182 310 1187
rect 353 1182 470 1187
rect 505 1182 614 1187
rect 625 1182 902 1187
rect 929 1182 1062 1187
rect 1073 1182 1390 1187
rect 1489 1182 1878 1187
rect 1969 1182 2030 1187
rect 2049 1182 2174 1187
rect 2305 1182 2342 1187
rect 2353 1182 2550 1187
rect 2625 1182 2774 1187
rect 2817 1182 2974 1187
rect 3057 1182 3134 1187
rect 3321 1182 3374 1187
rect 1057 1177 1062 1182
rect 185 1172 238 1177
rect 385 1172 414 1177
rect 585 1172 886 1177
rect 945 1172 998 1177
rect 1009 1172 1038 1177
rect 1057 1172 1854 1177
rect 1953 1172 2302 1177
rect 2361 1172 2598 1177
rect 2649 1172 2686 1177
rect 2713 1172 3078 1177
rect 3185 1172 3262 1177
rect 257 1167 366 1172
rect 993 1167 998 1172
rect 233 1162 262 1167
rect 361 1162 574 1167
rect 673 1162 710 1167
rect 737 1162 934 1167
rect 945 1162 982 1167
rect 993 1162 1054 1167
rect 1073 1162 1126 1167
rect 1369 1162 2766 1167
rect 3017 1162 3198 1167
rect 569 1157 678 1162
rect 1073 1157 1078 1162
rect 1145 1157 1246 1162
rect 241 1152 454 1157
rect 697 1152 854 1157
rect 897 1152 1078 1157
rect 1113 1152 1150 1157
rect 1241 1152 1270 1157
rect 1377 1152 1494 1157
rect 1649 1152 1806 1157
rect 1889 1152 1974 1157
rect 1993 1152 2150 1157
rect 2185 1152 2238 1157
rect 2337 1152 2438 1157
rect 2569 1152 2918 1157
rect 3129 1152 3198 1157
rect 1289 1147 1382 1152
rect 1649 1147 1654 1152
rect 1889 1147 1894 1152
rect 2457 1147 2550 1152
rect 105 1142 134 1147
rect 145 1142 214 1147
rect 361 1142 422 1147
rect 457 1142 486 1147
rect 593 1142 678 1147
rect 753 1142 862 1147
rect 953 1142 1294 1147
rect 1393 1142 1654 1147
rect 1665 1142 1894 1147
rect 1913 1142 2134 1147
rect 2153 1142 2214 1147
rect 2241 1142 2302 1147
rect 2313 1142 2358 1147
rect 2393 1142 2462 1147
rect 2545 1142 2718 1147
rect 2873 1142 2902 1147
rect 3073 1142 3222 1147
rect 233 1137 342 1142
rect 1393 1137 1398 1142
rect 2713 1137 2878 1142
rect 193 1132 238 1137
rect 337 1132 774 1137
rect 833 1132 974 1137
rect 1089 1132 1398 1137
rect 1409 1132 1446 1137
rect 1601 1132 1686 1137
rect 193 1127 198 1132
rect 1393 1127 1398 1132
rect 1697 1127 1702 1137
rect 1937 1127 1942 1137
rect 2009 1132 2390 1137
rect 2409 1132 2574 1137
rect 2609 1132 2654 1137
rect 2689 1127 2694 1137
rect 3201 1132 3254 1137
rect 161 1122 198 1127
rect 217 1122 254 1127
rect 289 1122 350 1127
rect 377 1122 518 1127
rect 641 1122 710 1127
rect 857 1122 886 1127
rect 993 1122 1254 1127
rect 1345 1122 1382 1127
rect 1393 1122 1414 1127
rect 1465 1122 1558 1127
rect 1569 1122 1598 1127
rect 1665 1122 1702 1127
rect 1713 1122 1782 1127
rect 1801 1122 1918 1127
rect 1937 1122 2022 1127
rect 2065 1122 2502 1127
rect 2521 1122 2606 1127
rect 2665 1122 3062 1127
rect 1345 1117 1350 1122
rect 1801 1117 1806 1122
rect 385 1112 414 1117
rect 897 1112 1014 1117
rect 1081 1112 1110 1117
rect 1345 1112 1806 1117
rect 1913 1117 1918 1122
rect 3057 1117 3062 1122
rect 3153 1122 3238 1127
rect 3153 1117 3158 1122
rect 1913 1112 2886 1117
rect 3057 1112 3158 1117
rect 3177 1112 3230 1117
rect 777 1107 870 1112
rect 1129 1107 1286 1112
rect 3249 1107 3254 1132
rect 3273 1112 3318 1117
rect 81 1102 134 1107
rect 177 1102 222 1107
rect 297 1102 430 1107
rect 657 1102 782 1107
rect 865 1102 934 1107
rect 929 1097 934 1102
rect 1017 1102 1134 1107
rect 1281 1102 1534 1107
rect 1641 1102 1974 1107
rect 1993 1102 2134 1107
rect 2177 1102 2406 1107
rect 2417 1102 2494 1107
rect 2505 1102 2622 1107
rect 2745 1102 2790 1107
rect 3185 1102 3254 1107
rect 1017 1097 1022 1102
rect 1529 1097 1646 1102
rect 473 1092 494 1097
rect 593 1092 726 1097
rect 793 1092 854 1097
rect 929 1092 1022 1097
rect 1041 1092 1174 1097
rect 1201 1092 1270 1097
rect 1433 1092 1510 1097
rect 1665 1092 1686 1097
rect 1697 1092 1806 1097
rect 1889 1092 2686 1097
rect 2769 1092 2838 1097
rect 1505 1087 1510 1092
rect 1697 1087 1702 1092
rect 81 1082 166 1087
rect 321 1082 774 1087
rect 817 1082 910 1087
rect 1041 1082 1070 1087
rect 1425 1082 1494 1087
rect 1505 1082 1558 1087
rect 1569 1082 1598 1087
rect 1649 1082 1702 1087
rect 1761 1082 2478 1087
rect 2593 1082 2670 1087
rect 2721 1082 2798 1087
rect 129 1072 1198 1077
rect 1345 1072 1718 1077
rect 1921 1072 2070 1077
rect 2257 1072 2502 1077
rect 2513 1072 2598 1077
rect 2609 1072 2654 1077
rect 2673 1072 2854 1077
rect 1801 1067 1926 1072
rect 2065 1067 2182 1072
rect 337 1062 438 1067
rect 489 1062 918 1067
rect 993 1062 1062 1067
rect 1129 1062 1286 1067
rect 1401 1062 1806 1067
rect 1945 1062 2046 1067
rect 2177 1062 2734 1067
rect 993 1057 998 1062
rect 553 1052 654 1057
rect 689 1052 998 1057
rect 1017 1052 1686 1057
rect 1817 1052 1990 1057
rect 2009 1052 2150 1057
rect 2217 1052 2278 1057
rect 2313 1052 2462 1057
rect 2489 1052 2630 1057
rect 393 1047 534 1052
rect 1705 1047 1798 1052
rect 2649 1047 2750 1052
rect 369 1042 398 1047
rect 529 1042 702 1047
rect 785 1042 1550 1047
rect 1585 1042 1710 1047
rect 1793 1042 1830 1047
rect 1849 1042 2654 1047
rect 2745 1042 2774 1047
rect 697 1037 790 1042
rect 345 1032 406 1037
rect 433 1032 486 1037
rect 529 1032 582 1037
rect 633 1032 678 1037
rect 809 1032 998 1037
rect 1009 1032 1118 1037
rect 1161 1032 1190 1037
rect 1209 1032 1270 1037
rect 1489 1032 2718 1037
rect 2857 1032 3014 1037
rect 1313 1027 1398 1032
rect 361 1022 798 1027
rect 1113 1022 1222 1027
rect 1281 1022 1318 1027
rect 1393 1022 1422 1027
rect 1449 1022 1478 1027
rect 1721 1022 1750 1027
rect 1769 1022 1806 1027
rect 1817 1022 1886 1027
rect 1905 1022 1934 1027
rect 2017 1022 2206 1027
rect 2273 1022 2590 1027
rect 2889 1022 2966 1027
rect 3137 1022 3174 1027
rect 3273 1022 3374 1027
rect 793 1017 1118 1022
rect 1217 1017 1286 1022
rect 1553 1017 1630 1022
rect 2273 1017 2278 1022
rect 433 1012 454 1017
rect 465 1012 494 1017
rect 585 1012 614 1017
rect 1137 1012 1198 1017
rect 1329 1012 1374 1017
rect 1433 1012 1558 1017
rect 1625 1012 2214 1017
rect 2225 1012 2278 1017
rect 2297 1012 2878 1017
rect 97 992 142 997
rect 201 992 326 997
rect 345 992 382 997
rect 433 992 438 1012
rect 489 1007 590 1012
rect 753 1002 846 1007
rect 865 1002 950 1007
rect 977 1002 1062 1007
rect 865 997 870 1002
rect 457 992 526 997
rect 673 992 870 997
rect 945 997 950 1002
rect 945 992 974 997
rect 201 987 206 992
rect 65 982 118 987
rect 177 982 206 987
rect 321 987 326 992
rect 457 987 462 992
rect 321 982 462 987
rect 521 987 526 992
rect 521 982 550 987
rect 681 982 710 987
rect 793 982 822 987
rect 881 982 934 987
rect 945 982 998 987
rect 705 977 798 982
rect 1137 977 1142 1012
rect 2209 1007 2214 1012
rect 2873 1007 2878 1012
rect 2953 1012 2982 1017
rect 3257 1012 3286 1017
rect 2953 1007 2958 1012
rect 1169 1002 1486 1007
rect 1569 1002 1614 1007
rect 1697 1002 1926 1007
rect 1937 1002 2054 1007
rect 2209 1002 2318 1007
rect 2385 1002 2526 1007
rect 2873 1002 2958 1007
rect 3281 1007 3286 1012
rect 3361 1012 3390 1017
rect 3361 1007 3366 1012
rect 3281 1002 3366 1007
rect 2073 997 2182 1002
rect 1265 992 1886 997
rect 1953 992 2078 997
rect 2177 992 2622 997
rect 2641 992 2726 997
rect 2985 992 3158 997
rect 3233 992 3262 997
rect 2641 987 2646 992
rect 1161 982 1318 987
rect 1329 982 1742 987
rect 1753 982 1798 987
rect 2001 982 2398 987
rect 2409 982 2478 987
rect 2497 982 2646 987
rect 2721 987 2726 992
rect 2721 982 2958 987
rect 3081 982 3206 987
rect 3225 982 3350 987
rect 425 972 526 977
rect 545 972 582 977
rect 1137 972 1214 977
rect 233 967 398 972
rect 601 967 686 972
rect 1313 967 1318 982
rect 1817 977 1926 982
rect 1345 972 1822 977
rect 1921 972 2710 977
rect 2921 972 2958 977
rect 2729 967 2902 972
rect 2977 967 3078 972
rect 209 962 238 967
rect 393 962 606 967
rect 681 962 798 967
rect 809 962 966 967
rect 1017 962 1110 967
rect 1129 962 1166 967
rect 1313 962 1342 967
rect 1441 962 1470 967
rect 1481 962 1566 967
rect 1609 962 1670 967
rect 1745 962 1790 967
rect 1825 962 1910 967
rect 2033 962 2078 967
rect 2137 962 2414 967
rect 2425 962 2454 967
rect 2473 962 2550 967
rect 2705 962 2734 967
rect 2897 962 2982 967
rect 3073 962 3102 967
rect 1017 957 1022 962
rect 81 952 382 957
rect 449 952 670 957
rect 937 952 1022 957
rect 1105 957 1110 962
rect 1337 957 1446 962
rect 1105 952 1278 957
rect 1625 952 2774 957
rect 2809 952 3094 957
rect 3193 952 3222 957
rect 201 942 278 947
rect 401 942 518 947
rect 561 942 590 947
rect 585 937 590 942
rect 665 942 694 947
rect 777 942 838 947
rect 849 942 1430 947
rect 1473 942 1694 947
rect 1777 942 1902 947
rect 1921 942 2030 947
rect 2049 942 2110 947
rect 2161 942 2270 947
rect 2289 942 2310 947
rect 2353 942 2550 947
rect 2577 942 2654 947
rect 2865 942 2974 947
rect 3073 942 3134 947
rect 3153 942 3270 947
rect 3337 942 3390 947
rect 665 937 670 942
rect 2289 937 2294 942
rect 2577 937 2582 942
rect 2969 937 3078 942
rect 3153 937 3158 942
rect 585 932 670 937
rect 841 932 1942 937
rect 1961 932 2006 937
rect 2017 932 2046 937
rect 2081 932 2374 937
rect 2441 932 2582 937
rect 2753 932 2942 937
rect 3097 932 3158 937
rect 3209 932 3374 937
rect 1937 927 1942 932
rect 105 922 230 927
rect 689 922 726 927
rect 793 922 854 927
rect 937 922 1366 927
rect 1465 922 1502 927
rect 1529 922 1670 927
rect 1793 922 1902 927
rect 1937 922 2038 927
rect 2225 922 2366 927
rect 2577 922 2606 927
rect 2833 922 3030 927
rect 225 917 230 922
rect 305 917 406 922
rect 2057 917 2206 922
rect 2385 917 2558 922
rect 3025 917 3030 922
rect 3113 922 3142 927
rect 3241 922 3294 927
rect 3321 922 3350 927
rect 3113 917 3118 922
rect 225 912 262 917
rect 281 912 310 917
rect 401 912 430 917
rect 513 912 534 917
rect 625 912 734 917
rect 833 912 870 917
rect 1009 912 1078 917
rect 1129 912 1198 917
rect 1217 912 1350 917
rect 1417 912 1638 917
rect 1713 912 2062 917
rect 2201 912 2390 917
rect 2553 912 2822 917
rect 3025 912 3118 917
rect 3137 912 3142 922
rect 345 902 374 907
rect 505 902 598 907
rect 633 902 1366 907
rect 1425 902 1526 907
rect 1641 902 1958 907
rect 1993 902 2094 907
rect 2129 902 2198 907
rect 2265 902 2630 907
rect 1521 897 1646 902
rect 2193 897 2198 902
rect 281 892 366 897
rect 577 892 886 897
rect 969 892 1070 897
rect 1081 892 1502 897
rect 1665 892 1766 897
rect 1905 892 2182 897
rect 2193 892 2334 897
rect 2385 892 2574 897
rect 2617 892 2686 897
rect 3297 892 3406 897
rect 1785 887 1886 892
rect 393 882 486 887
rect 521 882 774 887
rect 817 882 862 887
rect 945 882 1550 887
rect 1609 882 1790 887
rect 1881 882 2062 887
rect 2081 882 2222 887
rect 2305 882 2350 887
rect 2441 882 2670 887
rect 265 877 398 882
rect 481 877 486 882
rect 241 872 270 877
rect 481 872 958 877
rect 1089 872 2198 877
rect 2569 872 2726 877
rect 2905 872 2950 877
rect 953 867 1094 872
rect 2217 867 2414 872
rect 297 862 630 867
rect 673 862 934 867
rect 1113 862 1150 867
rect 1161 862 2222 867
rect 2409 862 2702 867
rect 2889 862 2942 867
rect 321 852 894 857
rect 1009 852 1086 857
rect 1105 852 1630 857
rect 1705 852 1814 857
rect 1825 852 2246 857
rect 2281 852 2398 857
rect 2505 852 2902 857
rect 1009 847 1014 852
rect 217 842 270 847
rect 321 842 582 847
rect 641 842 694 847
rect 753 842 798 847
rect 857 842 974 847
rect 985 842 1014 847
rect 1081 847 1086 852
rect 1081 842 1206 847
rect 1249 842 1574 847
rect 1625 842 1702 847
rect 1849 842 1942 847
rect 2057 842 2086 847
rect 2113 842 2518 847
rect 2609 842 2686 847
rect 2841 842 2926 847
rect 321 837 326 842
rect 641 837 646 842
rect 1721 837 1830 842
rect 2513 837 2614 842
rect 137 832 166 837
rect 225 832 326 837
rect 337 832 422 837
rect 441 832 470 837
rect 489 832 582 837
rect 609 832 646 837
rect 665 832 694 837
rect 825 832 1134 837
rect 1193 832 1534 837
rect 1585 832 1726 837
rect 1825 832 1878 837
rect 2049 832 2190 837
rect 2241 832 2278 837
rect 2313 832 2494 837
rect 3289 832 3406 837
rect 689 827 830 832
rect 401 822 510 827
rect 545 822 638 827
rect 849 822 1006 827
rect 1033 822 1390 827
rect 1449 822 2006 827
rect 2033 822 2462 827
rect 2513 822 2606 827
rect 2513 817 2518 822
rect 209 812 278 817
rect 313 812 358 817
rect 625 812 654 817
rect 273 807 278 812
rect 649 807 654 812
rect 761 812 1278 817
rect 1289 812 1310 817
rect 1321 812 2518 817
rect 2601 817 2606 822
rect 2601 812 2630 817
rect 761 807 766 812
rect 113 802 254 807
rect 273 802 374 807
rect 417 802 438 807
rect 457 802 542 807
rect 649 802 766 807
rect 785 802 894 807
rect 913 802 1254 807
rect 1273 802 1278 812
rect 1305 807 1310 812
rect 1305 802 1494 807
rect 1569 802 1846 807
rect 1945 802 2022 807
rect 2057 802 2134 807
rect 2185 802 2246 807
rect 2257 802 2622 807
rect 457 797 462 802
rect 153 792 182 797
rect 289 792 462 797
rect 537 797 542 802
rect 537 792 566 797
rect 993 792 1126 797
rect 1137 792 1950 797
rect 2057 792 2614 797
rect 2657 792 2662 817
rect 2729 812 2806 817
rect 2929 812 3126 817
rect 2929 807 2934 812
rect 2713 802 2774 807
rect 2905 802 2934 807
rect 3121 807 3126 812
rect 3121 802 3150 807
rect 3361 802 3390 807
rect 2777 792 2894 797
rect 3049 792 3094 797
rect 177 787 294 792
rect 1945 787 2062 792
rect 313 782 622 787
rect 889 782 974 787
rect 1089 782 1206 787
rect 1265 782 1486 787
rect 1529 782 1622 787
rect 1745 782 1854 787
rect 1881 782 1926 787
rect 2081 782 2190 787
rect 2249 782 2350 787
rect 2457 782 2478 787
rect 2585 782 2718 787
rect 2729 782 2758 787
rect 889 777 894 782
rect 169 772 398 777
rect 425 772 614 777
rect 633 772 670 777
rect 689 772 846 777
rect 865 772 894 777
rect 969 777 974 782
rect 2753 777 2758 782
rect 2873 782 3046 787
rect 3097 782 3206 787
rect 2873 777 2878 782
rect 969 772 1078 777
rect 1193 772 1518 777
rect 1569 772 1614 777
rect 1705 772 2398 777
rect 2753 772 2878 777
rect 3089 772 3142 777
rect 3265 772 3294 777
rect 689 767 694 772
rect 337 762 526 767
rect 625 762 694 767
rect 841 767 846 772
rect 1073 767 1198 772
rect 3089 767 3094 772
rect 841 762 966 767
rect 1217 762 1326 767
rect 1369 762 1702 767
rect 1825 762 1974 767
rect 2185 762 2462 767
rect 2913 762 3094 767
rect 3105 762 3270 767
rect 713 757 822 762
rect 1993 757 2166 762
rect 81 752 110 757
rect 409 752 478 757
rect 569 752 718 757
rect 817 752 934 757
rect 1009 752 1062 757
rect 1089 752 1406 757
rect 1481 752 1590 757
rect 1665 752 1998 757
rect 2161 752 2342 757
rect 2393 752 2510 757
rect 3113 752 3134 757
rect 1009 747 1014 752
rect 2881 747 3046 752
rect 113 742 166 747
rect 233 742 342 747
rect 393 742 422 747
rect 465 742 558 747
rect 649 742 678 747
rect 705 742 758 747
rect 801 742 1014 747
rect 1137 742 1310 747
rect 1601 742 2206 747
rect 2225 742 2294 747
rect 2305 742 2382 747
rect 2417 742 2438 747
rect 2449 742 2510 747
rect 2537 742 2566 747
rect 2689 742 2734 747
rect 2857 742 2886 747
rect 3041 742 3094 747
rect 3113 742 3190 747
rect 3225 742 3358 747
rect 337 737 342 742
rect 553 737 654 742
rect 1137 737 1142 742
rect 1329 737 1582 742
rect 2225 737 2230 742
rect 81 732 142 737
rect 337 732 510 737
rect 689 732 726 737
rect 1057 732 1142 737
rect 1161 732 1334 737
rect 1577 732 1646 737
rect 1681 732 1886 737
rect 1977 732 2030 737
rect 2081 732 2230 737
rect 2289 737 2294 742
rect 3089 737 3094 742
rect 2289 732 2454 737
rect 745 727 942 732
rect 2545 727 2550 737
rect 2737 732 3022 737
rect 3089 732 3166 737
rect 3281 732 3342 737
rect 377 722 422 727
rect 577 722 646 727
rect 681 722 750 727
rect 937 722 1358 727
rect 1385 722 1486 727
rect 1513 722 1598 727
rect 1825 722 2550 727
rect 3017 722 3022 732
rect 3137 722 3166 727
rect 1633 717 1806 722
rect 3161 717 3166 722
rect 3281 722 3350 727
rect 3281 717 3286 722
rect 65 712 134 717
rect 233 712 342 717
rect 353 712 430 717
rect 625 712 926 717
rect 1033 712 1150 717
rect 1201 712 1278 717
rect 1345 712 1526 717
rect 921 707 1038 712
rect 1521 707 1526 712
rect 1609 712 1638 717
rect 1801 712 2286 717
rect 2297 712 2382 717
rect 2473 712 2542 717
rect 3161 712 3286 717
rect 3321 712 3366 717
rect 1609 707 1614 712
rect 65 702 254 707
rect 489 702 510 707
rect 521 702 614 707
rect 713 702 822 707
rect 857 702 902 707
rect 1057 702 1126 707
rect 1177 702 1230 707
rect 1249 702 1334 707
rect 1409 702 1502 707
rect 1521 702 1614 707
rect 1657 702 2086 707
rect 2361 702 2446 707
rect 2457 702 2518 707
rect 2569 702 2742 707
rect 2969 702 3054 707
rect 3313 702 3358 707
rect 337 697 438 702
rect 609 697 718 702
rect 2209 697 2342 702
rect 313 692 342 697
rect 433 692 590 697
rect 737 692 870 697
rect 1009 692 1142 697
rect 1201 692 1470 697
rect 1713 692 1774 697
rect 1873 692 2062 697
rect 2153 692 2174 697
rect 2185 692 2214 697
rect 2337 692 2470 697
rect 2497 692 2550 697
rect 1201 687 1206 692
rect 209 682 422 687
rect 593 682 662 687
rect 737 682 774 687
rect 1041 682 1110 687
rect 1145 682 1206 687
rect 1217 682 1382 687
rect 1521 682 1566 687
rect 1657 682 1798 687
rect 2129 682 2406 687
rect 793 677 886 682
rect 2001 677 2110 682
rect 2465 677 2470 692
rect 2569 687 2574 702
rect 2489 682 2574 687
rect 2737 687 2742 702
rect 2737 682 2934 687
rect 313 672 494 677
rect 753 672 798 677
rect 881 672 910 677
rect 937 672 1206 677
rect 1225 672 1318 677
rect 1385 672 1430 677
rect 1489 672 1534 677
rect 1553 672 2006 677
rect 2105 672 2398 677
rect 2465 672 2590 677
rect 2601 672 2726 677
rect 513 667 734 672
rect 1553 667 1558 672
rect 329 662 398 667
rect 473 662 518 667
rect 729 662 1302 667
rect 1313 662 1558 667
rect 1569 662 1590 667
rect 1617 662 1766 667
rect 1985 662 2230 667
rect 2289 662 2358 667
rect 2521 662 2550 667
rect 1585 657 1590 662
rect 1785 657 1966 662
rect 2545 657 2550 662
rect 2609 662 2638 667
rect 2609 657 2614 662
rect 177 652 238 657
rect 505 652 1078 657
rect 1105 652 1574 657
rect 1585 652 1790 657
rect 1961 652 2006 657
rect 2073 652 2438 657
rect 2449 652 2494 657
rect 2545 652 2614 657
rect 409 647 510 652
rect 1105 647 1110 652
rect 129 642 230 647
rect 321 642 414 647
rect 641 642 1038 647
rect 1081 642 1110 647
rect 1121 642 1390 647
rect 1449 642 1902 647
rect 1921 642 2006 647
rect 2033 642 2118 647
rect 2169 642 2390 647
rect 137 632 222 637
rect 321 627 326 642
rect 561 637 646 642
rect 2449 637 2454 652
rect 3225 642 3326 647
rect 489 632 566 637
rect 665 632 702 637
rect 769 632 2454 637
rect 2537 632 2654 637
rect 2929 632 3014 637
rect 3297 632 3342 637
rect 161 622 230 627
rect 289 622 326 627
rect 361 622 510 627
rect 633 622 918 627
rect 1129 622 1286 627
rect 1329 622 1446 627
rect 1497 622 1558 627
rect 1609 622 1710 627
rect 1769 622 1942 627
rect 2073 622 2150 627
rect 2161 622 2198 627
rect 2329 622 2358 627
rect 1553 617 1558 622
rect 1953 617 2078 622
rect 2217 617 2310 622
rect 2353 617 2358 622
rect 2433 622 2566 627
rect 2433 617 2438 622
rect 2929 617 2934 632
rect 3169 622 3254 627
rect 209 612 270 617
rect 281 612 446 617
rect 641 612 694 617
rect 817 612 942 617
rect 1049 612 1150 617
rect 1169 612 1270 617
rect 1313 612 1342 617
rect 1353 612 1374 617
rect 1553 612 1606 617
rect 1665 612 1958 617
rect 2097 612 2222 617
rect 2305 612 2334 617
rect 2353 612 2438 617
rect 2449 612 2582 617
rect 2865 612 2934 617
rect 2953 612 3414 617
rect 2577 607 2582 612
rect 193 602 398 607
rect 545 602 630 607
rect 705 602 1502 607
rect 1761 602 1870 607
rect 1881 602 1958 607
rect 2033 602 2278 607
rect 2409 602 2494 607
rect 2577 602 2646 607
rect 2673 602 2702 607
rect 3385 602 3430 607
rect 625 597 710 602
rect 137 592 326 597
rect 729 592 806 597
rect 905 592 1206 597
rect 1217 592 1302 597
rect 1313 592 1494 597
rect 1585 592 1958 597
rect 2049 592 2134 597
rect 2233 592 2286 597
rect 2305 592 2438 597
rect 2529 592 2590 597
rect 2833 592 3030 597
rect 3049 592 3206 597
rect 801 587 910 592
rect 1297 587 1302 592
rect 2129 587 2134 592
rect 177 582 278 587
rect 337 582 526 587
rect 585 582 638 587
rect 657 582 694 587
rect 761 582 782 587
rect 929 582 1014 587
rect 1065 582 1286 587
rect 1297 582 1398 587
rect 1737 582 1798 587
rect 1857 582 2110 587
rect 2129 582 2342 587
rect 2353 582 2430 587
rect 2585 582 2614 587
rect 2977 582 3046 587
rect 273 577 342 582
rect 169 572 246 577
rect 497 572 526 577
rect 689 572 814 577
rect 833 572 1046 577
rect 1129 572 1254 577
rect 545 567 646 572
rect 1281 567 1286 582
rect 1441 577 1718 582
rect 3041 577 3046 582
rect 3153 582 3414 587
rect 3153 577 3158 582
rect 1329 572 1374 577
rect 1417 572 1446 577
rect 1713 572 1766 577
rect 1817 572 2094 577
rect 2201 572 2246 577
rect 2329 572 2542 577
rect 2577 572 2710 577
rect 2745 572 3022 577
rect 3041 572 3158 577
rect 369 562 550 567
rect 641 562 822 567
rect 1001 562 1062 567
rect 1089 562 1190 567
rect 1281 562 2462 567
rect 849 557 982 562
rect 329 552 366 557
rect 385 552 630 557
rect 825 552 854 557
rect 977 552 1030 557
rect 1049 552 1078 557
rect 1201 552 1246 557
rect 1257 552 2470 557
rect 2801 552 2870 557
rect 385 547 390 552
rect 649 547 806 552
rect 89 542 166 547
rect 313 542 390 547
rect 401 542 654 547
rect 801 542 1966 547
rect 2081 542 2134 547
rect 2153 542 2374 547
rect 2473 542 2502 547
rect 2537 542 2614 547
rect 2961 542 3046 547
rect 3217 542 3438 547
rect 393 532 582 537
rect 625 532 830 537
rect 905 532 1134 537
rect 1169 532 1622 537
rect 1641 532 1774 537
rect 1865 532 2166 537
rect 2177 532 2222 537
rect 2257 532 2462 537
rect 2545 532 2582 537
rect 1769 527 1870 532
rect 2177 527 2182 532
rect 2457 527 2550 532
rect 321 522 406 527
rect 633 522 838 527
rect 945 522 1430 527
rect 1553 522 1750 527
rect 1889 522 1982 527
rect 2009 522 2134 527
rect 2161 522 2182 527
rect 2569 522 2718 527
rect 425 517 614 522
rect 217 512 278 517
rect 313 512 430 517
rect 609 512 670 517
rect 865 512 1006 517
rect 1073 512 1142 517
rect 1193 512 1414 517
rect 689 507 790 512
rect 1425 507 1430 522
rect 2961 517 2966 542
rect 3041 537 3046 542
rect 3041 532 3310 537
rect 3025 522 3174 527
rect 3249 522 3310 527
rect 1441 512 1566 517
rect 1601 512 1686 517
rect 1865 512 1902 517
rect 1961 512 2030 517
rect 2081 512 2166 517
rect 2241 512 2278 517
rect 2345 512 2422 517
rect 2505 512 2638 517
rect 2697 512 2830 517
rect 2881 512 2966 517
rect 3009 512 3126 517
rect 1705 507 1822 512
rect 2241 507 2246 512
rect 3169 507 3174 522
rect 3273 512 3382 517
rect 3273 507 3278 512
rect 113 502 142 507
rect 441 502 694 507
rect 785 502 1342 507
rect 1425 502 1710 507
rect 1817 502 2086 507
rect 2153 502 2246 507
rect 2337 502 2406 507
rect 2457 502 2518 507
rect 2721 502 2750 507
rect 3169 502 3278 507
rect 3297 502 3430 507
rect 2513 497 2726 502
rect 193 492 254 497
rect 521 492 822 497
rect 833 492 2046 497
rect 2193 492 2222 497
rect 2385 492 2494 497
rect 249 487 254 492
rect 393 487 526 492
rect 2265 487 2366 492
rect 249 482 398 487
rect 561 482 1734 487
rect 1817 482 1974 487
rect 2177 482 2270 487
rect 2361 482 2438 487
rect 2489 482 2654 487
rect 417 472 1222 477
rect 1241 472 1414 477
rect 1457 472 1630 477
rect 1745 472 1958 477
rect 2137 472 2166 477
rect 2281 472 2342 477
rect 2929 472 3014 477
rect 2161 467 2286 472
rect 561 462 662 467
rect 721 462 886 467
rect 969 462 1270 467
rect 1385 462 1566 467
rect 1617 462 1814 467
rect 1921 462 2030 467
rect 2305 462 2558 467
rect 713 452 790 457
rect 801 452 950 457
rect 1089 452 1214 457
rect 1297 452 1542 457
rect 1569 452 1598 457
rect 1625 452 1886 457
rect 2073 452 2158 457
rect 2217 452 2390 457
rect 2529 452 2742 457
rect 609 447 718 452
rect 1569 447 1574 452
rect 1905 447 1982 452
rect 2073 447 2078 452
rect 153 442 286 447
rect 417 442 542 447
rect 417 437 422 442
rect 297 432 422 437
rect 537 437 542 442
rect 609 437 614 447
rect 737 442 766 447
rect 865 442 902 447
rect 985 442 1246 447
rect 1377 442 1422 447
rect 1441 442 1470 447
rect 1569 442 1910 447
rect 1977 442 2078 447
rect 2153 447 2158 452
rect 2153 442 2510 447
rect 1265 437 1358 442
rect 2505 437 2510 442
rect 537 432 614 437
rect 625 432 1174 437
rect 1225 432 1270 437
rect 1353 432 1638 437
rect 1729 432 1814 437
rect 1905 432 1966 437
rect 2089 432 2142 437
rect 2241 432 2334 437
rect 2505 432 2542 437
rect 1809 427 1910 432
rect 257 422 318 427
rect 625 422 734 427
rect 457 417 606 422
rect 753 417 758 427
rect 881 422 1790 427
rect 1929 422 2078 427
rect 2145 422 2230 427
rect 2313 422 2622 427
rect 3057 422 3206 427
rect 273 412 462 417
rect 601 412 838 417
rect 873 412 894 417
rect 905 412 942 417
rect 1201 412 1390 417
rect 1401 412 2422 417
rect 961 407 1142 412
rect 2417 407 2422 412
rect 2561 412 2590 417
rect 2601 412 2734 417
rect 2561 407 2566 412
rect 145 402 654 407
rect 689 402 966 407
rect 1137 402 1190 407
rect 1265 402 1294 407
rect 1377 402 1438 407
rect 1449 402 1606 407
rect 1617 402 1662 407
rect 1689 402 1846 407
rect 2417 402 2566 407
rect 3081 402 3238 407
rect 1185 397 1270 402
rect 1865 397 2230 402
rect 3081 397 3086 402
rect 297 392 358 397
rect 457 392 662 397
rect 681 392 806 397
rect 969 392 1126 397
rect 1385 392 1702 397
rect 1761 392 1870 397
rect 2225 392 2254 397
rect 2369 392 2398 397
rect 2809 392 2966 397
rect 3057 392 3086 397
rect 3233 397 3238 402
rect 3233 392 3262 397
rect 833 387 950 392
rect 2961 387 2966 392
rect 513 382 718 387
rect 817 382 838 387
rect 945 382 982 387
rect 1097 382 1206 387
rect 1233 382 1366 387
rect 1401 382 1686 387
rect 1785 382 2574 387
rect 2961 382 3342 387
rect 401 377 494 382
rect 713 377 822 382
rect 1681 377 1790 382
rect 217 372 310 377
rect 377 372 406 377
rect 489 372 694 377
rect 849 372 1382 377
rect 1425 372 1662 377
rect 1809 372 2038 377
rect 2145 372 2174 377
rect 2361 372 2478 377
rect 2593 372 2942 377
rect 2593 367 2598 372
rect 2937 367 3102 372
rect 409 362 502 367
rect 561 362 750 367
rect 809 362 1350 367
rect 1369 362 1478 367
rect 1561 362 1638 367
rect 1681 362 1782 367
rect 1801 362 2134 367
rect 2273 362 2318 367
rect 2377 362 2406 367
rect 2489 362 2598 367
rect 3097 362 3422 367
rect 305 352 390 357
rect 425 352 670 357
rect 801 352 886 357
rect 969 352 1334 357
rect 1345 352 1350 362
rect 1473 357 1478 362
rect 1681 357 1686 362
rect 1473 352 1686 357
rect 1777 357 1782 362
rect 2129 357 2214 362
rect 2273 357 2278 362
rect 2401 357 2494 362
rect 2817 357 2918 362
rect 1777 352 1806 357
rect 2017 352 2102 357
rect 2209 352 2278 357
rect 2713 352 2822 357
rect 2913 352 3086 357
rect 305 347 310 352
rect 73 342 310 347
rect 385 347 390 352
rect 665 347 806 352
rect 881 347 974 352
rect 1345 347 1454 352
rect 1825 347 1974 352
rect 2529 347 2638 352
rect 385 342 646 347
rect 825 342 862 347
rect 1105 342 1182 347
rect 1249 342 1310 347
rect 1449 342 1478 347
rect 1497 342 1542 347
rect 1601 342 1726 347
rect 1745 342 1830 347
rect 1969 342 1998 347
rect 2033 342 2190 347
rect 2417 342 2534 347
rect 2633 342 2662 347
rect 2857 342 3014 347
rect 1745 337 1750 342
rect 3009 337 3014 342
rect 3073 342 3342 347
rect 3073 337 3078 342
rect 321 332 414 337
rect 441 332 1302 337
rect 1313 332 1470 337
rect 1521 332 1558 337
rect 1569 332 1750 337
rect 1809 332 2030 337
rect 2465 332 2502 337
rect 2569 332 2718 337
rect 3009 332 3078 337
rect 3385 332 3438 337
rect 1553 327 1558 332
rect 353 322 462 327
rect 497 322 614 327
rect 761 322 854 327
rect 1105 322 1278 327
rect 1353 322 1534 327
rect 1553 322 1646 327
rect 1729 322 1934 327
rect 1985 322 2118 327
rect 1009 317 1086 322
rect 329 312 438 317
rect 745 312 1014 317
rect 1081 312 1678 317
rect 1697 307 1830 312
rect 2113 307 2118 322
rect 2177 312 2238 317
rect 65 302 886 307
rect 1025 302 1166 307
rect 1281 302 1494 307
rect 1529 302 1702 307
rect 1825 302 1854 307
rect 1897 302 1982 307
rect 2001 302 2094 307
rect 2113 302 2166 307
rect 1025 297 1030 302
rect 2001 297 2006 302
rect 89 292 134 297
rect 393 292 446 297
rect 649 292 678 297
rect 897 292 1030 297
rect 1049 292 1142 297
rect 1249 292 1446 297
rect 1489 292 1550 297
rect 1569 292 2006 297
rect 2089 297 2094 302
rect 2177 297 2182 312
rect 2089 292 2182 297
rect 673 287 814 292
rect 897 287 902 292
rect 1569 287 1574 292
rect 465 282 630 287
rect 809 282 902 287
rect 1161 282 1574 287
rect 1585 282 1806 287
rect 1905 282 2246 287
rect 345 277 470 282
rect 625 277 630 282
rect 2321 277 2326 327
rect 2377 322 2526 327
rect 2617 322 2718 327
rect 2737 322 2782 327
rect 2417 312 2502 317
rect 2681 312 3342 317
rect 2353 302 2510 307
rect 2721 302 2814 307
rect 2809 297 2814 302
rect 3161 302 3190 307
rect 2705 292 2734 297
rect 2809 292 2966 297
rect 2961 287 2966 292
rect 3161 287 3166 302
rect 2961 282 3166 287
rect 3241 282 3310 287
rect 257 272 350 277
rect 625 272 790 277
rect 1417 272 1622 277
rect 2297 272 2406 277
rect 2809 272 2910 277
rect 489 267 606 272
rect 1281 267 1398 272
rect 1641 267 2278 272
rect 2809 267 2814 272
rect 361 262 494 267
rect 601 262 638 267
rect 721 262 910 267
rect 929 262 1006 267
rect 1153 262 1286 267
rect 1393 262 1646 267
rect 2273 262 2382 267
rect 2785 262 2814 267
rect 2905 267 2910 272
rect 2905 262 2942 267
rect 633 257 726 262
rect 929 257 934 262
rect 305 252 614 257
rect 305 247 310 252
rect 609 247 614 252
rect 745 252 934 257
rect 1001 257 1006 262
rect 1001 252 1030 257
rect 1297 252 2446 257
rect 2465 252 2742 257
rect 2825 252 2894 257
rect 745 247 750 252
rect 2465 247 2470 252
rect 233 242 310 247
rect 353 242 398 247
rect 609 242 750 247
rect 769 242 798 247
rect 889 242 1286 247
rect 1361 242 2470 247
rect 2737 247 2742 252
rect 2737 242 2766 247
rect 353 237 358 242
rect 417 237 510 242
rect 793 237 894 242
rect 97 232 358 237
rect 377 232 422 237
rect 505 232 590 237
rect 913 232 958 237
rect 1217 232 1350 237
rect 1537 232 1606 237
rect 1665 232 1702 237
rect 1721 232 1782 237
rect 1793 232 1846 237
rect 1889 232 2430 237
rect 2449 232 2518 237
rect 2537 232 2638 237
rect 2737 232 2782 237
rect 2833 232 2942 237
rect 3089 232 3182 237
rect 1425 227 1518 232
rect 2449 227 2454 232
rect 2537 227 2542 232
rect 193 222 222 227
rect 385 222 542 227
rect 833 222 950 227
rect 985 222 1062 227
rect 1249 222 1286 227
rect 1329 222 1430 227
rect 1513 222 2182 227
rect 2425 222 2454 227
rect 2489 222 2542 227
rect 2633 227 2638 232
rect 2633 222 2678 227
rect 2961 222 3070 227
rect 217 217 390 222
rect 2177 217 2430 222
rect 409 212 622 217
rect 825 212 1022 217
rect 1265 212 1342 217
rect 1441 212 1470 217
rect 1497 212 2030 217
rect 2121 212 2150 217
rect 2545 212 2622 217
rect 2913 212 3030 217
rect 1441 207 1446 212
rect 2025 207 2126 212
rect 225 202 438 207
rect 705 202 814 207
rect 1305 202 1446 207
rect 1457 202 1534 207
rect 1769 202 1982 207
rect 2153 202 2174 207
rect 545 197 686 202
rect 921 197 1038 202
rect 1553 197 1750 202
rect 2153 197 2158 202
rect 521 192 550 197
rect 681 192 726 197
rect 761 192 926 197
rect 1033 192 1454 197
rect 1473 192 1558 197
rect 1745 192 2158 197
rect 2169 197 2174 202
rect 2233 202 2446 207
rect 2625 202 2726 207
rect 2889 202 3078 207
rect 3321 202 3438 207
rect 2233 197 2238 202
rect 2169 192 2238 197
rect 2529 192 2614 197
rect 2777 192 2878 197
rect 2937 192 2966 197
rect 3073 192 3174 197
rect 3193 192 3334 197
rect 225 187 478 192
rect 2961 187 3078 192
rect 129 182 230 187
rect 473 182 502 187
rect 513 182 782 187
rect 937 182 1126 187
rect 1289 182 1718 187
rect 1729 182 1902 187
rect 1953 182 1990 187
rect 801 177 894 182
rect 1729 177 1734 182
rect 1953 177 1958 182
rect 89 172 118 177
rect 113 167 118 172
rect 241 172 542 177
rect 241 167 246 172
rect 537 167 542 172
rect 641 172 686 177
rect 745 172 806 177
rect 889 172 926 177
rect 985 172 1086 177
rect 1321 172 1550 177
rect 1633 172 1734 177
rect 1785 172 1854 177
rect 1905 172 1958 177
rect 1969 172 2150 177
rect 2305 172 2454 177
rect 2577 172 2766 177
rect 641 167 646 172
rect 921 167 990 172
rect 113 162 246 167
rect 281 162 382 167
rect 401 162 518 167
rect 537 162 646 167
rect 689 162 878 167
rect 1049 162 1142 167
rect 1241 162 1574 167
rect 1601 162 1742 167
rect 1825 162 1974 167
rect 2177 162 2286 167
rect 2305 157 2310 172
rect 265 152 358 157
rect 665 152 766 157
rect 889 152 1030 157
rect 1177 152 2310 157
rect 2449 157 2454 172
rect 2761 167 2766 172
rect 2873 172 3222 177
rect 2873 167 2878 172
rect 2761 162 2878 167
rect 2449 152 2526 157
rect 2897 152 2926 157
rect 481 147 566 152
rect 1049 147 1158 152
rect 2921 147 2926 152
rect 3033 152 3382 157
rect 3033 147 3038 152
rect 321 142 486 147
rect 561 142 902 147
rect 1001 142 1054 147
rect 1153 142 1302 147
rect 1393 142 1862 147
rect 1945 142 1982 147
rect 2129 142 2238 147
rect 2337 142 2438 147
rect 2921 142 3038 147
rect 3057 142 3094 147
rect 321 137 326 142
rect 2001 137 2110 142
rect 2233 137 2326 142
rect 225 132 326 137
rect 337 132 422 137
rect 497 132 550 137
rect 545 127 550 132
rect 697 132 766 137
rect 857 132 1166 137
rect 1201 132 1510 137
rect 1713 132 2006 137
rect 2105 132 2198 137
rect 2321 132 2510 137
rect 697 127 702 132
rect 1593 127 1694 132
rect 169 122 214 127
rect 209 117 214 122
rect 305 122 526 127
rect 545 122 702 127
rect 873 122 1030 127
rect 1041 122 1526 127
rect 1569 122 1598 127
rect 1689 122 1750 127
rect 1977 122 2030 127
rect 2057 122 2486 127
rect 2745 122 2902 127
rect 305 117 310 122
rect 1041 117 1046 122
rect 1521 117 1526 122
rect 1745 117 1982 122
rect 209 112 310 117
rect 329 112 430 117
rect 721 112 862 117
rect 937 112 1046 117
rect 1113 112 1502 117
rect 1521 112 1606 117
rect 1665 112 1726 117
rect 2385 112 2414 117
rect 2721 112 2782 117
rect 2873 112 2966 117
rect 857 107 942 112
rect 1665 107 1670 112
rect 2001 107 2254 112
rect 2385 107 2390 112
rect 1017 102 1110 107
rect 1161 102 1214 107
rect 1289 102 1318 107
rect 1401 102 1590 107
rect 1601 102 1670 107
rect 1697 102 1806 107
rect 1825 102 1966 107
rect 1985 102 2006 107
rect 2249 102 2390 107
rect 2849 102 2878 107
rect 1313 97 1406 102
rect 1601 97 1606 102
rect 1825 97 1830 102
rect 489 92 710 97
rect 705 87 710 92
rect 873 92 1046 97
rect 1425 92 1606 97
rect 1625 92 1830 97
rect 1961 97 1966 102
rect 2873 97 2878 102
rect 2961 102 2990 107
rect 2961 97 2966 102
rect 1961 92 2230 97
rect 2873 92 2966 97
rect 873 87 878 92
rect 1129 87 1262 92
rect 705 82 878 87
rect 1033 82 1134 87
rect 1257 82 1438 87
rect 1505 82 2350 87
rect 2417 82 2502 87
rect 921 77 998 82
rect 2417 77 2422 82
rect 897 72 926 77
rect 993 72 1022 77
rect 1145 72 1246 77
rect 1017 67 1150 72
rect 1241 67 1246 72
rect 1417 72 1766 77
rect 1953 72 2294 77
rect 1417 67 1422 72
rect 1761 67 1942 72
rect 2289 67 2294 72
rect 2361 72 2422 77
rect 2361 67 2366 72
rect 953 62 982 67
rect 977 57 982 62
rect 1177 62 1206 67
rect 1241 62 1422 67
rect 1937 62 1966 67
rect 2065 62 2142 67
rect 2241 62 2270 67
rect 2289 62 2366 67
rect 1177 57 1182 62
rect 1961 57 2070 62
rect 2137 57 2246 62
rect 569 52 942 57
rect 977 52 1182 57
rect 1537 52 1926 57
rect 937 37 942 52
rect 1537 47 1542 52
rect 1921 47 1926 52
rect 2089 52 2118 57
rect 2089 47 2094 52
rect 1217 42 1542 47
rect 1561 42 1590 47
rect 1921 42 2094 47
rect 2209 42 2238 47
rect 1217 37 1222 42
rect 937 32 1222 37
rect 1585 27 1590 42
rect 2209 37 2214 42
rect 2129 32 2214 37
rect 2129 27 2134 32
rect 1585 22 2134 27
use AND2X2  AND2X2_0
timestamp 1712256841
transform 1 0 2664 0 -1 1170
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1712256841
transform 1 0 1416 0 -1 1170
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1712256841
transform 1 0 2840 0 -1 170
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1712256841
transform 1 0 1440 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1712256841
transform 1 0 1400 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1712256841
transform 1 0 1320 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1712256841
transform 1 0 2304 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1712256841
transform 1 0 1584 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1712256841
transform 1 0 1024 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1712256841
transform 1 0 2608 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1712256841
transform 1 0 1000 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1712256841
transform 1 0 2672 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1712256841
transform 1 0 2688 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1712256841
transform 1 0 872 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1712256841
transform 1 0 2104 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1712256841
transform 1 0 1536 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1712256841
transform 1 0 1424 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1712256841
transform 1 0 1776 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1712256841
transform 1 0 80 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1712256841
transform 1 0 1112 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_20
timestamp 1712256841
transform 1 0 1712 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1712256841
transform 1 0 1000 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1712256841
transform 1 0 1560 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_23
timestamp 1712256841
transform 1 0 3128 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1712256841
transform 1 0 3216 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_25
timestamp 1712256841
transform 1 0 2704 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_26
timestamp 1712256841
transform 1 0 2752 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_27
timestamp 1712256841
transform 1 0 2048 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_28
timestamp 1712256841
transform 1 0 848 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_29
timestamp 1712256841
transform 1 0 2032 0 -1 3170
box -8 -3 40 105
use AND2X2  AND2X2_30
timestamp 1712256841
transform 1 0 3048 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_31
timestamp 1712256841
transform 1 0 2928 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_32
timestamp 1712256841
transform 1 0 1760 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_33
timestamp 1712256841
transform 1 0 688 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_34
timestamp 1712256841
transform 1 0 1192 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_35
timestamp 1712256841
transform 1 0 1488 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_36
timestamp 1712256841
transform 1 0 3280 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_37
timestamp 1712256841
transform 1 0 3248 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_38
timestamp 1712256841
transform 1 0 3240 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_39
timestamp 1712256841
transform 1 0 3336 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_40
timestamp 1712256841
transform 1 0 2872 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_41
timestamp 1712256841
transform 1 0 2928 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_42
timestamp 1712256841
transform 1 0 3056 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_43
timestamp 1712256841
transform 1 0 3296 0 1 570
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1712256841
transform 1 0 3192 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1712256841
transform 1 0 272 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1712256841
transform 1 0 480 0 -1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1712256841
transform 1 0 1712 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1712256841
transform 1 0 536 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1712256841
transform 1 0 2320 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1712256841
transform 1 0 624 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1712256841
transform 1 0 720 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1712256841
transform 1 0 392 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1712256841
transform 1 0 1952 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1712256841
transform 1 0 768 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1712256841
transform 1 0 2304 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1712256841
transform 1 0 96 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1712256841
transform 1 0 1192 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1712256841
transform 1 0 1928 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1712256841
transform 1 0 1128 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1712256841
transform 1 0 1264 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1712256841
transform 1 0 912 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1712256841
transform 1 0 824 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1712256841
transform 1 0 816 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1712256841
transform 1 0 1024 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1712256841
transform 1 0 1272 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1712256841
transform 1 0 1672 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1712256841
transform 1 0 1816 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1712256841
transform 1 0 1656 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1712256841
transform 1 0 1624 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1712256841
transform 1 0 1392 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_27
timestamp 1712256841
transform 1 0 2160 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_28
timestamp 1712256841
transform 1 0 2392 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_29
timestamp 1712256841
transform 1 0 2536 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_30
timestamp 1712256841
transform 1 0 2064 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_31
timestamp 1712256841
transform 1 0 3056 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_32
timestamp 1712256841
transform 1 0 2968 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_33
timestamp 1712256841
transform 1 0 2880 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_34
timestamp 1712256841
transform 1 0 2584 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_35
timestamp 1712256841
transform 1 0 2760 0 1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_36
timestamp 1712256841
transform 1 0 2528 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_37
timestamp 1712256841
transform 1 0 2624 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_38
timestamp 1712256841
transform 1 0 1800 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_39
timestamp 1712256841
transform 1 0 1752 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_40
timestamp 1712256841
transform 1 0 880 0 1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_41
timestamp 1712256841
transform 1 0 864 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_42
timestamp 1712256841
transform 1 0 2616 0 1 2970
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1712256841
transform 1 0 1472 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1712256841
transform 1 0 1000 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1712256841
transform 1 0 648 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1712256841
transform 1 0 1024 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1712256841
transform 1 0 272 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1712256841
transform 1 0 176 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1712256841
transform 1 0 200 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1712256841
transform 1 0 2232 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1712256841
transform 1 0 2312 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1712256841
transform 1 0 2072 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1712256841
transform 1 0 1000 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1712256841
transform 1 0 2208 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1712256841
transform 1 0 1592 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1712256841
transform 1 0 776 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1712256841
transform 1 0 392 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1712256841
transform 1 0 384 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1712256841
transform 1 0 432 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1712256841
transform 1 0 960 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1712256841
transform 1 0 424 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1712256841
transform 1 0 2120 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1712256841
transform 1 0 1720 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1712256841
transform 1 0 1960 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1712256841
transform 1 0 2520 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1712256841
transform 1 0 2616 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1712256841
transform 1 0 1008 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1712256841
transform 1 0 496 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1712256841
transform 1 0 464 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1712256841
transform 1 0 704 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1712256841
transform 1 0 984 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1712256841
transform 1 0 512 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1712256841
transform 1 0 1936 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1712256841
transform 1 0 2440 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1712256841
transform 1 0 2416 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1712256841
transform 1 0 2136 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1712256841
transform 1 0 1608 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1712256841
transform 1 0 1240 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1712256841
transform 1 0 864 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1712256841
transform 1 0 672 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1712256841
transform 1 0 928 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1712256841
transform 1 0 552 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1712256841
transform 1 0 568 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1712256841
transform 1 0 1384 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1712256841
transform 1 0 2208 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1712256841
transform 1 0 1928 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1712256841
transform 1 0 2384 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1712256841
transform 1 0 2000 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1712256841
transform 1 0 1592 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1712256841
transform 1 0 400 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1712256841
transform 1 0 1448 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1712256841
transform 1 0 368 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1712256841
transform 1 0 328 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1712256841
transform 1 0 352 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1712256841
transform 1 0 2592 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1712256841
transform 1 0 2128 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1712256841
transform 1 0 1816 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_55
timestamp 1712256841
transform 1 0 1240 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1712256841
transform 1 0 2472 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_57
timestamp 1712256841
transform 1 0 1600 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_58
timestamp 1712256841
transform 1 0 2200 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_59
timestamp 1712256841
transform 1 0 1984 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_60
timestamp 1712256841
transform 1 0 2224 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_61
timestamp 1712256841
transform 1 0 2008 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_62
timestamp 1712256841
transform 1 0 200 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_63
timestamp 1712256841
transform 1 0 688 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_64
timestamp 1712256841
transform 1 0 240 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_65
timestamp 1712256841
transform 1 0 88 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_66
timestamp 1712256841
transform 1 0 392 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_67
timestamp 1712256841
transform 1 0 280 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_68
timestamp 1712256841
transform 1 0 344 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_69
timestamp 1712256841
transform 1 0 408 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_70
timestamp 1712256841
transform 1 0 1456 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_71
timestamp 1712256841
transform 1 0 1312 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1712256841
transform 1 0 2392 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_73
timestamp 1712256841
transform 1 0 1800 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_74
timestamp 1712256841
transform 1 0 2256 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_75
timestamp 1712256841
transform 1 0 2384 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_76
timestamp 1712256841
transform 1 0 144 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_77
timestamp 1712256841
transform 1 0 720 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_78
timestamp 1712256841
transform 1 0 136 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_79
timestamp 1712256841
transform 1 0 176 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_80
timestamp 1712256841
transform 1 0 1096 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_81
timestamp 1712256841
transform 1 0 1904 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_82
timestamp 1712256841
transform 1 0 2136 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_83
timestamp 1712256841
transform 1 0 2208 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_84
timestamp 1712256841
transform 1 0 1576 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_85
timestamp 1712256841
transform 1 0 1880 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_86
timestamp 1712256841
transform 1 0 1496 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_87
timestamp 1712256841
transform 1 0 1592 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_88
timestamp 1712256841
transform 1 0 1208 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_89
timestamp 1712256841
transform 1 0 1408 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_90
timestamp 1712256841
transform 1 0 1128 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_91
timestamp 1712256841
transform 1 0 1352 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_92
timestamp 1712256841
transform 1 0 920 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_93
timestamp 1712256841
transform 1 0 1008 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_94
timestamp 1712256841
transform 1 0 1352 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_95
timestamp 1712256841
transform 1 0 1296 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_96
timestamp 1712256841
transform 1 0 720 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_97
timestamp 1712256841
transform 1 0 936 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_98
timestamp 1712256841
transform 1 0 576 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_99
timestamp 1712256841
transform 1 0 576 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_100
timestamp 1712256841
transform 1 0 416 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_101
timestamp 1712256841
transform 1 0 552 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_102
timestamp 1712256841
transform 1 0 344 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_103
timestamp 1712256841
transform 1 0 232 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_104
timestamp 1712256841
transform 1 0 344 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_105
timestamp 1712256841
transform 1 0 544 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_106
timestamp 1712256841
transform 1 0 168 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_107
timestamp 1712256841
transform 1 0 88 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_108
timestamp 1712256841
transform 1 0 416 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_109
timestamp 1712256841
transform 1 0 552 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_110
timestamp 1712256841
transform 1 0 192 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_111
timestamp 1712256841
transform 1 0 88 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_112
timestamp 1712256841
transform 1 0 1064 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_113
timestamp 1712256841
transform 1 0 416 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_114
timestamp 1712256841
transform 1 0 552 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_115
timestamp 1712256841
transform 1 0 272 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_116
timestamp 1712256841
transform 1 0 88 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_117
timestamp 1712256841
transform 1 0 456 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_118
timestamp 1712256841
transform 1 0 496 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_119
timestamp 1712256841
transform 1 0 208 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_120
timestamp 1712256841
transform 1 0 88 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_121
timestamp 1712256841
transform 1 0 432 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_122
timestamp 1712256841
transform 1 0 496 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_123
timestamp 1712256841
transform 1 0 144 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_124
timestamp 1712256841
transform 1 0 88 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_125
timestamp 1712256841
transform 1 0 392 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_126
timestamp 1712256841
transform 1 0 600 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_127
timestamp 1712256841
transform 1 0 200 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_128
timestamp 1712256841
transform 1 0 88 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_129
timestamp 1712256841
transform 1 0 392 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_130
timestamp 1712256841
transform 1 0 768 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_131
timestamp 1712256841
transform 1 0 232 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_132
timestamp 1712256841
transform 1 0 136 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_133
timestamp 1712256841
transform 1 0 472 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_134
timestamp 1712256841
transform 1 0 616 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_135
timestamp 1712256841
transform 1 0 320 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_136
timestamp 1712256841
transform 1 0 496 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_137
timestamp 1712256841
transform 1 0 960 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_138
timestamp 1712256841
transform 1 0 920 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_139
timestamp 1712256841
transform 1 0 920 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_140
timestamp 1712256841
transform 1 0 808 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_141
timestamp 1712256841
transform 1 0 1096 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_142
timestamp 1712256841
transform 1 0 1096 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_143
timestamp 1712256841
transform 1 0 1168 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_144
timestamp 1712256841
transform 1 0 1120 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_145
timestamp 1712256841
transform 1 0 1040 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_146
timestamp 1712256841
transform 1 0 1296 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_147
timestamp 1712256841
transform 1 0 1448 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_148
timestamp 1712256841
transform 1 0 1440 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_149
timestamp 1712256841
transform 1 0 1488 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_150
timestamp 1712256841
transform 1 0 1848 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_151
timestamp 1712256841
transform 1 0 1808 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_152
timestamp 1712256841
transform 1 0 1760 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_153
timestamp 1712256841
transform 1 0 1720 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_154
timestamp 1712256841
transform 1 0 2120 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_155
timestamp 1712256841
transform 1 0 2040 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_156
timestamp 1712256841
transform 1 0 2312 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_157
timestamp 1712256841
transform 1 0 2144 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_158
timestamp 1712256841
transform 1 0 2480 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_159
timestamp 1712256841
transform 1 0 2280 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_160
timestamp 1712256841
transform 1 0 2288 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_161
timestamp 1712256841
transform 1 0 2200 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_162
timestamp 1712256841
transform 1 0 2504 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_163
timestamp 1712256841
transform 1 0 2344 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_164
timestamp 1712256841
transform 1 0 2384 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_165
timestamp 1712256841
transform 1 0 2216 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_166
timestamp 1712256841
transform 1 0 2456 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_167
timestamp 1712256841
transform 1 0 2368 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_168
timestamp 1712256841
transform 1 0 2160 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_169
timestamp 1712256841
transform 1 0 2080 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_170
timestamp 1712256841
transform 1 0 2592 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_171
timestamp 1712256841
transform 1 0 2400 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_172
timestamp 1712256841
transform 1 0 2248 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_173
timestamp 1712256841
transform 1 0 2128 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_174
timestamp 1712256841
transform 1 0 1600 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_175
timestamp 1712256841
transform 1 0 1720 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_176
timestamp 1712256841
transform 1 0 1664 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_177
timestamp 1712256841
transform 1 0 1816 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_178
timestamp 1712256841
transform 1 0 1776 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_179
timestamp 1712256841
transform 1 0 1768 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_180
timestamp 1712256841
transform 1 0 1896 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_181
timestamp 1712256841
transform 1 0 1984 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_182
timestamp 1712256841
transform 1 0 1864 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_183
timestamp 1712256841
transform 1 0 1808 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_184
timestamp 1712256841
transform 1 0 2200 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_185
timestamp 1712256841
transform 1 0 2240 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_186
timestamp 1712256841
transform 1 0 2168 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_187
timestamp 1712256841
transform 1 0 2144 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_188
timestamp 1712256841
transform 1 0 2312 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_189
timestamp 1712256841
transform 1 0 2344 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_190
timestamp 1712256841
transform 1 0 2392 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_191
timestamp 1712256841
transform 1 0 2288 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_192
timestamp 1712256841
transform 1 0 2472 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_193
timestamp 1712256841
transform 1 0 2008 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_194
timestamp 1712256841
transform 1 0 1648 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_195
timestamp 1712256841
transform 1 0 2648 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_196
timestamp 1712256841
transform 1 0 2976 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_197
timestamp 1712256841
transform 1 0 2944 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_198
timestamp 1712256841
transform 1 0 3080 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_199
timestamp 1712256841
transform 1 0 3064 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_200
timestamp 1712256841
transform 1 0 2952 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_201
timestamp 1712256841
transform 1 0 2832 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_202
timestamp 1712256841
transform 1 0 2752 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_203
timestamp 1712256841
transform 1 0 2736 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_204
timestamp 1712256841
transform 1 0 2904 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_205
timestamp 1712256841
transform 1 0 2968 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_206
timestamp 1712256841
transform 1 0 3152 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_207
timestamp 1712256841
transform 1 0 3320 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_208
timestamp 1712256841
transform 1 0 3368 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_209
timestamp 1712256841
transform 1 0 3232 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_210
timestamp 1712256841
transform 1 0 2536 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_211
timestamp 1712256841
transform 1 0 2392 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_212
timestamp 1712256841
transform 1 0 2008 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_213
timestamp 1712256841
transform 1 0 2328 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_214
timestamp 1712256841
transform 1 0 2288 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_215
timestamp 1712256841
transform 1 0 2304 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_216
timestamp 1712256841
transform 1 0 2208 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_217
timestamp 1712256841
transform 1 0 2248 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_218
timestamp 1712256841
transform 1 0 2072 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_219
timestamp 1712256841
transform 1 0 2152 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_220
timestamp 1712256841
transform 1 0 1792 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_221
timestamp 1712256841
transform 1 0 1792 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_222
timestamp 1712256841
transform 1 0 1888 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_223
timestamp 1712256841
transform 1 0 1896 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_224
timestamp 1712256841
transform 1 0 1648 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_225
timestamp 1712256841
transform 1 0 1688 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_226
timestamp 1712256841
transform 1 0 1592 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_227
timestamp 1712256841
transform 1 0 1688 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_228
timestamp 1712256841
transform 1 0 1432 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_229
timestamp 1712256841
transform 1 0 1624 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_230
timestamp 1712256841
transform 1 0 1328 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_231
timestamp 1712256841
transform 1 0 1584 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_232
timestamp 1712256841
transform 1 0 1304 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_233
timestamp 1712256841
transform 1 0 1592 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_234
timestamp 1712256841
transform 1 0 1224 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_235
timestamp 1712256841
transform 1 0 1520 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_236
timestamp 1712256841
transform 1 0 1200 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_237
timestamp 1712256841
transform 1 0 1168 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_238
timestamp 1712256841
transform 1 0 1000 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_239
timestamp 1712256841
transform 1 0 1064 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_240
timestamp 1712256841
transform 1 0 608 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_241
timestamp 1712256841
transform 1 0 1144 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_242
timestamp 1712256841
transform 1 0 736 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_243
timestamp 1712256841
transform 1 0 1040 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_244
timestamp 1712256841
transform 1 0 584 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_245
timestamp 1712256841
transform 1 0 720 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_246
timestamp 1712256841
transform 1 0 512 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_247
timestamp 1712256841
transform 1 0 648 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_248
timestamp 1712256841
transform 1 0 504 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_249
timestamp 1712256841
transform 1 0 616 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_250
timestamp 1712256841
transform 1 0 544 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_251
timestamp 1712256841
transform 1 0 664 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_252
timestamp 1712256841
transform 1 0 720 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_253
timestamp 1712256841
transform 1 0 792 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_254
timestamp 1712256841
transform 1 0 624 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_255
timestamp 1712256841
transform 1 0 720 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_256
timestamp 1712256841
transform 1 0 880 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_257
timestamp 1712256841
transform 1 0 784 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_258
timestamp 1712256841
transform 1 0 968 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_259
timestamp 1712256841
transform 1 0 824 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_260
timestamp 1712256841
transform 1 0 3304 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_261
timestamp 1712256841
transform 1 0 2344 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_262
timestamp 1712256841
transform 1 0 2008 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_263
timestamp 1712256841
transform 1 0 2184 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_264
timestamp 1712256841
transform 1 0 2400 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_265
timestamp 1712256841
transform 1 0 2488 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_266
timestamp 1712256841
transform 1 0 2600 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_267
timestamp 1712256841
transform 1 0 2776 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_268
timestamp 1712256841
transform 1 0 1200 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_269
timestamp 1712256841
transform 1 0 792 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_270
timestamp 1712256841
transform 1 0 2856 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_271
timestamp 1712256841
transform 1 0 704 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_272
timestamp 1712256841
transform 1 0 608 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_273
timestamp 1712256841
transform 1 0 512 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_274
timestamp 1712256841
transform 1 0 424 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_275
timestamp 1712256841
transform 1 0 360 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_276
timestamp 1712256841
transform 1 0 288 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_277
timestamp 1712256841
transform 1 0 224 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_278
timestamp 1712256841
transform 1 0 80 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_279
timestamp 1712256841
transform 1 0 152 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_280
timestamp 1712256841
transform 1 0 856 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_281
timestamp 1712256841
transform 1 0 2816 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_282
timestamp 1712256841
transform 1 0 1032 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_283
timestamp 1712256841
transform 1 0 1248 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_284
timestamp 1712256841
transform 1 0 1400 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_285
timestamp 1712256841
transform 1 0 1560 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_286
timestamp 1712256841
transform 1 0 1608 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_287
timestamp 1712256841
transform 1 0 1688 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_288
timestamp 1712256841
transform 1 0 1784 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_289
timestamp 1712256841
transform 1 0 1880 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_290
timestamp 1712256841
transform 1 0 2088 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_291
timestamp 1712256841
transform 1 0 2272 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_292
timestamp 1712256841
transform 1 0 2688 0 -1 2570
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1712256841
transform 1 0 2160 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1712256841
transform 1 0 2152 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1712256841
transform 1 0 3336 0 1 1970
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1712256841
transform 1 0 3120 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1712256841
transform 1 0 2640 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1712256841
transform 1 0 2592 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1712256841
transform 1 0 3168 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1712256841
transform 1 0 3104 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1712256841
transform 1 0 1760 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1712256841
transform 1 0 2944 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1712256841
transform 1 0 3128 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1712256841
transform 1 0 3192 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1712256841
transform 1 0 3240 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1712256841
transform 1 0 2360 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1712256841
transform 1 0 2184 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1712256841
transform 1 0 2336 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1712256841
transform 1 0 1976 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1712256841
transform 1 0 1856 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1712256841
transform 1 0 1952 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1712256841
transform 1 0 3160 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1712256841
transform 1 0 2624 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_21
timestamp 1712256841
transform 1 0 2792 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_22
timestamp 1712256841
transform 1 0 2976 0 1 2770
box -5 -3 28 105
use BUFX2  BUFX2_23
timestamp 1712256841
transform 1 0 3136 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1712256841
transform 1 0 3056 0 -1 2970
box -5 -3 28 105
use BUFX2  BUFX2_25
timestamp 1712256841
transform 1 0 2504 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_26
timestamp 1712256841
transform 1 0 2600 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_27
timestamp 1712256841
transform 1 0 2448 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_28
timestamp 1712256841
transform 1 0 2528 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_29
timestamp 1712256841
transform 1 0 2408 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_30
timestamp 1712256841
transform 1 0 2480 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_31
timestamp 1712256841
transform 1 0 1648 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_32
timestamp 1712256841
transform 1 0 3176 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_33
timestamp 1712256841
transform 1 0 1616 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_34
timestamp 1712256841
transform 1 0 3072 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_35
timestamp 1712256841
transform 1 0 2632 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_36
timestamp 1712256841
transform 1 0 1736 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_37
timestamp 1712256841
transform 1 0 1904 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_38
timestamp 1712256841
transform 1 0 2864 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_39
timestamp 1712256841
transform 1 0 1728 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_40
timestamp 1712256841
transform 1 0 1512 0 -1 2970
box -5 -3 28 105
use BUFX2  BUFX2_41
timestamp 1712256841
transform 1 0 1464 0 -1 2970
box -5 -3 28 105
use BUFX2  BUFX2_42
timestamp 1712256841
transform 1 0 1696 0 1 1770
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1712256841
transform 1 0 3336 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1712256841
transform 1 0 3336 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1712256841
transform 1 0 3120 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1712256841
transform 1 0 3120 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1712256841
transform 1 0 2848 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1712256841
transform 1 0 2976 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1712256841
transform 1 0 3088 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1712256841
transform 1 0 3216 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1712256841
transform 1 0 3328 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1712256841
transform 1 0 2720 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1712256841
transform 1 0 2680 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1712256841
transform 1 0 2992 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1712256841
transform 1 0 3040 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1712256841
transform 1 0 3024 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1712256841
transform 1 0 3328 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1712256841
transform 1 0 3224 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1712256841
transform 1 0 3112 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1712256841
transform 1 0 2920 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1712256841
transform 1 0 2800 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1712256841
transform 1 0 3168 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1712256841
transform 1 0 3336 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1712256841
transform 1 0 1192 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1712256841
transform 1 0 880 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1712256841
transform 1 0 656 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1712256841
transform 1 0 544 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1712256841
transform 1 0 432 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1712256841
transform 1 0 320 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1712256841
transform 1 0 288 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1712256841
transform 1 0 208 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1712256841
transform 1 0 88 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1712256841
transform 1 0 80 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1712256841
transform 1 0 128 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1712256841
transform 1 0 768 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1712256841
transform 1 0 928 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1712256841
transform 1 0 1088 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1712256841
transform 1 0 1304 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1712256841
transform 1 0 1456 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1712256841
transform 1 0 1472 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1712256841
transform 1 0 1584 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1712256841
transform 1 0 1696 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1712256841
transform 1 0 1800 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1712256841
transform 1 0 1992 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1712256841
transform 1 0 2184 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1712256841
transform 1 0 2280 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1712256841
transform 1 0 1896 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1712256841
transform 1 0 2088 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1712256841
transform 1 0 2376 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1712256841
transform 1 0 2472 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1712256841
transform 1 0 2568 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1712256841
transform 1 0 2760 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1712256841
transform 1 0 2952 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1712256841
transform 1 0 2856 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1712256841
transform 1 0 2664 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1712256841
transform 1 0 2936 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1712256841
transform 1 0 928 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1712256841
transform 1 0 728 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1712256841
transform 1 0 360 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1712256841
transform 1 0 520 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1712256841
transform 1 0 408 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1712256841
transform 1 0 296 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1712256841
transform 1 0 344 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1712256841
transform 1 0 240 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1712256841
transform 1 0 160 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1712256841
transform 1 0 80 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1712256841
transform 1 0 80 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1712256841
transform 1 0 1048 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1712256841
transform 1 0 1104 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1712256841
transform 1 0 1304 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1712256841
transform 1 0 1280 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1712256841
transform 1 0 1360 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1712256841
transform 1 0 1520 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1712256841
transform 1 0 1576 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1712256841
transform 1 0 1792 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1712256841
transform 1 0 1664 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1712256841
transform 1 0 1936 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1712256841
transform 1 0 2104 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1712256841
transform 1 0 2272 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1712256841
transform 1 0 2048 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1712256841
transform 1 0 2464 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1712256841
transform 1 0 2704 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1712256841
transform 1 0 2576 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1712256841
transform 1 0 2584 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1712256841
transform 1 0 2808 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1712256841
transform 1 0 3136 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1712256841
transform 1 0 2912 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1712256841
transform 1 0 2704 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1712256841
transform 1 0 3104 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1712256841
transform 1 0 3040 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1712256841
transform 1 0 1104 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1712256841
transform 1 0 776 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1712256841
transform 1 0 664 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1712256841
transform 1 0 560 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1712256841
transform 1 0 424 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1712256841
transform 1 0 408 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1712256841
transform 1 0 288 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1712256841
transform 1 0 296 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1712256841
transform 1 0 184 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1712256841
transform 1 0 72 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1712256841
transform 1 0 128 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1712256841
transform 1 0 888 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1712256841
transform 1 0 992 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1712256841
transform 1 0 1216 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1712256841
transform 1 0 1320 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1712256841
transform 1 0 1432 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1712256841
transform 1 0 1536 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1712256841
transform 1 0 1648 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1712256841
transform 1 0 1744 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1712256841
transform 1 0 1848 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1712256841
transform 1 0 2056 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1712256841
transform 1 0 2104 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1712256841
transform 1 0 2208 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1712256841
transform 1 0 1952 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1712256841
transform 1 0 2256 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1712256841
transform 1 0 2408 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1712256841
transform 1 0 2640 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1712256841
transform 1 0 2528 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1712256841
transform 1 0 2760 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1712256841
transform 1 0 2888 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1712256841
transform 1 0 2880 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1712256841
transform 1 0 2680 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1712256841
transform 1 0 3240 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1712256841
transform 1 0 3328 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1712256841
transform 1 0 3248 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1712256841
transform 1 0 3336 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1712256841
transform 1 0 3256 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1712256841
transform 1 0 3048 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1712256841
transform 1 0 3144 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1712256841
transform 1 0 3328 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_128
timestamp 1712256841
transform 1 0 3328 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1712256841
transform 1 0 3328 0 -1 2570
box -8 -3 104 105
use FILL  FILL_0
timestamp 1712256841
transform 1 0 3424 0 1 3170
box -8 -3 16 105
use FILL  FILL_1
timestamp 1712256841
transform 1 0 3416 0 1 3170
box -8 -3 16 105
use FILL  FILL_2
timestamp 1712256841
transform 1 0 3360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3
timestamp 1712256841
transform 1 0 3352 0 1 3170
box -8 -3 16 105
use FILL  FILL_4
timestamp 1712256841
transform 1 0 3344 0 1 3170
box -8 -3 16 105
use FILL  FILL_5
timestamp 1712256841
transform 1 0 3240 0 1 3170
box -8 -3 16 105
use FILL  FILL_6
timestamp 1712256841
transform 1 0 3232 0 1 3170
box -8 -3 16 105
use FILL  FILL_7
timestamp 1712256841
transform 1 0 3128 0 1 3170
box -8 -3 16 105
use FILL  FILL_8
timestamp 1712256841
transform 1 0 3120 0 1 3170
box -8 -3 16 105
use FILL  FILL_9
timestamp 1712256841
transform 1 0 3096 0 1 3170
box -8 -3 16 105
use FILL  FILL_10
timestamp 1712256841
transform 1 0 3016 0 1 3170
box -8 -3 16 105
use FILL  FILL_11
timestamp 1712256841
transform 1 0 3008 0 1 3170
box -8 -3 16 105
use FILL  FILL_12
timestamp 1712256841
transform 1 0 3000 0 1 3170
box -8 -3 16 105
use FILL  FILL_13
timestamp 1712256841
transform 1 0 2992 0 1 3170
box -8 -3 16 105
use FILL  FILL_14
timestamp 1712256841
transform 1 0 2936 0 1 3170
box -8 -3 16 105
use FILL  FILL_15
timestamp 1712256841
transform 1 0 2928 0 1 3170
box -8 -3 16 105
use FILL  FILL_16
timestamp 1712256841
transform 1 0 2920 0 1 3170
box -8 -3 16 105
use FILL  FILL_17
timestamp 1712256841
transform 1 0 2912 0 1 3170
box -8 -3 16 105
use FILL  FILL_18
timestamp 1712256841
transform 1 0 2840 0 1 3170
box -8 -3 16 105
use FILL  FILL_19
timestamp 1712256841
transform 1 0 2832 0 1 3170
box -8 -3 16 105
use FILL  FILL_20
timestamp 1712256841
transform 1 0 2824 0 1 3170
box -8 -3 16 105
use FILL  FILL_21
timestamp 1712256841
transform 1 0 2816 0 1 3170
box -8 -3 16 105
use FILL  FILL_22
timestamp 1712256841
transform 1 0 2752 0 1 3170
box -8 -3 16 105
use FILL  FILL_23
timestamp 1712256841
transform 1 0 2744 0 1 3170
box -8 -3 16 105
use FILL  FILL_24
timestamp 1712256841
transform 1 0 2688 0 1 3170
box -8 -3 16 105
use FILL  FILL_25
timestamp 1712256841
transform 1 0 2680 0 1 3170
box -8 -3 16 105
use FILL  FILL_26
timestamp 1712256841
transform 1 0 2672 0 1 3170
box -8 -3 16 105
use FILL  FILL_27
timestamp 1712256841
transform 1 0 2568 0 1 3170
box -8 -3 16 105
use FILL  FILL_28
timestamp 1712256841
transform 1 0 2560 0 1 3170
box -8 -3 16 105
use FILL  FILL_29
timestamp 1712256841
transform 1 0 2496 0 1 3170
box -8 -3 16 105
use FILL  FILL_30
timestamp 1712256841
transform 1 0 2488 0 1 3170
box -8 -3 16 105
use FILL  FILL_31
timestamp 1712256841
transform 1 0 2480 0 1 3170
box -8 -3 16 105
use FILL  FILL_32
timestamp 1712256841
transform 1 0 2432 0 1 3170
box -8 -3 16 105
use FILL  FILL_33
timestamp 1712256841
transform 1 0 2392 0 1 3170
box -8 -3 16 105
use FILL  FILL_34
timestamp 1712256841
transform 1 0 2384 0 1 3170
box -8 -3 16 105
use FILL  FILL_35
timestamp 1712256841
transform 1 0 2376 0 1 3170
box -8 -3 16 105
use FILL  FILL_36
timestamp 1712256841
transform 1 0 2312 0 1 3170
box -8 -3 16 105
use FILL  FILL_37
timestamp 1712256841
transform 1 0 2304 0 1 3170
box -8 -3 16 105
use FILL  FILL_38
timestamp 1712256841
transform 1 0 2296 0 1 3170
box -8 -3 16 105
use FILL  FILL_39
timestamp 1712256841
transform 1 0 2256 0 1 3170
box -8 -3 16 105
use FILL  FILL_40
timestamp 1712256841
transform 1 0 2248 0 1 3170
box -8 -3 16 105
use FILL  FILL_41
timestamp 1712256841
transform 1 0 2240 0 1 3170
box -8 -3 16 105
use FILL  FILL_42
timestamp 1712256841
transform 1 0 2232 0 1 3170
box -8 -3 16 105
use FILL  FILL_43
timestamp 1712256841
transform 1 0 2144 0 1 3170
box -8 -3 16 105
use FILL  FILL_44
timestamp 1712256841
transform 1 0 2136 0 1 3170
box -8 -3 16 105
use FILL  FILL_45
timestamp 1712256841
transform 1 0 2128 0 1 3170
box -8 -3 16 105
use FILL  FILL_46
timestamp 1712256841
transform 1 0 2040 0 1 3170
box -8 -3 16 105
use FILL  FILL_47
timestamp 1712256841
transform 1 0 2032 0 1 3170
box -8 -3 16 105
use FILL  FILL_48
timestamp 1712256841
transform 1 0 2024 0 1 3170
box -8 -3 16 105
use FILL  FILL_49
timestamp 1712256841
transform 1 0 1952 0 1 3170
box -8 -3 16 105
use FILL  FILL_50
timestamp 1712256841
transform 1 0 1944 0 1 3170
box -8 -3 16 105
use FILL  FILL_51
timestamp 1712256841
transform 1 0 1880 0 1 3170
box -8 -3 16 105
use FILL  FILL_52
timestamp 1712256841
transform 1 0 1872 0 1 3170
box -8 -3 16 105
use FILL  FILL_53
timestamp 1712256841
transform 1 0 1808 0 1 3170
box -8 -3 16 105
use FILL  FILL_54
timestamp 1712256841
transform 1 0 1800 0 1 3170
box -8 -3 16 105
use FILL  FILL_55
timestamp 1712256841
transform 1 0 1792 0 1 3170
box -8 -3 16 105
use FILL  FILL_56
timestamp 1712256841
transform 1 0 1728 0 1 3170
box -8 -3 16 105
use FILL  FILL_57
timestamp 1712256841
transform 1 0 1720 0 1 3170
box -8 -3 16 105
use FILL  FILL_58
timestamp 1712256841
transform 1 0 1712 0 1 3170
box -8 -3 16 105
use FILL  FILL_59
timestamp 1712256841
transform 1 0 1704 0 1 3170
box -8 -3 16 105
use FILL  FILL_60
timestamp 1712256841
transform 1 0 1680 0 1 3170
box -8 -3 16 105
use FILL  FILL_61
timestamp 1712256841
transform 1 0 1624 0 1 3170
box -8 -3 16 105
use FILL  FILL_62
timestamp 1712256841
transform 1 0 1616 0 1 3170
box -8 -3 16 105
use FILL  FILL_63
timestamp 1712256841
transform 1 0 1608 0 1 3170
box -8 -3 16 105
use FILL  FILL_64
timestamp 1712256841
transform 1 0 1600 0 1 3170
box -8 -3 16 105
use FILL  FILL_65
timestamp 1712256841
transform 1 0 1552 0 1 3170
box -8 -3 16 105
use FILL  FILL_66
timestamp 1712256841
transform 1 0 1512 0 1 3170
box -8 -3 16 105
use FILL  FILL_67
timestamp 1712256841
transform 1 0 1504 0 1 3170
box -8 -3 16 105
use FILL  FILL_68
timestamp 1712256841
transform 1 0 1464 0 1 3170
box -8 -3 16 105
use FILL  FILL_69
timestamp 1712256841
transform 1 0 1456 0 1 3170
box -8 -3 16 105
use FILL  FILL_70
timestamp 1712256841
transform 1 0 1448 0 1 3170
box -8 -3 16 105
use FILL  FILL_71
timestamp 1712256841
transform 1 0 1440 0 1 3170
box -8 -3 16 105
use FILL  FILL_72
timestamp 1712256841
transform 1 0 1376 0 1 3170
box -8 -3 16 105
use FILL  FILL_73
timestamp 1712256841
transform 1 0 1368 0 1 3170
box -8 -3 16 105
use FILL  FILL_74
timestamp 1712256841
transform 1 0 1360 0 1 3170
box -8 -3 16 105
use FILL  FILL_75
timestamp 1712256841
transform 1 0 1352 0 1 3170
box -8 -3 16 105
use FILL  FILL_76
timestamp 1712256841
transform 1 0 1344 0 1 3170
box -8 -3 16 105
use FILL  FILL_77
timestamp 1712256841
transform 1 0 1272 0 1 3170
box -8 -3 16 105
use FILL  FILL_78
timestamp 1712256841
transform 1 0 1264 0 1 3170
box -8 -3 16 105
use FILL  FILL_79
timestamp 1712256841
transform 1 0 1256 0 1 3170
box -8 -3 16 105
use FILL  FILL_80
timestamp 1712256841
transform 1 0 1184 0 1 3170
box -8 -3 16 105
use FILL  FILL_81
timestamp 1712256841
transform 1 0 1176 0 1 3170
box -8 -3 16 105
use FILL  FILL_82
timestamp 1712256841
transform 1 0 1168 0 1 3170
box -8 -3 16 105
use FILL  FILL_83
timestamp 1712256841
transform 1 0 1160 0 1 3170
box -8 -3 16 105
use FILL  FILL_84
timestamp 1712256841
transform 1 0 1104 0 1 3170
box -8 -3 16 105
use FILL  FILL_85
timestamp 1712256841
transform 1 0 1096 0 1 3170
box -8 -3 16 105
use FILL  FILL_86
timestamp 1712256841
transform 1 0 1056 0 1 3170
box -8 -3 16 105
use FILL  FILL_87
timestamp 1712256841
transform 1 0 1048 0 1 3170
box -8 -3 16 105
use FILL  FILL_88
timestamp 1712256841
transform 1 0 1024 0 1 3170
box -8 -3 16 105
use FILL  FILL_89
timestamp 1712256841
transform 1 0 1016 0 1 3170
box -8 -3 16 105
use FILL  FILL_90
timestamp 1712256841
transform 1 0 952 0 1 3170
box -8 -3 16 105
use FILL  FILL_91
timestamp 1712256841
transform 1 0 944 0 1 3170
box -8 -3 16 105
use FILL  FILL_92
timestamp 1712256841
transform 1 0 920 0 1 3170
box -8 -3 16 105
use FILL  FILL_93
timestamp 1712256841
transform 1 0 912 0 1 3170
box -8 -3 16 105
use FILL  FILL_94
timestamp 1712256841
transform 1 0 840 0 1 3170
box -8 -3 16 105
use FILL  FILL_95
timestamp 1712256841
transform 1 0 832 0 1 3170
box -8 -3 16 105
use FILL  FILL_96
timestamp 1712256841
transform 1 0 824 0 1 3170
box -8 -3 16 105
use FILL  FILL_97
timestamp 1712256841
transform 1 0 776 0 1 3170
box -8 -3 16 105
use FILL  FILL_98
timestamp 1712256841
transform 1 0 744 0 1 3170
box -8 -3 16 105
use FILL  FILL_99
timestamp 1712256841
transform 1 0 720 0 1 3170
box -8 -3 16 105
use FILL  FILL_100
timestamp 1712256841
transform 1 0 712 0 1 3170
box -8 -3 16 105
use FILL  FILL_101
timestamp 1712256841
transform 1 0 704 0 1 3170
box -8 -3 16 105
use FILL  FILL_102
timestamp 1712256841
transform 1 0 656 0 1 3170
box -8 -3 16 105
use FILL  FILL_103
timestamp 1712256841
transform 1 0 608 0 1 3170
box -8 -3 16 105
use FILL  FILL_104
timestamp 1712256841
transform 1 0 600 0 1 3170
box -8 -3 16 105
use FILL  FILL_105
timestamp 1712256841
transform 1 0 592 0 1 3170
box -8 -3 16 105
use FILL  FILL_106
timestamp 1712256841
transform 1 0 520 0 1 3170
box -8 -3 16 105
use FILL  FILL_107
timestamp 1712256841
transform 1 0 512 0 1 3170
box -8 -3 16 105
use FILL  FILL_108
timestamp 1712256841
transform 1 0 504 0 1 3170
box -8 -3 16 105
use FILL  FILL_109
timestamp 1712256841
transform 1 0 400 0 1 3170
box -8 -3 16 105
use FILL  FILL_110
timestamp 1712256841
transform 1 0 392 0 1 3170
box -8 -3 16 105
use FILL  FILL_111
timestamp 1712256841
transform 1 0 288 0 1 3170
box -8 -3 16 105
use FILL  FILL_112
timestamp 1712256841
transform 1 0 280 0 1 3170
box -8 -3 16 105
use FILL  FILL_113
timestamp 1712256841
transform 1 0 256 0 1 3170
box -8 -3 16 105
use FILL  FILL_114
timestamp 1712256841
transform 1 0 152 0 1 3170
box -8 -3 16 105
use FILL  FILL_115
timestamp 1712256841
transform 1 0 144 0 1 3170
box -8 -3 16 105
use FILL  FILL_116
timestamp 1712256841
transform 1 0 136 0 1 3170
box -8 -3 16 105
use FILL  FILL_117
timestamp 1712256841
transform 1 0 128 0 1 3170
box -8 -3 16 105
use FILL  FILL_118
timestamp 1712256841
transform 1 0 120 0 1 3170
box -8 -3 16 105
use FILL  FILL_119
timestamp 1712256841
transform 1 0 112 0 1 3170
box -8 -3 16 105
use FILL  FILL_120
timestamp 1712256841
transform 1 0 104 0 1 3170
box -8 -3 16 105
use FILL  FILL_121
timestamp 1712256841
transform 1 0 96 0 1 3170
box -8 -3 16 105
use FILL  FILL_122
timestamp 1712256841
transform 1 0 88 0 1 3170
box -8 -3 16 105
use FILL  FILL_123
timestamp 1712256841
transform 1 0 80 0 1 3170
box -8 -3 16 105
use FILL  FILL_124
timestamp 1712256841
transform 1 0 72 0 1 3170
box -8 -3 16 105
use FILL  FILL_125
timestamp 1712256841
transform 1 0 3424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_126
timestamp 1712256841
transform 1 0 3416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_127
timestamp 1712256841
transform 1 0 3408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_128
timestamp 1712256841
transform 1 0 3352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_129
timestamp 1712256841
transform 1 0 3320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_130
timestamp 1712256841
transform 1 0 3312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_131
timestamp 1712256841
transform 1 0 3304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_132
timestamp 1712256841
transform 1 0 3296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_133
timestamp 1712256841
transform 1 0 3232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_134
timestamp 1712256841
transform 1 0 3224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_135
timestamp 1712256841
transform 1 0 3216 0 -1 3170
box -8 -3 16 105
use FILL  FILL_136
timestamp 1712256841
transform 1 0 3168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_137
timestamp 1712256841
transform 1 0 3160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_138
timestamp 1712256841
transform 1 0 3152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_139
timestamp 1712256841
transform 1 0 3112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_140
timestamp 1712256841
transform 1 0 3104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_141
timestamp 1712256841
transform 1 0 3096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_142
timestamp 1712256841
transform 1 0 3064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_143
timestamp 1712256841
transform 1 0 3032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_144
timestamp 1712256841
transform 1 0 3024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_145
timestamp 1712256841
transform 1 0 3016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_146
timestamp 1712256841
transform 1 0 3008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_147
timestamp 1712256841
transform 1 0 3000 0 -1 3170
box -8 -3 16 105
use FILL  FILL_148
timestamp 1712256841
transform 1 0 2936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_149
timestamp 1712256841
transform 1 0 2928 0 -1 3170
box -8 -3 16 105
use FILL  FILL_150
timestamp 1712256841
transform 1 0 2920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_151
timestamp 1712256841
transform 1 0 2912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_152
timestamp 1712256841
transform 1 0 2840 0 -1 3170
box -8 -3 16 105
use FILL  FILL_153
timestamp 1712256841
transform 1 0 2832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_154
timestamp 1712256841
transform 1 0 2824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_155
timestamp 1712256841
transform 1 0 2816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_156
timestamp 1712256841
transform 1 0 2808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_157
timestamp 1712256841
transform 1 0 2784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_158
timestamp 1712256841
transform 1 0 2736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_159
timestamp 1712256841
transform 1 0 2728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_160
timestamp 1712256841
transform 1 0 2680 0 -1 3170
box -8 -3 16 105
use FILL  FILL_161
timestamp 1712256841
transform 1 0 2672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_162
timestamp 1712256841
transform 1 0 2664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_163
timestamp 1712256841
transform 1 0 2656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_164
timestamp 1712256841
transform 1 0 2584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_165
timestamp 1712256841
transform 1 0 2576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_166
timestamp 1712256841
transform 1 0 2568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_167
timestamp 1712256841
transform 1 0 2560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_168
timestamp 1712256841
transform 1 0 2504 0 -1 3170
box -8 -3 16 105
use FILL  FILL_169
timestamp 1712256841
transform 1 0 2496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_170
timestamp 1712256841
transform 1 0 2488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_171
timestamp 1712256841
transform 1 0 2424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_172
timestamp 1712256841
transform 1 0 2416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_173
timestamp 1712256841
transform 1 0 2408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_174
timestamp 1712256841
transform 1 0 2352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_175
timestamp 1712256841
transform 1 0 2344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_176
timestamp 1712256841
transform 1 0 2296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_177
timestamp 1712256841
transform 1 0 2288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_178
timestamp 1712256841
transform 1 0 2240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_179
timestamp 1712256841
transform 1 0 2232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_180
timestamp 1712256841
transform 1 0 2192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_181
timestamp 1712256841
transform 1 0 2144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_182
timestamp 1712256841
transform 1 0 2136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_183
timestamp 1712256841
transform 1 0 2128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_184
timestamp 1712256841
transform 1 0 2088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_185
timestamp 1712256841
transform 1 0 2080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_186
timestamp 1712256841
transform 1 0 2024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_187
timestamp 1712256841
transform 1 0 1984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_188
timestamp 1712256841
transform 1 0 1976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_189
timestamp 1712256841
transform 1 0 1968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_190
timestamp 1712256841
transform 1 0 1904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_191
timestamp 1712256841
transform 1 0 1896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_192
timestamp 1712256841
transform 1 0 1888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_193
timestamp 1712256841
transform 1 0 1880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_194
timestamp 1712256841
transform 1 0 1840 0 -1 3170
box -8 -3 16 105
use FILL  FILL_195
timestamp 1712256841
transform 1 0 1832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_196
timestamp 1712256841
transform 1 0 1792 0 -1 3170
box -8 -3 16 105
use FILL  FILL_197
timestamp 1712256841
transform 1 0 1784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_198
timestamp 1712256841
transform 1 0 1744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_199
timestamp 1712256841
transform 1 0 1736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_200
timestamp 1712256841
transform 1 0 1728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_201
timestamp 1712256841
transform 1 0 1680 0 -1 3170
box -8 -3 16 105
use FILL  FILL_202
timestamp 1712256841
transform 1 0 1672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_203
timestamp 1712256841
transform 1 0 1664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_204
timestamp 1712256841
transform 1 0 1632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_205
timestamp 1712256841
transform 1 0 1584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_206
timestamp 1712256841
transform 1 0 1576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_207
timestamp 1712256841
transform 1 0 1568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_208
timestamp 1712256841
transform 1 0 1560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_209
timestamp 1712256841
transform 1 0 1512 0 -1 3170
box -8 -3 16 105
use FILL  FILL_210
timestamp 1712256841
transform 1 0 1472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_211
timestamp 1712256841
transform 1 0 1464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_212
timestamp 1712256841
transform 1 0 1456 0 -1 3170
box -8 -3 16 105
use FILL  FILL_213
timestamp 1712256841
transform 1 0 1448 0 -1 3170
box -8 -3 16 105
use FILL  FILL_214
timestamp 1712256841
transform 1 0 1440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_215
timestamp 1712256841
transform 1 0 1368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_216
timestamp 1712256841
transform 1 0 1360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_217
timestamp 1712256841
transform 1 0 1352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_218
timestamp 1712256841
transform 1 0 1344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_219
timestamp 1712256841
transform 1 0 1296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_220
timestamp 1712256841
transform 1 0 1288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_221
timestamp 1712256841
transform 1 0 1280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_222
timestamp 1712256841
transform 1 0 1216 0 -1 3170
box -8 -3 16 105
use FILL  FILL_223
timestamp 1712256841
transform 1 0 1208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_224
timestamp 1712256841
transform 1 0 1200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_225
timestamp 1712256841
transform 1 0 1192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_226
timestamp 1712256841
transform 1 0 1184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_227
timestamp 1712256841
transform 1 0 1104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_228
timestamp 1712256841
transform 1 0 1096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_229
timestamp 1712256841
transform 1 0 1088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_230
timestamp 1712256841
transform 1 0 1080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_231
timestamp 1712256841
transform 1 0 1032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_232
timestamp 1712256841
transform 1 0 1024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_233
timestamp 1712256841
transform 1 0 1016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_234
timestamp 1712256841
transform 1 0 960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_235
timestamp 1712256841
transform 1 0 952 0 -1 3170
box -8 -3 16 105
use FILL  FILL_236
timestamp 1712256841
transform 1 0 944 0 -1 3170
box -8 -3 16 105
use FILL  FILL_237
timestamp 1712256841
transform 1 0 904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_238
timestamp 1712256841
transform 1 0 896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_239
timestamp 1712256841
transform 1 0 832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_240
timestamp 1712256841
transform 1 0 824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_241
timestamp 1712256841
transform 1 0 816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_242
timestamp 1712256841
transform 1 0 808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_243
timestamp 1712256841
transform 1 0 800 0 -1 3170
box -8 -3 16 105
use FILL  FILL_244
timestamp 1712256841
transform 1 0 792 0 -1 3170
box -8 -3 16 105
use FILL  FILL_245
timestamp 1712256841
transform 1 0 696 0 -1 3170
box -8 -3 16 105
use FILL  FILL_246
timestamp 1712256841
transform 1 0 688 0 -1 3170
box -8 -3 16 105
use FILL  FILL_247
timestamp 1712256841
transform 1 0 680 0 -1 3170
box -8 -3 16 105
use FILL  FILL_248
timestamp 1712256841
transform 1 0 672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_249
timestamp 1712256841
transform 1 0 664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_250
timestamp 1712256841
transform 1 0 600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_251
timestamp 1712256841
transform 1 0 592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_252
timestamp 1712256841
transform 1 0 584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_253
timestamp 1712256841
transform 1 0 496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_254
timestamp 1712256841
transform 1 0 488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_255
timestamp 1712256841
transform 1 0 480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_256
timestamp 1712256841
transform 1 0 472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_257
timestamp 1712256841
transform 1 0 464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_258
timestamp 1712256841
transform 1 0 408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_259
timestamp 1712256841
transform 1 0 400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_260
timestamp 1712256841
transform 1 0 392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_261
timestamp 1712256841
transform 1 0 384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_262
timestamp 1712256841
transform 1 0 376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_263
timestamp 1712256841
transform 1 0 320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_264
timestamp 1712256841
transform 1 0 312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_265
timestamp 1712256841
transform 1 0 272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_266
timestamp 1712256841
transform 1 0 264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_267
timestamp 1712256841
transform 1 0 256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_268
timestamp 1712256841
transform 1 0 200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_269
timestamp 1712256841
transform 1 0 192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_270
timestamp 1712256841
transform 1 0 184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_271
timestamp 1712256841
transform 1 0 176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_272
timestamp 1712256841
transform 1 0 72 0 -1 3170
box -8 -3 16 105
use FILL  FILL_273
timestamp 1712256841
transform 1 0 3424 0 1 2970
box -8 -3 16 105
use FILL  FILL_274
timestamp 1712256841
transform 1 0 3320 0 1 2970
box -8 -3 16 105
use FILL  FILL_275
timestamp 1712256841
transform 1 0 3312 0 1 2970
box -8 -3 16 105
use FILL  FILL_276
timestamp 1712256841
transform 1 0 3240 0 1 2970
box -8 -3 16 105
use FILL  FILL_277
timestamp 1712256841
transform 1 0 3216 0 1 2970
box -8 -3 16 105
use FILL  FILL_278
timestamp 1712256841
transform 1 0 3208 0 1 2970
box -8 -3 16 105
use FILL  FILL_279
timestamp 1712256841
transform 1 0 3200 0 1 2970
box -8 -3 16 105
use FILL  FILL_280
timestamp 1712256841
transform 1 0 3096 0 1 2970
box -8 -3 16 105
use FILL  FILL_281
timestamp 1712256841
transform 1 0 3088 0 1 2970
box -8 -3 16 105
use FILL  FILL_282
timestamp 1712256841
transform 1 0 3080 0 1 2970
box -8 -3 16 105
use FILL  FILL_283
timestamp 1712256841
transform 1 0 3072 0 1 2970
box -8 -3 16 105
use FILL  FILL_284
timestamp 1712256841
transform 1 0 3008 0 1 2970
box -8 -3 16 105
use FILL  FILL_285
timestamp 1712256841
transform 1 0 3000 0 1 2970
box -8 -3 16 105
use FILL  FILL_286
timestamp 1712256841
transform 1 0 2992 0 1 2970
box -8 -3 16 105
use FILL  FILL_287
timestamp 1712256841
transform 1 0 2984 0 1 2970
box -8 -3 16 105
use FILL  FILL_288
timestamp 1712256841
transform 1 0 2976 0 1 2970
box -8 -3 16 105
use FILL  FILL_289
timestamp 1712256841
transform 1 0 2928 0 1 2970
box -8 -3 16 105
use FILL  FILL_290
timestamp 1712256841
transform 1 0 2920 0 1 2970
box -8 -3 16 105
use FILL  FILL_291
timestamp 1712256841
transform 1 0 2912 0 1 2970
box -8 -3 16 105
use FILL  FILL_292
timestamp 1712256841
transform 1 0 2904 0 1 2970
box -8 -3 16 105
use FILL  FILL_293
timestamp 1712256841
transform 1 0 2896 0 1 2970
box -8 -3 16 105
use FILL  FILL_294
timestamp 1712256841
transform 1 0 2824 0 1 2970
box -8 -3 16 105
use FILL  FILL_295
timestamp 1712256841
transform 1 0 2816 0 1 2970
box -8 -3 16 105
use FILL  FILL_296
timestamp 1712256841
transform 1 0 2808 0 1 2970
box -8 -3 16 105
use FILL  FILL_297
timestamp 1712256841
transform 1 0 2800 0 1 2970
box -8 -3 16 105
use FILL  FILL_298
timestamp 1712256841
transform 1 0 2696 0 1 2970
box -8 -3 16 105
use FILL  FILL_299
timestamp 1712256841
transform 1 0 2688 0 1 2970
box -8 -3 16 105
use FILL  FILL_300
timestamp 1712256841
transform 1 0 2680 0 1 2970
box -8 -3 16 105
use FILL  FILL_301
timestamp 1712256841
transform 1 0 2672 0 1 2970
box -8 -3 16 105
use FILL  FILL_302
timestamp 1712256841
transform 1 0 2664 0 1 2970
box -8 -3 16 105
use FILL  FILL_303
timestamp 1712256841
transform 1 0 2608 0 1 2970
box -8 -3 16 105
use FILL  FILL_304
timestamp 1712256841
transform 1 0 2600 0 1 2970
box -8 -3 16 105
use FILL  FILL_305
timestamp 1712256841
transform 1 0 2592 0 1 2970
box -8 -3 16 105
use FILL  FILL_306
timestamp 1712256841
transform 1 0 2584 0 1 2970
box -8 -3 16 105
use FILL  FILL_307
timestamp 1712256841
transform 1 0 2576 0 1 2970
box -8 -3 16 105
use FILL  FILL_308
timestamp 1712256841
transform 1 0 2504 0 1 2970
box -8 -3 16 105
use FILL  FILL_309
timestamp 1712256841
transform 1 0 2496 0 1 2970
box -8 -3 16 105
use FILL  FILL_310
timestamp 1712256841
transform 1 0 2488 0 1 2970
box -8 -3 16 105
use FILL  FILL_311
timestamp 1712256841
transform 1 0 2480 0 1 2970
box -8 -3 16 105
use FILL  FILL_312
timestamp 1712256841
transform 1 0 2456 0 1 2970
box -8 -3 16 105
use FILL  FILL_313
timestamp 1712256841
transform 1 0 2400 0 1 2970
box -8 -3 16 105
use FILL  FILL_314
timestamp 1712256841
transform 1 0 2392 0 1 2970
box -8 -3 16 105
use FILL  FILL_315
timestamp 1712256841
transform 1 0 2384 0 1 2970
box -8 -3 16 105
use FILL  FILL_316
timestamp 1712256841
transform 1 0 2376 0 1 2970
box -8 -3 16 105
use FILL  FILL_317
timestamp 1712256841
transform 1 0 2368 0 1 2970
box -8 -3 16 105
use FILL  FILL_318
timestamp 1712256841
transform 1 0 2288 0 1 2970
box -8 -3 16 105
use FILL  FILL_319
timestamp 1712256841
transform 1 0 2280 0 1 2970
box -8 -3 16 105
use FILL  FILL_320
timestamp 1712256841
transform 1 0 2272 0 1 2970
box -8 -3 16 105
use FILL  FILL_321
timestamp 1712256841
transform 1 0 2264 0 1 2970
box -8 -3 16 105
use FILL  FILL_322
timestamp 1712256841
transform 1 0 2200 0 1 2970
box -8 -3 16 105
use FILL  FILL_323
timestamp 1712256841
transform 1 0 2192 0 1 2970
box -8 -3 16 105
use FILL  FILL_324
timestamp 1712256841
transform 1 0 2160 0 1 2970
box -8 -3 16 105
use FILL  FILL_325
timestamp 1712256841
transform 1 0 2152 0 1 2970
box -8 -3 16 105
use FILL  FILL_326
timestamp 1712256841
transform 1 0 2112 0 1 2970
box -8 -3 16 105
use FILL  FILL_327
timestamp 1712256841
transform 1 0 2064 0 1 2970
box -8 -3 16 105
use FILL  FILL_328
timestamp 1712256841
transform 1 0 2056 0 1 2970
box -8 -3 16 105
use FILL  FILL_329
timestamp 1712256841
transform 1 0 2048 0 1 2970
box -8 -3 16 105
use FILL  FILL_330
timestamp 1712256841
transform 1 0 1984 0 1 2970
box -8 -3 16 105
use FILL  FILL_331
timestamp 1712256841
transform 1 0 1976 0 1 2970
box -8 -3 16 105
use FILL  FILL_332
timestamp 1712256841
transform 1 0 1968 0 1 2970
box -8 -3 16 105
use FILL  FILL_333
timestamp 1712256841
transform 1 0 1888 0 1 2970
box -8 -3 16 105
use FILL  FILL_334
timestamp 1712256841
transform 1 0 1880 0 1 2970
box -8 -3 16 105
use FILL  FILL_335
timestamp 1712256841
transform 1 0 1872 0 1 2970
box -8 -3 16 105
use FILL  FILL_336
timestamp 1712256841
transform 1 0 1864 0 1 2970
box -8 -3 16 105
use FILL  FILL_337
timestamp 1712256841
transform 1 0 1784 0 1 2970
box -8 -3 16 105
use FILL  FILL_338
timestamp 1712256841
transform 1 0 1776 0 1 2970
box -8 -3 16 105
use FILL  FILL_339
timestamp 1712256841
transform 1 0 1768 0 1 2970
box -8 -3 16 105
use FILL  FILL_340
timestamp 1712256841
transform 1 0 1760 0 1 2970
box -8 -3 16 105
use FILL  FILL_341
timestamp 1712256841
transform 1 0 1680 0 1 2970
box -8 -3 16 105
use FILL  FILL_342
timestamp 1712256841
transform 1 0 1672 0 1 2970
box -8 -3 16 105
use FILL  FILL_343
timestamp 1712256841
transform 1 0 1664 0 1 2970
box -8 -3 16 105
use FILL  FILL_344
timestamp 1712256841
transform 1 0 1576 0 1 2970
box -8 -3 16 105
use FILL  FILL_345
timestamp 1712256841
transform 1 0 1568 0 1 2970
box -8 -3 16 105
use FILL  FILL_346
timestamp 1712256841
transform 1 0 1560 0 1 2970
box -8 -3 16 105
use FILL  FILL_347
timestamp 1712256841
transform 1 0 1552 0 1 2970
box -8 -3 16 105
use FILL  FILL_348
timestamp 1712256841
transform 1 0 1480 0 1 2970
box -8 -3 16 105
use FILL  FILL_349
timestamp 1712256841
transform 1 0 1472 0 1 2970
box -8 -3 16 105
use FILL  FILL_350
timestamp 1712256841
transform 1 0 1424 0 1 2970
box -8 -3 16 105
use FILL  FILL_351
timestamp 1712256841
transform 1 0 1384 0 1 2970
box -8 -3 16 105
use FILL  FILL_352
timestamp 1712256841
transform 1 0 1376 0 1 2970
box -8 -3 16 105
use FILL  FILL_353
timestamp 1712256841
transform 1 0 1368 0 1 2970
box -8 -3 16 105
use FILL  FILL_354
timestamp 1712256841
transform 1 0 1320 0 1 2970
box -8 -3 16 105
use FILL  FILL_355
timestamp 1712256841
transform 1 0 1296 0 1 2970
box -8 -3 16 105
use FILL  FILL_356
timestamp 1712256841
transform 1 0 1288 0 1 2970
box -8 -3 16 105
use FILL  FILL_357
timestamp 1712256841
transform 1 0 1256 0 1 2970
box -8 -3 16 105
use FILL  FILL_358
timestamp 1712256841
transform 1 0 1248 0 1 2970
box -8 -3 16 105
use FILL  FILL_359
timestamp 1712256841
transform 1 0 1240 0 1 2970
box -8 -3 16 105
use FILL  FILL_360
timestamp 1712256841
transform 1 0 1160 0 1 2970
box -8 -3 16 105
use FILL  FILL_361
timestamp 1712256841
transform 1 0 1152 0 1 2970
box -8 -3 16 105
use FILL  FILL_362
timestamp 1712256841
transform 1 0 1144 0 1 2970
box -8 -3 16 105
use FILL  FILL_363
timestamp 1712256841
transform 1 0 1136 0 1 2970
box -8 -3 16 105
use FILL  FILL_364
timestamp 1712256841
transform 1 0 1056 0 1 2970
box -8 -3 16 105
use FILL  FILL_365
timestamp 1712256841
transform 1 0 1048 0 1 2970
box -8 -3 16 105
use FILL  FILL_366
timestamp 1712256841
transform 1 0 1040 0 1 2970
box -8 -3 16 105
use FILL  FILL_367
timestamp 1712256841
transform 1 0 960 0 1 2970
box -8 -3 16 105
use FILL  FILL_368
timestamp 1712256841
transform 1 0 952 0 1 2970
box -8 -3 16 105
use FILL  FILL_369
timestamp 1712256841
transform 1 0 944 0 1 2970
box -8 -3 16 105
use FILL  FILL_370
timestamp 1712256841
transform 1 0 880 0 1 2970
box -8 -3 16 105
use FILL  FILL_371
timestamp 1712256841
transform 1 0 872 0 1 2970
box -8 -3 16 105
use FILL  FILL_372
timestamp 1712256841
transform 1 0 864 0 1 2970
box -8 -3 16 105
use FILL  FILL_373
timestamp 1712256841
transform 1 0 776 0 1 2970
box -8 -3 16 105
use FILL  FILL_374
timestamp 1712256841
transform 1 0 768 0 1 2970
box -8 -3 16 105
use FILL  FILL_375
timestamp 1712256841
transform 1 0 760 0 1 2970
box -8 -3 16 105
use FILL  FILL_376
timestamp 1712256841
transform 1 0 640 0 1 2970
box -8 -3 16 105
use FILL  FILL_377
timestamp 1712256841
transform 1 0 632 0 1 2970
box -8 -3 16 105
use FILL  FILL_378
timestamp 1712256841
transform 1 0 560 0 1 2970
box -8 -3 16 105
use FILL  FILL_379
timestamp 1712256841
transform 1 0 552 0 1 2970
box -8 -3 16 105
use FILL  FILL_380
timestamp 1712256841
transform 1 0 504 0 1 2970
box -8 -3 16 105
use FILL  FILL_381
timestamp 1712256841
transform 1 0 496 0 1 2970
box -8 -3 16 105
use FILL  FILL_382
timestamp 1712256841
transform 1 0 440 0 1 2970
box -8 -3 16 105
use FILL  FILL_383
timestamp 1712256841
transform 1 0 336 0 1 2970
box -8 -3 16 105
use FILL  FILL_384
timestamp 1712256841
transform 1 0 232 0 1 2970
box -8 -3 16 105
use FILL  FILL_385
timestamp 1712256841
transform 1 0 224 0 1 2970
box -8 -3 16 105
use FILL  FILL_386
timestamp 1712256841
transform 1 0 72 0 1 2970
box -8 -3 16 105
use FILL  FILL_387
timestamp 1712256841
transform 1 0 3232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_388
timestamp 1712256841
transform 1 0 3224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_389
timestamp 1712256841
transform 1 0 3200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_390
timestamp 1712256841
transform 1 0 3192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_391
timestamp 1712256841
transform 1 0 3128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_392
timestamp 1712256841
transform 1 0 3120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_393
timestamp 1712256841
transform 1 0 3112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_394
timestamp 1712256841
transform 1 0 3016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_395
timestamp 1712256841
transform 1 0 3008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_396
timestamp 1712256841
transform 1 0 2904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_397
timestamp 1712256841
transform 1 0 2800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_398
timestamp 1712256841
transform 1 0 2680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_399
timestamp 1712256841
transform 1 0 2576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_400
timestamp 1712256841
transform 1 0 2568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_401
timestamp 1712256841
transform 1 0 2560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_402
timestamp 1712256841
transform 1 0 2504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_403
timestamp 1712256841
transform 1 0 2480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_404
timestamp 1712256841
transform 1 0 2472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_405
timestamp 1712256841
transform 1 0 2440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_406
timestamp 1712256841
transform 1 0 2432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_407
timestamp 1712256841
transform 1 0 2368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_408
timestamp 1712256841
transform 1 0 2360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_409
timestamp 1712256841
transform 1 0 2352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_410
timestamp 1712256841
transform 1 0 2344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_411
timestamp 1712256841
transform 1 0 2280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_412
timestamp 1712256841
transform 1 0 2272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_413
timestamp 1712256841
transform 1 0 2264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_414
timestamp 1712256841
transform 1 0 2200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_415
timestamp 1712256841
transform 1 0 2144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_416
timestamp 1712256841
transform 1 0 2040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_417
timestamp 1712256841
transform 1 0 2032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_418
timestamp 1712256841
transform 1 0 2024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_419
timestamp 1712256841
transform 1 0 1968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_420
timestamp 1712256841
transform 1 0 1960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_421
timestamp 1712256841
transform 1 0 1880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_422
timestamp 1712256841
transform 1 0 1872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_423
timestamp 1712256841
transform 1 0 1864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_424
timestamp 1712256841
transform 1 0 1840 0 -1 2970
box -8 -3 16 105
use FILL  FILL_425
timestamp 1712256841
transform 1 0 1832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_426
timestamp 1712256841
transform 1 0 1752 0 -1 2970
box -8 -3 16 105
use FILL  FILL_427
timestamp 1712256841
transform 1 0 1744 0 -1 2970
box -8 -3 16 105
use FILL  FILL_428
timestamp 1712256841
transform 1 0 1736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_429
timestamp 1712256841
transform 1 0 1696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_430
timestamp 1712256841
transform 1 0 1688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_431
timestamp 1712256841
transform 1 0 1640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_432
timestamp 1712256841
transform 1 0 1632 0 -1 2970
box -8 -3 16 105
use FILL  FILL_433
timestamp 1712256841
transform 1 0 1584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_434
timestamp 1712256841
transform 1 0 1576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_435
timestamp 1712256841
transform 1 0 1568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_436
timestamp 1712256841
transform 1 0 1504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_437
timestamp 1712256841
transform 1 0 1496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_438
timestamp 1712256841
transform 1 0 1488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_439
timestamp 1712256841
transform 1 0 1424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_440
timestamp 1712256841
transform 1 0 1384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_441
timestamp 1712256841
transform 1 0 1376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_442
timestamp 1712256841
transform 1 0 1272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_443
timestamp 1712256841
transform 1 0 1248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_444
timestamp 1712256841
transform 1 0 1240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_445
timestamp 1712256841
transform 1 0 1160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_446
timestamp 1712256841
transform 1 0 1152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_447
timestamp 1712256841
transform 1 0 1144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_448
timestamp 1712256841
transform 1 0 1040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_449
timestamp 1712256841
transform 1 0 1032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_450
timestamp 1712256841
transform 1 0 1024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_451
timestamp 1712256841
transform 1 0 960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_452
timestamp 1712256841
transform 1 0 920 0 -1 2970
box -8 -3 16 105
use FILL  FILL_453
timestamp 1712256841
transform 1 0 872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_454
timestamp 1712256841
transform 1 0 864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_455
timestamp 1712256841
transform 1 0 784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_456
timestamp 1712256841
transform 1 0 776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_457
timestamp 1712256841
transform 1 0 768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_458
timestamp 1712256841
transform 1 0 760 0 -1 2970
box -8 -3 16 105
use FILL  FILL_459
timestamp 1712256841
transform 1 0 680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_460
timestamp 1712256841
transform 1 0 672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_461
timestamp 1712256841
transform 1 0 664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_462
timestamp 1712256841
transform 1 0 576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_463
timestamp 1712256841
transform 1 0 568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_464
timestamp 1712256841
transform 1 0 560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_465
timestamp 1712256841
transform 1 0 552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_466
timestamp 1712256841
transform 1 0 544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_467
timestamp 1712256841
transform 1 0 472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_468
timestamp 1712256841
transform 1 0 464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_469
timestamp 1712256841
transform 1 0 456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_470
timestamp 1712256841
transform 1 0 352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_471
timestamp 1712256841
transform 1 0 344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_472
timestamp 1712256841
transform 1 0 336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_473
timestamp 1712256841
transform 1 0 328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_474
timestamp 1712256841
transform 1 0 248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_475
timestamp 1712256841
transform 1 0 240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_476
timestamp 1712256841
transform 1 0 232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_477
timestamp 1712256841
transform 1 0 224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_478
timestamp 1712256841
transform 1 0 216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_479
timestamp 1712256841
transform 1 0 184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_480
timestamp 1712256841
transform 1 0 128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_481
timestamp 1712256841
transform 1 0 120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_482
timestamp 1712256841
transform 1 0 112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_483
timestamp 1712256841
transform 1 0 104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_484
timestamp 1712256841
transform 1 0 96 0 -1 2970
box -8 -3 16 105
use FILL  FILL_485
timestamp 1712256841
transform 1 0 88 0 -1 2970
box -8 -3 16 105
use FILL  FILL_486
timestamp 1712256841
transform 1 0 80 0 -1 2970
box -8 -3 16 105
use FILL  FILL_487
timestamp 1712256841
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_488
timestamp 1712256841
transform 1 0 3424 0 1 2770
box -8 -3 16 105
use FILL  FILL_489
timestamp 1712256841
transform 1 0 3320 0 1 2770
box -8 -3 16 105
use FILL  FILL_490
timestamp 1712256841
transform 1 0 3312 0 1 2770
box -8 -3 16 105
use FILL  FILL_491
timestamp 1712256841
transform 1 0 3256 0 1 2770
box -8 -3 16 105
use FILL  FILL_492
timestamp 1712256841
transform 1 0 3248 0 1 2770
box -8 -3 16 105
use FILL  FILL_493
timestamp 1712256841
transform 1 0 3240 0 1 2770
box -8 -3 16 105
use FILL  FILL_494
timestamp 1712256841
transform 1 0 3232 0 1 2770
box -8 -3 16 105
use FILL  FILL_495
timestamp 1712256841
transform 1 0 3224 0 1 2770
box -8 -3 16 105
use FILL  FILL_496
timestamp 1712256841
transform 1 0 3216 0 1 2770
box -8 -3 16 105
use FILL  FILL_497
timestamp 1712256841
transform 1 0 3152 0 1 2770
box -8 -3 16 105
use FILL  FILL_498
timestamp 1712256841
transform 1 0 3144 0 1 2770
box -8 -3 16 105
use FILL  FILL_499
timestamp 1712256841
transform 1 0 3136 0 1 2770
box -8 -3 16 105
use FILL  FILL_500
timestamp 1712256841
transform 1 0 3128 0 1 2770
box -8 -3 16 105
use FILL  FILL_501
timestamp 1712256841
transform 1 0 3120 0 1 2770
box -8 -3 16 105
use FILL  FILL_502
timestamp 1712256841
transform 1 0 3112 0 1 2770
box -8 -3 16 105
use FILL  FILL_503
timestamp 1712256841
transform 1 0 3040 0 1 2770
box -8 -3 16 105
use FILL  FILL_504
timestamp 1712256841
transform 1 0 3032 0 1 2770
box -8 -3 16 105
use FILL  FILL_505
timestamp 1712256841
transform 1 0 3024 0 1 2770
box -8 -3 16 105
use FILL  FILL_506
timestamp 1712256841
transform 1 0 3016 0 1 2770
box -8 -3 16 105
use FILL  FILL_507
timestamp 1712256841
transform 1 0 2920 0 1 2770
box -8 -3 16 105
use FILL  FILL_508
timestamp 1712256841
transform 1 0 2912 0 1 2770
box -8 -3 16 105
use FILL  FILL_509
timestamp 1712256841
transform 1 0 2904 0 1 2770
box -8 -3 16 105
use FILL  FILL_510
timestamp 1712256841
transform 1 0 2896 0 1 2770
box -8 -3 16 105
use FILL  FILL_511
timestamp 1712256841
transform 1 0 2888 0 1 2770
box -8 -3 16 105
use FILL  FILL_512
timestamp 1712256841
transform 1 0 2800 0 1 2770
box -8 -3 16 105
use FILL  FILL_513
timestamp 1712256841
transform 1 0 2792 0 1 2770
box -8 -3 16 105
use FILL  FILL_514
timestamp 1712256841
transform 1 0 2784 0 1 2770
box -8 -3 16 105
use FILL  FILL_515
timestamp 1712256841
transform 1 0 2776 0 1 2770
box -8 -3 16 105
use FILL  FILL_516
timestamp 1712256841
transform 1 0 2768 0 1 2770
box -8 -3 16 105
use FILL  FILL_517
timestamp 1712256841
transform 1 0 2696 0 1 2770
box -8 -3 16 105
use FILL  FILL_518
timestamp 1712256841
transform 1 0 2688 0 1 2770
box -8 -3 16 105
use FILL  FILL_519
timestamp 1712256841
transform 1 0 2680 0 1 2770
box -8 -3 16 105
use FILL  FILL_520
timestamp 1712256841
transform 1 0 2672 0 1 2770
box -8 -3 16 105
use FILL  FILL_521
timestamp 1712256841
transform 1 0 2640 0 1 2770
box -8 -3 16 105
use FILL  FILL_522
timestamp 1712256841
transform 1 0 2632 0 1 2770
box -8 -3 16 105
use FILL  FILL_523
timestamp 1712256841
transform 1 0 2600 0 1 2770
box -8 -3 16 105
use FILL  FILL_524
timestamp 1712256841
transform 1 0 2568 0 1 2770
box -8 -3 16 105
use FILL  FILL_525
timestamp 1712256841
transform 1 0 2560 0 1 2770
box -8 -3 16 105
use FILL  FILL_526
timestamp 1712256841
transform 1 0 2456 0 1 2770
box -8 -3 16 105
use FILL  FILL_527
timestamp 1712256841
transform 1 0 2448 0 1 2770
box -8 -3 16 105
use FILL  FILL_528
timestamp 1712256841
transform 1 0 2440 0 1 2770
box -8 -3 16 105
use FILL  FILL_529
timestamp 1712256841
transform 1 0 2432 0 1 2770
box -8 -3 16 105
use FILL  FILL_530
timestamp 1712256841
transform 1 0 2376 0 1 2770
box -8 -3 16 105
use FILL  FILL_531
timestamp 1712256841
transform 1 0 2368 0 1 2770
box -8 -3 16 105
use FILL  FILL_532
timestamp 1712256841
transform 1 0 2264 0 1 2770
box -8 -3 16 105
use FILL  FILL_533
timestamp 1712256841
transform 1 0 2256 0 1 2770
box -8 -3 16 105
use FILL  FILL_534
timestamp 1712256841
transform 1 0 2200 0 1 2770
box -8 -3 16 105
use FILL  FILL_535
timestamp 1712256841
transform 1 0 2096 0 1 2770
box -8 -3 16 105
use FILL  FILL_536
timestamp 1712256841
transform 1 0 2088 0 1 2770
box -8 -3 16 105
use FILL  FILL_537
timestamp 1712256841
transform 1 0 2032 0 1 2770
box -8 -3 16 105
use FILL  FILL_538
timestamp 1712256841
transform 1 0 1928 0 1 2770
box -8 -3 16 105
use FILL  FILL_539
timestamp 1712256841
transform 1 0 1920 0 1 2770
box -8 -3 16 105
use FILL  FILL_540
timestamp 1712256841
transform 1 0 1784 0 1 2770
box -8 -3 16 105
use FILL  FILL_541
timestamp 1712256841
transform 1 0 1776 0 1 2770
box -8 -3 16 105
use FILL  FILL_542
timestamp 1712256841
transform 1 0 1624 0 1 2770
box -8 -3 16 105
use FILL  FILL_543
timestamp 1712256841
transform 1 0 1616 0 1 2770
box -8 -3 16 105
use FILL  FILL_544
timestamp 1712256841
transform 1 0 1512 0 1 2770
box -8 -3 16 105
use FILL  FILL_545
timestamp 1712256841
transform 1 0 1504 0 1 2770
box -8 -3 16 105
use FILL  FILL_546
timestamp 1712256841
transform 1 0 1480 0 1 2770
box -8 -3 16 105
use FILL  FILL_547
timestamp 1712256841
transform 1 0 1456 0 1 2770
box -8 -3 16 105
use FILL  FILL_548
timestamp 1712256841
transform 1 0 1352 0 1 2770
box -8 -3 16 105
use FILL  FILL_549
timestamp 1712256841
transform 1 0 1344 0 1 2770
box -8 -3 16 105
use FILL  FILL_550
timestamp 1712256841
transform 1 0 1336 0 1 2770
box -8 -3 16 105
use FILL  FILL_551
timestamp 1712256841
transform 1 0 1328 0 1 2770
box -8 -3 16 105
use FILL  FILL_552
timestamp 1712256841
transform 1 0 1272 0 1 2770
box -8 -3 16 105
use FILL  FILL_553
timestamp 1712256841
transform 1 0 1264 0 1 2770
box -8 -3 16 105
use FILL  FILL_554
timestamp 1712256841
transform 1 0 1256 0 1 2770
box -8 -3 16 105
use FILL  FILL_555
timestamp 1712256841
transform 1 0 1216 0 1 2770
box -8 -3 16 105
use FILL  FILL_556
timestamp 1712256841
transform 1 0 1208 0 1 2770
box -8 -3 16 105
use FILL  FILL_557
timestamp 1712256841
transform 1 0 1200 0 1 2770
box -8 -3 16 105
use FILL  FILL_558
timestamp 1712256841
transform 1 0 1096 0 1 2770
box -8 -3 16 105
use FILL  FILL_559
timestamp 1712256841
transform 1 0 1088 0 1 2770
box -8 -3 16 105
use FILL  FILL_560
timestamp 1712256841
transform 1 0 1080 0 1 2770
box -8 -3 16 105
use FILL  FILL_561
timestamp 1712256841
transform 1 0 1072 0 1 2770
box -8 -3 16 105
use FILL  FILL_562
timestamp 1712256841
transform 1 0 1048 0 1 2770
box -8 -3 16 105
use FILL  FILL_563
timestamp 1712256841
transform 1 0 1008 0 1 2770
box -8 -3 16 105
use FILL  FILL_564
timestamp 1712256841
transform 1 0 1000 0 1 2770
box -8 -3 16 105
use FILL  FILL_565
timestamp 1712256841
transform 1 0 992 0 1 2770
box -8 -3 16 105
use FILL  FILL_566
timestamp 1712256841
transform 1 0 984 0 1 2770
box -8 -3 16 105
use FILL  FILL_567
timestamp 1712256841
transform 1 0 976 0 1 2770
box -8 -3 16 105
use FILL  FILL_568
timestamp 1712256841
transform 1 0 968 0 1 2770
box -8 -3 16 105
use FILL  FILL_569
timestamp 1712256841
transform 1 0 944 0 1 2770
box -8 -3 16 105
use FILL  FILL_570
timestamp 1712256841
transform 1 0 912 0 1 2770
box -8 -3 16 105
use FILL  FILL_571
timestamp 1712256841
transform 1 0 904 0 1 2770
box -8 -3 16 105
use FILL  FILL_572
timestamp 1712256841
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_573
timestamp 1712256841
transform 1 0 856 0 1 2770
box -8 -3 16 105
use FILL  FILL_574
timestamp 1712256841
transform 1 0 848 0 1 2770
box -8 -3 16 105
use FILL  FILL_575
timestamp 1712256841
transform 1 0 840 0 1 2770
box -8 -3 16 105
use FILL  FILL_576
timestamp 1712256841
transform 1 0 800 0 1 2770
box -8 -3 16 105
use FILL  FILL_577
timestamp 1712256841
transform 1 0 792 0 1 2770
box -8 -3 16 105
use FILL  FILL_578
timestamp 1712256841
transform 1 0 768 0 1 2770
box -8 -3 16 105
use FILL  FILL_579
timestamp 1712256841
transform 1 0 760 0 1 2770
box -8 -3 16 105
use FILL  FILL_580
timestamp 1712256841
transform 1 0 712 0 1 2770
box -8 -3 16 105
use FILL  FILL_581
timestamp 1712256841
transform 1 0 704 0 1 2770
box -8 -3 16 105
use FILL  FILL_582
timestamp 1712256841
transform 1 0 696 0 1 2770
box -8 -3 16 105
use FILL  FILL_583
timestamp 1712256841
transform 1 0 688 0 1 2770
box -8 -3 16 105
use FILL  FILL_584
timestamp 1712256841
transform 1 0 632 0 1 2770
box -8 -3 16 105
use FILL  FILL_585
timestamp 1712256841
transform 1 0 624 0 1 2770
box -8 -3 16 105
use FILL  FILL_586
timestamp 1712256841
transform 1 0 616 0 1 2770
box -8 -3 16 105
use FILL  FILL_587
timestamp 1712256841
transform 1 0 512 0 1 2770
box -8 -3 16 105
use FILL  FILL_588
timestamp 1712256841
transform 1 0 504 0 1 2770
box -8 -3 16 105
use FILL  FILL_589
timestamp 1712256841
transform 1 0 496 0 1 2770
box -8 -3 16 105
use FILL  FILL_590
timestamp 1712256841
transform 1 0 488 0 1 2770
box -8 -3 16 105
use FILL  FILL_591
timestamp 1712256841
transform 1 0 408 0 1 2770
box -8 -3 16 105
use FILL  FILL_592
timestamp 1712256841
transform 1 0 400 0 1 2770
box -8 -3 16 105
use FILL  FILL_593
timestamp 1712256841
transform 1 0 392 0 1 2770
box -8 -3 16 105
use FILL  FILL_594
timestamp 1712256841
transform 1 0 288 0 1 2770
box -8 -3 16 105
use FILL  FILL_595
timestamp 1712256841
transform 1 0 280 0 1 2770
box -8 -3 16 105
use FILL  FILL_596
timestamp 1712256841
transform 1 0 176 0 1 2770
box -8 -3 16 105
use FILL  FILL_597
timestamp 1712256841
transform 1 0 168 0 1 2770
box -8 -3 16 105
use FILL  FILL_598
timestamp 1712256841
transform 1 0 3424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_599
timestamp 1712256841
transform 1 0 3320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_600
timestamp 1712256841
transform 1 0 3312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_601
timestamp 1712256841
transform 1 0 3304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_602
timestamp 1712256841
transform 1 0 3296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_603
timestamp 1712256841
transform 1 0 3248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_604
timestamp 1712256841
transform 1 0 3240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_605
timestamp 1712256841
transform 1 0 3232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_606
timestamp 1712256841
transform 1 0 3224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_607
timestamp 1712256841
transform 1 0 3216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_608
timestamp 1712256841
transform 1 0 3208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_609
timestamp 1712256841
transform 1 0 3152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_610
timestamp 1712256841
transform 1 0 3144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_611
timestamp 1712256841
transform 1 0 3136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_612
timestamp 1712256841
transform 1 0 3032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_613
timestamp 1712256841
transform 1 0 3024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_614
timestamp 1712256841
transform 1 0 3016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_615
timestamp 1712256841
transform 1 0 2984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_616
timestamp 1712256841
transform 1 0 2976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_617
timestamp 1712256841
transform 1 0 2872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_618
timestamp 1712256841
transform 1 0 2864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_619
timestamp 1712256841
transform 1 0 2856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_620
timestamp 1712256841
transform 1 0 2752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_621
timestamp 1712256841
transform 1 0 2744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_622
timestamp 1712256841
transform 1 0 2736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_623
timestamp 1712256841
transform 1 0 2632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_624
timestamp 1712256841
transform 1 0 2624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_625
timestamp 1712256841
transform 1 0 2520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_626
timestamp 1712256841
transform 1 0 2512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_627
timestamp 1712256841
transform 1 0 2504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_628
timestamp 1712256841
transform 1 0 2400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_629
timestamp 1712256841
transform 1 0 2368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_630
timestamp 1712256841
transform 1 0 2360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_631
timestamp 1712256841
transform 1 0 2352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_632
timestamp 1712256841
transform 1 0 2248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_633
timestamp 1712256841
transform 1 0 2240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_634
timestamp 1712256841
transform 1 0 2208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_635
timestamp 1712256841
transform 1 0 2200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_636
timestamp 1712256841
transform 1 0 2096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_637
timestamp 1712256841
transform 1 0 2088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_638
timestamp 1712256841
transform 1 0 2080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_639
timestamp 1712256841
transform 1 0 2072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_640
timestamp 1712256841
transform 1 0 2016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_641
timestamp 1712256841
transform 1 0 2008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_642
timestamp 1712256841
transform 1 0 2000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_643
timestamp 1712256841
transform 1 0 1992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_644
timestamp 1712256841
transform 1 0 1944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_645
timestamp 1712256841
transform 1 0 1936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_646
timestamp 1712256841
transform 1 0 1928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_647
timestamp 1712256841
transform 1 0 1920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_648
timestamp 1712256841
transform 1 0 1912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_649
timestamp 1712256841
transform 1 0 1904 0 -1 2770
box -8 -3 16 105
use FILL  FILL_650
timestamp 1712256841
transform 1 0 1856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_651
timestamp 1712256841
transform 1 0 1848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_652
timestamp 1712256841
transform 1 0 1816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_653
timestamp 1712256841
transform 1 0 1808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_654
timestamp 1712256841
transform 1 0 1800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_655
timestamp 1712256841
transform 1 0 1776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_656
timestamp 1712256841
transform 1 0 1768 0 -1 2770
box -8 -3 16 105
use FILL  FILL_657
timestamp 1712256841
transform 1 0 1760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_658
timestamp 1712256841
transform 1 0 1752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_659
timestamp 1712256841
transform 1 0 1744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_660
timestamp 1712256841
transform 1 0 1696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_661
timestamp 1712256841
transform 1 0 1688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_662
timestamp 1712256841
transform 1 0 1680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_663
timestamp 1712256841
transform 1 0 1672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_664
timestamp 1712256841
transform 1 0 1568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_665
timestamp 1712256841
transform 1 0 1560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_666
timestamp 1712256841
transform 1 0 1552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_667
timestamp 1712256841
transform 1 0 1544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_668
timestamp 1712256841
transform 1 0 1496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_669
timestamp 1712256841
transform 1 0 1488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_670
timestamp 1712256841
transform 1 0 1480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_671
timestamp 1712256841
transform 1 0 1424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_672
timestamp 1712256841
transform 1 0 1416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_673
timestamp 1712256841
transform 1 0 1408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_674
timestamp 1712256841
transform 1 0 1400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_675
timestamp 1712256841
transform 1 0 1296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_676
timestamp 1712256841
transform 1 0 1288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_677
timestamp 1712256841
transform 1 0 1280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_678
timestamp 1712256841
transform 1 0 1272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_679
timestamp 1712256841
transform 1 0 1224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_680
timestamp 1712256841
transform 1 0 1216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_681
timestamp 1712256841
transform 1 0 1208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_682
timestamp 1712256841
transform 1 0 1160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_683
timestamp 1712256841
transform 1 0 1152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_684
timestamp 1712256841
transform 1 0 1144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_685
timestamp 1712256841
transform 1 0 1136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_686
timestamp 1712256841
transform 1 0 1128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_687
timestamp 1712256841
transform 1 0 1120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_688
timestamp 1712256841
transform 1 0 1088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_689
timestamp 1712256841
transform 1 0 1040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_690
timestamp 1712256841
transform 1 0 1032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_691
timestamp 1712256841
transform 1 0 1024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_692
timestamp 1712256841
transform 1 0 920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_693
timestamp 1712256841
transform 1 0 912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_694
timestamp 1712256841
transform 1 0 904 0 -1 2770
box -8 -3 16 105
use FILL  FILL_695
timestamp 1712256841
transform 1 0 896 0 -1 2770
box -8 -3 16 105
use FILL  FILL_696
timestamp 1712256841
transform 1 0 888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_697
timestamp 1712256841
transform 1 0 840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_698
timestamp 1712256841
transform 1 0 832 0 -1 2770
box -8 -3 16 105
use FILL  FILL_699
timestamp 1712256841
transform 1 0 824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_700
timestamp 1712256841
transform 1 0 720 0 -1 2770
box -8 -3 16 105
use FILL  FILL_701
timestamp 1712256841
transform 1 0 712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_702
timestamp 1712256841
transform 1 0 704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_703
timestamp 1712256841
transform 1 0 696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_704
timestamp 1712256841
transform 1 0 688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_705
timestamp 1712256841
transform 1 0 648 0 -1 2770
box -8 -3 16 105
use FILL  FILL_706
timestamp 1712256841
transform 1 0 640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_707
timestamp 1712256841
transform 1 0 608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_708
timestamp 1712256841
transform 1 0 600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_709
timestamp 1712256841
transform 1 0 592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_710
timestamp 1712256841
transform 1 0 584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_711
timestamp 1712256841
transform 1 0 576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_712
timestamp 1712256841
transform 1 0 528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_713
timestamp 1712256841
transform 1 0 520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_714
timestamp 1712256841
transform 1 0 512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_715
timestamp 1712256841
transform 1 0 504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_716
timestamp 1712256841
transform 1 0 400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_717
timestamp 1712256841
transform 1 0 392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_718
timestamp 1712256841
transform 1 0 384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_719
timestamp 1712256841
transform 1 0 280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_720
timestamp 1712256841
transform 1 0 272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_721
timestamp 1712256841
transform 1 0 264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_722
timestamp 1712256841
transform 1 0 256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_723
timestamp 1712256841
transform 1 0 248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_724
timestamp 1712256841
transform 1 0 240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_725
timestamp 1712256841
transform 1 0 232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_726
timestamp 1712256841
transform 1 0 224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_727
timestamp 1712256841
transform 1 0 120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_728
timestamp 1712256841
transform 1 0 112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_729
timestamp 1712256841
transform 1 0 104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_730
timestamp 1712256841
transform 1 0 96 0 -1 2770
box -8 -3 16 105
use FILL  FILL_731
timestamp 1712256841
transform 1 0 88 0 -1 2770
box -8 -3 16 105
use FILL  FILL_732
timestamp 1712256841
transform 1 0 80 0 -1 2770
box -8 -3 16 105
use FILL  FILL_733
timestamp 1712256841
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_734
timestamp 1712256841
transform 1 0 3424 0 1 2570
box -8 -3 16 105
use FILL  FILL_735
timestamp 1712256841
transform 1 0 3416 0 1 2570
box -8 -3 16 105
use FILL  FILL_736
timestamp 1712256841
transform 1 0 3408 0 1 2570
box -8 -3 16 105
use FILL  FILL_737
timestamp 1712256841
transform 1 0 3376 0 1 2570
box -8 -3 16 105
use FILL  FILL_738
timestamp 1712256841
transform 1 0 3368 0 1 2570
box -8 -3 16 105
use FILL  FILL_739
timestamp 1712256841
transform 1 0 3360 0 1 2570
box -8 -3 16 105
use FILL  FILL_740
timestamp 1712256841
transform 1 0 3352 0 1 2570
box -8 -3 16 105
use FILL  FILL_741
timestamp 1712256841
transform 1 0 3344 0 1 2570
box -8 -3 16 105
use FILL  FILL_742
timestamp 1712256841
transform 1 0 3296 0 1 2570
box -8 -3 16 105
use FILL  FILL_743
timestamp 1712256841
transform 1 0 3288 0 1 2570
box -8 -3 16 105
use FILL  FILL_744
timestamp 1712256841
transform 1 0 3280 0 1 2570
box -8 -3 16 105
use FILL  FILL_745
timestamp 1712256841
transform 1 0 3272 0 1 2570
box -8 -3 16 105
use FILL  FILL_746
timestamp 1712256841
transform 1 0 3264 0 1 2570
box -8 -3 16 105
use FILL  FILL_747
timestamp 1712256841
transform 1 0 3216 0 1 2570
box -8 -3 16 105
use FILL  FILL_748
timestamp 1712256841
transform 1 0 3208 0 1 2570
box -8 -3 16 105
use FILL  FILL_749
timestamp 1712256841
transform 1 0 3200 0 1 2570
box -8 -3 16 105
use FILL  FILL_750
timestamp 1712256841
transform 1 0 3192 0 1 2570
box -8 -3 16 105
use FILL  FILL_751
timestamp 1712256841
transform 1 0 3184 0 1 2570
box -8 -3 16 105
use FILL  FILL_752
timestamp 1712256841
transform 1 0 3176 0 1 2570
box -8 -3 16 105
use FILL  FILL_753
timestamp 1712256841
transform 1 0 3136 0 1 2570
box -8 -3 16 105
use FILL  FILL_754
timestamp 1712256841
transform 1 0 3128 0 1 2570
box -8 -3 16 105
use FILL  FILL_755
timestamp 1712256841
transform 1 0 3120 0 1 2570
box -8 -3 16 105
use FILL  FILL_756
timestamp 1712256841
transform 1 0 3112 0 1 2570
box -8 -3 16 105
use FILL  FILL_757
timestamp 1712256841
transform 1 0 3104 0 1 2570
box -8 -3 16 105
use FILL  FILL_758
timestamp 1712256841
transform 1 0 3064 0 1 2570
box -8 -3 16 105
use FILL  FILL_759
timestamp 1712256841
transform 1 0 3056 0 1 2570
box -8 -3 16 105
use FILL  FILL_760
timestamp 1712256841
transform 1 0 3016 0 1 2570
box -8 -3 16 105
use FILL  FILL_761
timestamp 1712256841
transform 1 0 3008 0 1 2570
box -8 -3 16 105
use FILL  FILL_762
timestamp 1712256841
transform 1 0 3000 0 1 2570
box -8 -3 16 105
use FILL  FILL_763
timestamp 1712256841
transform 1 0 2992 0 1 2570
box -8 -3 16 105
use FILL  FILL_764
timestamp 1712256841
transform 1 0 2984 0 1 2570
box -8 -3 16 105
use FILL  FILL_765
timestamp 1712256841
transform 1 0 2880 0 1 2570
box -8 -3 16 105
use FILL  FILL_766
timestamp 1712256841
transform 1 0 2872 0 1 2570
box -8 -3 16 105
use FILL  FILL_767
timestamp 1712256841
transform 1 0 2864 0 1 2570
box -8 -3 16 105
use FILL  FILL_768
timestamp 1712256841
transform 1 0 2856 0 1 2570
box -8 -3 16 105
use FILL  FILL_769
timestamp 1712256841
transform 1 0 2808 0 1 2570
box -8 -3 16 105
use FILL  FILL_770
timestamp 1712256841
transform 1 0 2800 0 1 2570
box -8 -3 16 105
use FILL  FILL_771
timestamp 1712256841
transform 1 0 2792 0 1 2570
box -8 -3 16 105
use FILL  FILL_772
timestamp 1712256841
transform 1 0 2784 0 1 2570
box -8 -3 16 105
use FILL  FILL_773
timestamp 1712256841
transform 1 0 2776 0 1 2570
box -8 -3 16 105
use FILL  FILL_774
timestamp 1712256841
transform 1 0 2672 0 1 2570
box -8 -3 16 105
use FILL  FILL_775
timestamp 1712256841
transform 1 0 2664 0 1 2570
box -8 -3 16 105
use FILL  FILL_776
timestamp 1712256841
transform 1 0 2656 0 1 2570
box -8 -3 16 105
use FILL  FILL_777
timestamp 1712256841
transform 1 0 2648 0 1 2570
box -8 -3 16 105
use FILL  FILL_778
timestamp 1712256841
transform 1 0 2640 0 1 2570
box -8 -3 16 105
use FILL  FILL_779
timestamp 1712256841
transform 1 0 2592 0 1 2570
box -8 -3 16 105
use FILL  FILL_780
timestamp 1712256841
transform 1 0 2584 0 1 2570
box -8 -3 16 105
use FILL  FILL_781
timestamp 1712256841
transform 1 0 2576 0 1 2570
box -8 -3 16 105
use FILL  FILL_782
timestamp 1712256841
transform 1 0 2552 0 1 2570
box -8 -3 16 105
use FILL  FILL_783
timestamp 1712256841
transform 1 0 2544 0 1 2570
box -8 -3 16 105
use FILL  FILL_784
timestamp 1712256841
transform 1 0 2536 0 1 2570
box -8 -3 16 105
use FILL  FILL_785
timestamp 1712256841
transform 1 0 2528 0 1 2570
box -8 -3 16 105
use FILL  FILL_786
timestamp 1712256841
transform 1 0 2480 0 1 2570
box -8 -3 16 105
use FILL  FILL_787
timestamp 1712256841
transform 1 0 2472 0 1 2570
box -8 -3 16 105
use FILL  FILL_788
timestamp 1712256841
transform 1 0 2464 0 1 2570
box -8 -3 16 105
use FILL  FILL_789
timestamp 1712256841
transform 1 0 2456 0 1 2570
box -8 -3 16 105
use FILL  FILL_790
timestamp 1712256841
transform 1 0 2448 0 1 2570
box -8 -3 16 105
use FILL  FILL_791
timestamp 1712256841
transform 1 0 2440 0 1 2570
box -8 -3 16 105
use FILL  FILL_792
timestamp 1712256841
transform 1 0 2392 0 1 2570
box -8 -3 16 105
use FILL  FILL_793
timestamp 1712256841
transform 1 0 2384 0 1 2570
box -8 -3 16 105
use FILL  FILL_794
timestamp 1712256841
transform 1 0 2328 0 1 2570
box -8 -3 16 105
use FILL  FILL_795
timestamp 1712256841
transform 1 0 2320 0 1 2570
box -8 -3 16 105
use FILL  FILL_796
timestamp 1712256841
transform 1 0 2312 0 1 2570
box -8 -3 16 105
use FILL  FILL_797
timestamp 1712256841
transform 1 0 2304 0 1 2570
box -8 -3 16 105
use FILL  FILL_798
timestamp 1712256841
transform 1 0 2152 0 1 2570
box -8 -3 16 105
use FILL  FILL_799
timestamp 1712256841
transform 1 0 2048 0 1 2570
box -8 -3 16 105
use FILL  FILL_800
timestamp 1712256841
transform 1 0 1944 0 1 2570
box -8 -3 16 105
use FILL  FILL_801
timestamp 1712256841
transform 1 0 1840 0 1 2570
box -8 -3 16 105
use FILL  FILL_802
timestamp 1712256841
transform 1 0 1640 0 1 2570
box -8 -3 16 105
use FILL  FILL_803
timestamp 1712256841
transform 1 0 1632 0 1 2570
box -8 -3 16 105
use FILL  FILL_804
timestamp 1712256841
transform 1 0 1528 0 1 2570
box -8 -3 16 105
use FILL  FILL_805
timestamp 1712256841
transform 1 0 1424 0 1 2570
box -8 -3 16 105
use FILL  FILL_806
timestamp 1712256841
transform 1 0 1416 0 1 2570
box -8 -3 16 105
use FILL  FILL_807
timestamp 1712256841
transform 1 0 1312 0 1 2570
box -8 -3 16 105
use FILL  FILL_808
timestamp 1712256841
transform 1 0 1208 0 1 2570
box -8 -3 16 105
use FILL  FILL_809
timestamp 1712256841
transform 1 0 1200 0 1 2570
box -8 -3 16 105
use FILL  FILL_810
timestamp 1712256841
transform 1 0 1096 0 1 2570
box -8 -3 16 105
use FILL  FILL_811
timestamp 1712256841
transform 1 0 1088 0 1 2570
box -8 -3 16 105
use FILL  FILL_812
timestamp 1712256841
transform 1 0 984 0 1 2570
box -8 -3 16 105
use FILL  FILL_813
timestamp 1712256841
transform 1 0 880 0 1 2570
box -8 -3 16 105
use FILL  FILL_814
timestamp 1712256841
transform 1 0 872 0 1 2570
box -8 -3 16 105
use FILL  FILL_815
timestamp 1712256841
transform 1 0 768 0 1 2570
box -8 -3 16 105
use FILL  FILL_816
timestamp 1712256841
transform 1 0 760 0 1 2570
box -8 -3 16 105
use FILL  FILL_817
timestamp 1712256841
transform 1 0 656 0 1 2570
box -8 -3 16 105
use FILL  FILL_818
timestamp 1712256841
transform 1 0 552 0 1 2570
box -8 -3 16 105
use FILL  FILL_819
timestamp 1712256841
transform 1 0 528 0 1 2570
box -8 -3 16 105
use FILL  FILL_820
timestamp 1712256841
transform 1 0 520 0 1 2570
box -8 -3 16 105
use FILL  FILL_821
timestamp 1712256841
transform 1 0 416 0 1 2570
box -8 -3 16 105
use FILL  FILL_822
timestamp 1712256841
transform 1 0 408 0 1 2570
box -8 -3 16 105
use FILL  FILL_823
timestamp 1712256841
transform 1 0 400 0 1 2570
box -8 -3 16 105
use FILL  FILL_824
timestamp 1712256841
transform 1 0 352 0 1 2570
box -8 -3 16 105
use FILL  FILL_825
timestamp 1712256841
transform 1 0 344 0 1 2570
box -8 -3 16 105
use FILL  FILL_826
timestamp 1712256841
transform 1 0 336 0 1 2570
box -8 -3 16 105
use FILL  FILL_827
timestamp 1712256841
transform 1 0 328 0 1 2570
box -8 -3 16 105
use FILL  FILL_828
timestamp 1712256841
transform 1 0 280 0 1 2570
box -8 -3 16 105
use FILL  FILL_829
timestamp 1712256841
transform 1 0 272 0 1 2570
box -8 -3 16 105
use FILL  FILL_830
timestamp 1712256841
transform 1 0 264 0 1 2570
box -8 -3 16 105
use FILL  FILL_831
timestamp 1712256841
transform 1 0 216 0 1 2570
box -8 -3 16 105
use FILL  FILL_832
timestamp 1712256841
transform 1 0 208 0 1 2570
box -8 -3 16 105
use FILL  FILL_833
timestamp 1712256841
transform 1 0 200 0 1 2570
box -8 -3 16 105
use FILL  FILL_834
timestamp 1712256841
transform 1 0 192 0 1 2570
box -8 -3 16 105
use FILL  FILL_835
timestamp 1712256841
transform 1 0 144 0 1 2570
box -8 -3 16 105
use FILL  FILL_836
timestamp 1712256841
transform 1 0 136 0 1 2570
box -8 -3 16 105
use FILL  FILL_837
timestamp 1712256841
transform 1 0 128 0 1 2570
box -8 -3 16 105
use FILL  FILL_838
timestamp 1712256841
transform 1 0 120 0 1 2570
box -8 -3 16 105
use FILL  FILL_839
timestamp 1712256841
transform 1 0 72 0 1 2570
box -8 -3 16 105
use FILL  FILL_840
timestamp 1712256841
transform 1 0 3424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_841
timestamp 1712256841
transform 1 0 3320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_842
timestamp 1712256841
transform 1 0 3312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_843
timestamp 1712256841
transform 1 0 3304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_844
timestamp 1712256841
transform 1 0 3296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_845
timestamp 1712256841
transform 1 0 3232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_846
timestamp 1712256841
transform 1 0 3224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_847
timestamp 1712256841
transform 1 0 3216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_848
timestamp 1712256841
transform 1 0 3208 0 -1 2570
box -8 -3 16 105
use FILL  FILL_849
timestamp 1712256841
transform 1 0 3200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_850
timestamp 1712256841
transform 1 0 3160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_851
timestamp 1712256841
transform 1 0 3152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_852
timestamp 1712256841
transform 1 0 3112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_853
timestamp 1712256841
transform 1 0 3104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_854
timestamp 1712256841
transform 1 0 3096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_855
timestamp 1712256841
transform 1 0 3056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_856
timestamp 1712256841
transform 1 0 3048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_857
timestamp 1712256841
transform 1 0 3040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_858
timestamp 1712256841
transform 1 0 3032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_859
timestamp 1712256841
transform 1 0 2928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_860
timestamp 1712256841
transform 1 0 2920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_861
timestamp 1712256841
transform 1 0 2912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_862
timestamp 1712256841
transform 1 0 2904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_863
timestamp 1712256841
transform 1 0 2896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_864
timestamp 1712256841
transform 1 0 2848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_865
timestamp 1712256841
transform 1 0 2840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_866
timestamp 1712256841
transform 1 0 2832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_867
timestamp 1712256841
transform 1 0 2824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_868
timestamp 1712256841
transform 1 0 2816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_869
timestamp 1712256841
transform 1 0 2768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_870
timestamp 1712256841
transform 1 0 2760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_871
timestamp 1712256841
transform 1 0 2752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_872
timestamp 1712256841
transform 1 0 2744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_873
timestamp 1712256841
transform 1 0 2736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_874
timestamp 1712256841
transform 1 0 2728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_875
timestamp 1712256841
transform 1 0 2680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_876
timestamp 1712256841
transform 1 0 2672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_877
timestamp 1712256841
transform 1 0 2664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_878
timestamp 1712256841
transform 1 0 2656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_879
timestamp 1712256841
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_880
timestamp 1712256841
transform 1 0 2576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_881
timestamp 1712256841
transform 1 0 2568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_882
timestamp 1712256841
transform 1 0 2560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_883
timestamp 1712256841
transform 1 0 2552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_884
timestamp 1712256841
transform 1 0 2472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_885
timestamp 1712256841
transform 1 0 2440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_886
timestamp 1712256841
transform 1 0 2432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_887
timestamp 1712256841
transform 1 0 2400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_888
timestamp 1712256841
transform 1 0 2392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_889
timestamp 1712256841
transform 1 0 2384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_890
timestamp 1712256841
transform 1 0 2336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_891
timestamp 1712256841
transform 1 0 2328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_892
timestamp 1712256841
transform 1 0 2320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_893
timestamp 1712256841
transform 1 0 2312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_894
timestamp 1712256841
transform 1 0 2264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_895
timestamp 1712256841
transform 1 0 2256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_896
timestamp 1712256841
transform 1 0 2248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_897
timestamp 1712256841
transform 1 0 2240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_898
timestamp 1712256841
transform 1 0 2232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_899
timestamp 1712256841
transform 1 0 2224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_900
timestamp 1712256841
transform 1 0 2176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_901
timestamp 1712256841
transform 1 0 2144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_902
timestamp 1712256841
transform 1 0 2136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_903
timestamp 1712256841
transform 1 0 2128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_904
timestamp 1712256841
transform 1 0 2080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_905
timestamp 1712256841
transform 1 0 2072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_906
timestamp 1712256841
transform 1 0 2064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_907
timestamp 1712256841
transform 1 0 2056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_908
timestamp 1712256841
transform 1 0 2048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_909
timestamp 1712256841
transform 1 0 2000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_910
timestamp 1712256841
transform 1 0 1944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_911
timestamp 1712256841
transform 1 0 1936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_912
timestamp 1712256841
transform 1 0 1928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_913
timestamp 1712256841
transform 1 0 1920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_914
timestamp 1712256841
transform 1 0 1848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_915
timestamp 1712256841
transform 1 0 1840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_916
timestamp 1712256841
transform 1 0 1832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_917
timestamp 1712256841
transform 1 0 1824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_918
timestamp 1712256841
transform 1 0 1776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_919
timestamp 1712256841
transform 1 0 1768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_920
timestamp 1712256841
transform 1 0 1760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_921
timestamp 1712256841
transform 1 0 1752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_922
timestamp 1712256841
transform 1 0 1744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_923
timestamp 1712256841
transform 1 0 1680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_924
timestamp 1712256841
transform 1 0 1672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_925
timestamp 1712256841
transform 1 0 1664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_926
timestamp 1712256841
transform 1 0 1656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_927
timestamp 1712256841
transform 1 0 1648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_928
timestamp 1712256841
transform 1 0 1600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_929
timestamp 1712256841
transform 1 0 1552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_930
timestamp 1712256841
transform 1 0 1448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_931
timestamp 1712256841
transform 1 0 1440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_932
timestamp 1712256841
transform 1 0 1296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_933
timestamp 1712256841
transform 1 0 1288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_934
timestamp 1712256841
transform 1 0 1240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_935
timestamp 1712256841
transform 1 0 1192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_936
timestamp 1712256841
transform 1 0 1184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_937
timestamp 1712256841
transform 1 0 1080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_938
timestamp 1712256841
transform 1 0 1072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_939
timestamp 1712256841
transform 1 0 1024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_940
timestamp 1712256841
transform 1 0 920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_941
timestamp 1712256841
transform 1 0 912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_942
timestamp 1712256841
transform 1 0 904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_943
timestamp 1712256841
transform 1 0 896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_944
timestamp 1712256841
transform 1 0 848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_945
timestamp 1712256841
transform 1 0 840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_946
timestamp 1712256841
transform 1 0 832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_947
timestamp 1712256841
transform 1 0 784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_948
timestamp 1712256841
transform 1 0 776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_949
timestamp 1712256841
transform 1 0 768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_950
timestamp 1712256841
transform 1 0 760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_951
timestamp 1712256841
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_952
timestamp 1712256841
transform 1 0 744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_953
timestamp 1712256841
transform 1 0 696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_954
timestamp 1712256841
transform 1 0 688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_955
timestamp 1712256841
transform 1 0 680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_956
timestamp 1712256841
transform 1 0 672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_957
timestamp 1712256841
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_958
timestamp 1712256841
transform 1 0 656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_959
timestamp 1712256841
transform 1 0 648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_960
timestamp 1712256841
transform 1 0 600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_961
timestamp 1712256841
transform 1 0 592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_962
timestamp 1712256841
transform 1 0 584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_963
timestamp 1712256841
transform 1 0 576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_964
timestamp 1712256841
transform 1 0 568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_965
timestamp 1712256841
transform 1 0 560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_966
timestamp 1712256841
transform 1 0 552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_967
timestamp 1712256841
transform 1 0 504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_968
timestamp 1712256841
transform 1 0 496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_969
timestamp 1712256841
transform 1 0 488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_970
timestamp 1712256841
transform 1 0 480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_971
timestamp 1712256841
transform 1 0 472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_972
timestamp 1712256841
transform 1 0 464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_973
timestamp 1712256841
transform 1 0 416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_974
timestamp 1712256841
transform 1 0 408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_975
timestamp 1712256841
transform 1 0 400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_976
timestamp 1712256841
transform 1 0 392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_977
timestamp 1712256841
transform 1 0 384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_978
timestamp 1712256841
transform 1 0 280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_979
timestamp 1712256841
transform 1 0 272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_980
timestamp 1712256841
transform 1 0 264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_981
timestamp 1712256841
transform 1 0 256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_982
timestamp 1712256841
transform 1 0 248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_983
timestamp 1712256841
transform 1 0 240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_984
timestamp 1712256841
transform 1 0 232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_985
timestamp 1712256841
transform 1 0 224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_986
timestamp 1712256841
transform 1 0 120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_987
timestamp 1712256841
transform 1 0 112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_988
timestamp 1712256841
transform 1 0 104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_989
timestamp 1712256841
transform 1 0 96 0 -1 2570
box -8 -3 16 105
use FILL  FILL_990
timestamp 1712256841
transform 1 0 88 0 -1 2570
box -8 -3 16 105
use FILL  FILL_991
timestamp 1712256841
transform 1 0 80 0 -1 2570
box -8 -3 16 105
use FILL  FILL_992
timestamp 1712256841
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_993
timestamp 1712256841
transform 1 0 3424 0 1 2370
box -8 -3 16 105
use FILL  FILL_994
timestamp 1712256841
transform 1 0 3416 0 1 2370
box -8 -3 16 105
use FILL  FILL_995
timestamp 1712256841
transform 1 0 1792 0 1 2370
box -8 -3 16 105
use FILL  FILL_996
timestamp 1712256841
transform 1 0 1688 0 1 2370
box -8 -3 16 105
use FILL  FILL_997
timestamp 1712256841
transform 1 0 1680 0 1 2370
box -8 -3 16 105
use FILL  FILL_998
timestamp 1712256841
transform 1 0 1576 0 1 2370
box -8 -3 16 105
use FILL  FILL_999
timestamp 1712256841
transform 1 0 1568 0 1 2370
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1712256841
transform 1 0 1464 0 1 2370
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1712256841
transform 1 0 1456 0 1 2370
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1712256841
transform 1 0 1448 0 1 2370
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1712256841
transform 1 0 1408 0 1 2370
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1712256841
transform 1 0 1400 0 1 2370
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1712256841
transform 1 0 1392 0 1 2370
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1712256841
transform 1 0 1352 0 1 2370
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1712256841
transform 1 0 1344 0 1 2370
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1712256841
transform 1 0 1304 0 1 2370
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1712256841
transform 1 0 1296 0 1 2370
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1712256841
transform 1 0 1288 0 1 2370
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1712256841
transform 1 0 1184 0 1 2370
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1712256841
transform 1 0 1176 0 1 2370
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1712256841
transform 1 0 1168 0 1 2370
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1712256841
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1712256841
transform 1 0 1152 0 1 2370
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1712256841
transform 1 0 1112 0 1 2370
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1712256841
transform 1 0 1104 0 1 2370
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1712256841
transform 1 0 1096 0 1 2370
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1712256841
transform 1 0 1056 0 1 2370
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1712256841
transform 1 0 1048 0 1 2370
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1712256841
transform 1 0 1040 0 1 2370
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1712256841
transform 1 0 1032 0 1 2370
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1712256841
transform 1 0 992 0 1 2370
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1712256841
transform 1 0 984 0 1 2370
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1712256841
transform 1 0 976 0 1 2370
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1712256841
transform 1 0 872 0 1 2370
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1712256841
transform 1 0 864 0 1 2370
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1712256841
transform 1 0 760 0 1 2370
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1712256841
transform 1 0 752 0 1 2370
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1712256841
transform 1 0 648 0 1 2370
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1712256841
transform 1 0 640 0 1 2370
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1712256841
transform 1 0 536 0 1 2370
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1712256841
transform 1 0 528 0 1 2370
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1712256841
transform 1 0 424 0 1 2370
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1712256841
transform 1 0 416 0 1 2370
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1712256841
transform 1 0 312 0 1 2370
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1712256841
transform 1 0 304 0 1 2370
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1712256841
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1712256841
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1712256841
transform 1 0 184 0 1 2370
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1712256841
transform 1 0 80 0 1 2370
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1712256841
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1712256841
transform 1 0 3424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1712256841
transform 1 0 3416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1712256841
transform 1 0 3408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1712256841
transform 1 0 3352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1712256841
transform 1 0 3344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1712256841
transform 1 0 3304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1712256841
transform 1 0 3296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1712256841
transform 1 0 3288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1712256841
transform 1 0 3280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1712256841
transform 1 0 3224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1712256841
transform 1 0 3216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1712256841
transform 1 0 3208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1712256841
transform 1 0 3200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1712256841
transform 1 0 3192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1712256841
transform 1 0 3184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1712256841
transform 1 0 3176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1712256841
transform 1 0 3120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1712256841
transform 1 0 3112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1712256841
transform 1 0 3104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1712256841
transform 1 0 3096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1712256841
transform 1 0 3032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1712256841
transform 1 0 3024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1712256841
transform 1 0 3016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1712256841
transform 1 0 3008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1712256841
transform 1 0 3000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1712256841
transform 1 0 2960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1712256841
transform 1 0 2936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1712256841
transform 1 0 2928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1712256841
transform 1 0 2920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1712256841
transform 1 0 2912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1712256841
transform 1 0 2904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1712256841
transform 1 0 2896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1712256841
transform 1 0 2856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1712256841
transform 1 0 2848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1712256841
transform 1 0 2808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1712256841
transform 1 0 2800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1712256841
transform 1 0 2792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1712256841
transform 1 0 2784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1712256841
transform 1 0 2776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1712256841
transform 1 0 2736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1712256841
transform 1 0 2728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1712256841
transform 1 0 2688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1712256841
transform 1 0 2680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1712256841
transform 1 0 2672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1712256841
transform 1 0 2664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1712256841
transform 1 0 2656 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1712256841
transform 1 0 2592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1712256841
transform 1 0 2584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1712256841
transform 1 0 2576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1712256841
transform 1 0 2568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1712256841
transform 1 0 2528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1712256841
transform 1 0 2520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1712256841
transform 1 0 2512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1712256841
transform 1 0 2472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1712256841
transform 1 0 2464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1712256841
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1712256841
transform 1 0 2448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1712256841
transform 1 0 2408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1712256841
transform 1 0 2400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1712256841
transform 1 0 2392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1712256841
transform 1 0 2352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1712256841
transform 1 0 2344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1712256841
transform 1 0 2336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1712256841
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1712256841
transform 1 0 2288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1712256841
transform 1 0 2280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1712256841
transform 1 0 2272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1712256841
transform 1 0 2232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1712256841
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1712256841
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1712256841
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1712256841
transform 1 0 2168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1712256841
transform 1 0 2160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1712256841
transform 1 0 2152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1712256841
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1712256841
transform 1 0 2104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1712256841
transform 1 0 2096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1712256841
transform 1 0 2088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1712256841
transform 1 0 2048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1712256841
transform 1 0 2040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1712256841
transform 1 0 2032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1712256841
transform 1 0 2024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1712256841
transform 1 0 2016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1712256841
transform 1 0 1976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1712256841
transform 1 0 1968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1712256841
transform 1 0 1960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1712256841
transform 1 0 1920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1712256841
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1712256841
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1712256841
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1712256841
transform 1 0 1856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1712256841
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1712256841
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1712256841
transform 1 0 1832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1712256841
transform 1 0 1792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1712256841
transform 1 0 1784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1712256841
transform 1 0 1728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1712256841
transform 1 0 1720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1712256841
transform 1 0 1712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1712256841
transform 1 0 1704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1712256841
transform 1 0 1640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1712256841
transform 1 0 1632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1712256841
transform 1 0 1624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1712256841
transform 1 0 1616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1712256841
transform 1 0 1576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1712256841
transform 1 0 1568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1712256841
transform 1 0 1528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1712256841
transform 1 0 1520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1712256841
transform 1 0 1512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1712256841
transform 1 0 1504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1712256841
transform 1 0 1496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1712256841
transform 1 0 1424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1712256841
transform 1 0 1416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1712256841
transform 1 0 1408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1712256841
transform 1 0 1400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1712256841
transform 1 0 1392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1712256841
transform 1 0 1384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1712256841
transform 1 0 1376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1712256841
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1712256841
transform 1 0 1296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1712256841
transform 1 0 1288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1712256841
transform 1 0 1280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1712256841
transform 1 0 1272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1712256841
transform 1 0 1232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1712256841
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1712256841
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1712256841
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1712256841
transform 1 0 1168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1712256841
transform 1 0 1160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1712256841
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1712256841
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1712256841
transform 1 0 1072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1712256841
transform 1 0 1064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1712256841
transform 1 0 1056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1712256841
transform 1 0 1048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1712256841
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1712256841
transform 1 0 984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1712256841
transform 1 0 976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1712256841
transform 1 0 968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1712256841
transform 1 0 960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1712256841
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1712256841
transform 1 0 944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1712256841
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1712256841
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1712256841
transform 1 0 872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1712256841
transform 1 0 864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1712256841
transform 1 0 856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1712256841
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1712256841
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1712256841
transform 1 0 800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1712256841
transform 1 0 760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1712256841
transform 1 0 752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1712256841
transform 1 0 744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1712256841
transform 1 0 736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1712256841
transform 1 0 728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1712256841
transform 1 0 688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1712256841
transform 1 0 680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1712256841
transform 1 0 672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1712256841
transform 1 0 648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1712256841
transform 1 0 640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1712256841
transform 1 0 632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1712256841
transform 1 0 624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1712256841
transform 1 0 584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1712256841
transform 1 0 576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1712256841
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1712256841
transform 1 0 560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1712256841
transform 1 0 520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1712256841
transform 1 0 512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1712256841
transform 1 0 504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1712256841
transform 1 0 496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1712256841
transform 1 0 456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1712256841
transform 1 0 448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1712256841
transform 1 0 440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1712256841
transform 1 0 432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1712256841
transform 1 0 424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1712256841
transform 1 0 384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1712256841
transform 1 0 376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1712256841
transform 1 0 368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1712256841
transform 1 0 328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1712256841
transform 1 0 320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1712256841
transform 1 0 312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1712256841
transform 1 0 304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1712256841
transform 1 0 296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1712256841
transform 1 0 288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1712256841
transform 1 0 248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1712256841
transform 1 0 208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1712256841
transform 1 0 200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1712256841
transform 1 0 192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1712256841
transform 1 0 184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1712256841
transform 1 0 176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1712256841
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1712256841
transform 1 0 3424 0 1 2170
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1712256841
transform 1 0 3392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1712256841
transform 1 0 3384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1712256841
transform 1 0 3376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1712256841
transform 1 0 3368 0 1 2170
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1712256841
transform 1 0 3320 0 1 2170
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1712256841
transform 1 0 3312 0 1 2170
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1712256841
transform 1 0 3272 0 1 2170
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1712256841
transform 1 0 3264 0 1 2170
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1712256841
transform 1 0 3256 0 1 2170
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1712256841
transform 1 0 3184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1712256841
transform 1 0 3176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1712256841
transform 1 0 3152 0 1 2170
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1712256841
transform 1 0 3144 0 1 2170
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1712256841
transform 1 0 3136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1712256841
transform 1 0 3128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1712256841
transform 1 0 3064 0 1 2170
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1712256841
transform 1 0 3056 0 1 2170
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1712256841
transform 1 0 3048 0 1 2170
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1712256841
transform 1 0 3040 0 1 2170
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1712256841
transform 1 0 3000 0 1 2170
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1712256841
transform 1 0 2960 0 1 2170
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1712256841
transform 1 0 2952 0 1 2170
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1712256841
transform 1 0 2944 0 1 2170
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1712256841
transform 1 0 2936 0 1 2170
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1712256841
transform 1 0 2928 0 1 2170
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1712256841
transform 1 0 2888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1712256841
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1712256841
transform 1 0 2840 0 1 2170
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1712256841
transform 1 0 2832 0 1 2170
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1712256841
transform 1 0 2824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1712256841
transform 1 0 2816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1712256841
transform 1 0 2752 0 1 2170
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1712256841
transform 1 0 2744 0 1 2170
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1712256841
transform 1 0 2736 0 1 2170
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1712256841
transform 1 0 2696 0 1 2170
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1712256841
transform 1 0 2688 0 1 2170
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1712256841
transform 1 0 2680 0 1 2170
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1712256841
transform 1 0 2640 0 1 2170
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1712256841
transform 1 0 2632 0 1 2170
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1712256841
transform 1 0 2584 0 1 2170
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1712256841
transform 1 0 2576 0 1 2170
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1712256841
transform 1 0 2568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1712256841
transform 1 0 2560 0 1 2170
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1712256841
transform 1 0 2512 0 1 2170
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1712256841
transform 1 0 2504 0 1 2170
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1712256841
transform 1 0 2496 0 1 2170
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1712256841
transform 1 0 2472 0 1 2170
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1712256841
transform 1 0 2464 0 1 2170
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1712256841
transform 1 0 2456 0 1 2170
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1712256841
transform 1 0 2408 0 1 2170
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1712256841
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1712256841
transform 1 0 2392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1712256841
transform 1 0 2384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1712256841
transform 1 0 2376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1712256841
transform 1 0 2304 0 1 2170
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1712256841
transform 1 0 2296 0 1 2170
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1712256841
transform 1 0 2288 0 1 2170
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1712256841
transform 1 0 2280 0 1 2170
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1712256841
transform 1 0 2272 0 1 2170
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1712256841
transform 1 0 2240 0 1 2170
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1712256841
transform 1 0 2192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1712256841
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1712256841
transform 1 0 2176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1712256841
transform 1 0 2168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1712256841
transform 1 0 2160 0 1 2170
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1712256841
transform 1 0 2112 0 1 2170
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1712256841
transform 1 0 2104 0 1 2170
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1712256841
transform 1 0 2072 0 1 2170
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1712256841
transform 1 0 2064 0 1 2170
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1712256841
transform 1 0 2056 0 1 2170
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1712256841
transform 1 0 2048 0 1 2170
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1712256841
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1712256841
transform 1 0 1992 0 1 2170
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1712256841
transform 1 0 1984 0 1 2170
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1712256841
transform 1 0 1976 0 1 2170
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1712256841
transform 1 0 1944 0 1 2170
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1712256841
transform 1 0 1936 0 1 2170
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1712256841
transform 1 0 1888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1712256841
transform 1 0 1880 0 1 2170
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1712256841
transform 1 0 1872 0 1 2170
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1712256841
transform 1 0 1864 0 1 2170
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1712256841
transform 1 0 1856 0 1 2170
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1712256841
transform 1 0 1816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1712256841
transform 1 0 1808 0 1 2170
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1712256841
transform 1 0 1776 0 1 2170
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1712256841
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1712256841
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1712256841
transform 1 0 1712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1712256841
transform 1 0 1704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1712256841
transform 1 0 1680 0 1 2170
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1712256841
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1712256841
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1712256841
transform 1 0 1656 0 1 2170
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1712256841
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1712256841
transform 1 0 1584 0 1 2170
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1712256841
transform 1 0 1576 0 1 2170
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1712256841
transform 1 0 1568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1712256841
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1712256841
transform 1 0 1504 0 1 2170
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1712256841
transform 1 0 1496 0 1 2170
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1712256841
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1712256841
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1712256841
transform 1 0 1472 0 1 2170
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1712256841
transform 1 0 1448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1712256841
transform 1 0 1400 0 1 2170
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1712256841
transform 1 0 1392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1712256841
transform 1 0 1384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1712256841
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1712256841
transform 1 0 1344 0 1 2170
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1712256841
transform 1 0 1312 0 1 2170
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1712256841
transform 1 0 1272 0 1 2170
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1712256841
transform 1 0 1264 0 1 2170
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1712256841
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1712256841
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1712256841
transform 1 0 1200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1712256841
transform 1 0 1192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1712256841
transform 1 0 1184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1712256841
transform 1 0 1144 0 1 2170
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1712256841
transform 1 0 1136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1712256841
transform 1 0 1088 0 1 2170
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1712256841
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1712256841
transform 1 0 1072 0 1 2170
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1712256841
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1712256841
transform 1 0 1000 0 1 2170
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1712256841
transform 1 0 992 0 1 2170
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1712256841
transform 1 0 984 0 1 2170
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1712256841
transform 1 0 976 0 1 2170
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1712256841
transform 1 0 968 0 1 2170
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1712256841
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1712256841
transform 1 0 904 0 1 2170
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1712256841
transform 1 0 856 0 1 2170
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1712256841
transform 1 0 848 0 1 2170
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1712256841
transform 1 0 840 0 1 2170
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1712256841
transform 1 0 816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1712256841
transform 1 0 808 0 1 2170
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1712256841
transform 1 0 776 0 1 2170
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1712256841
transform 1 0 768 0 1 2170
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1712256841
transform 1 0 760 0 1 2170
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1712256841
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1712256841
transform 1 0 704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1712256841
transform 1 0 696 0 1 2170
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1712256841
transform 1 0 688 0 1 2170
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1712256841
transform 1 0 640 0 1 2170
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1712256841
transform 1 0 632 0 1 2170
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1712256841
transform 1 0 624 0 1 2170
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1712256841
transform 1 0 616 0 1 2170
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1712256841
transform 1 0 568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1712256841
transform 1 0 560 0 1 2170
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1712256841
transform 1 0 552 0 1 2170
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1712256841
transform 1 0 544 0 1 2170
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1712256841
transform 1 0 536 0 1 2170
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1712256841
transform 1 0 504 0 1 2170
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1712256841
transform 1 0 472 0 1 2170
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1712256841
transform 1 0 464 0 1 2170
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1712256841
transform 1 0 456 0 1 2170
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1712256841
transform 1 0 448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1712256841
transform 1 0 440 0 1 2170
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1712256841
transform 1 0 408 0 1 2170
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1712256841
transform 1 0 400 0 1 2170
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1712256841
transform 1 0 392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1712256841
transform 1 0 352 0 1 2170
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1712256841
transform 1 0 344 0 1 2170
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1712256841
transform 1 0 336 0 1 2170
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1712256841
transform 1 0 328 0 1 2170
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1712256841
transform 1 0 296 0 1 2170
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1712256841
transform 1 0 288 0 1 2170
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1712256841
transform 1 0 280 0 1 2170
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1712256841
transform 1 0 272 0 1 2170
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1712256841
transform 1 0 224 0 1 2170
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1712256841
transform 1 0 216 0 1 2170
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1712256841
transform 1 0 208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1712256841
transform 1 0 200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1712256841
transform 1 0 192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1712256841
transform 1 0 184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1712256841
transform 1 0 144 0 1 2170
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1712256841
transform 1 0 136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1712256841
transform 1 0 128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1712256841
transform 1 0 120 0 1 2170
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1712256841
transform 1 0 80 0 1 2170
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1712256841
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1712256841
transform 1 0 3424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1712256841
transform 1 0 3416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1712256841
transform 1 0 3344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1712256841
transform 1 0 3336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1712256841
transform 1 0 3272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1712256841
transform 1 0 3264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1712256841
transform 1 0 3224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1712256841
transform 1 0 3216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1712256841
transform 1 0 3208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1712256841
transform 1 0 3200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1712256841
transform 1 0 3112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1712256841
transform 1 0 3104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1712256841
transform 1 0 3096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1712256841
transform 1 0 3088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1712256841
transform 1 0 3080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1712256841
transform 1 0 3000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1712256841
transform 1 0 2992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1712256841
transform 1 0 2984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1712256841
transform 1 0 2976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1712256841
transform 1 0 2968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1712256841
transform 1 0 2896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1712256841
transform 1 0 2888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1712256841
transform 1 0 2848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1712256841
transform 1 0 2840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1712256841
transform 1 0 2808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1712256841
transform 1 0 2800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1712256841
transform 1 0 2792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1712256841
transform 1 0 2728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1712256841
transform 1 0 2720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1712256841
transform 1 0 2712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1712256841
transform 1 0 2704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1712256841
transform 1 0 2696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1712256841
transform 1 0 2616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1712256841
transform 1 0 2608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1712256841
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1712256841
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1712256841
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1712256841
transform 1 0 2536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1712256841
transform 1 0 2528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1712256841
transform 1 0 2488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1712256841
transform 1 0 2480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1712256841
transform 1 0 2472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1712256841
transform 1 0 2448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1712256841
transform 1 0 2408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1712256841
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1712256841
transform 1 0 2392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1712256841
transform 1 0 2384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1712256841
transform 1 0 2336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1712256841
transform 1 0 2312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1712256841
transform 1 0 2304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1712256841
transform 1 0 2296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1712256841
transform 1 0 2288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1712256841
transform 1 0 2280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1712256841
transform 1 0 2232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1712256841
transform 1 0 2224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1712256841
transform 1 0 2192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1712256841
transform 1 0 2184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1712256841
transform 1 0 2176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1712256841
transform 1 0 2168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1712256841
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1712256841
transform 1 0 2112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1712256841
transform 1 0 2104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1712256841
transform 1 0 2096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1712256841
transform 1 0 2056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1712256841
transform 1 0 2048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1712256841
transform 1 0 2040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1712256841
transform 1 0 2032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1712256841
transform 1 0 2024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1712256841
transform 1 0 1976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1712256841
transform 1 0 1968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1712256841
transform 1 0 1960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1712256841
transform 1 0 1952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1712256841
transform 1 0 1920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1712256841
transform 1 0 1888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1712256841
transform 1 0 1880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1712256841
transform 1 0 1872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1712256841
transform 1 0 1864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1712256841
transform 1 0 1856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1712256841
transform 1 0 1808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1712256841
transform 1 0 1800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1712256841
transform 1 0 1792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1712256841
transform 1 0 1760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1712256841
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1712256841
transform 1 0 1744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1712256841
transform 1 0 1704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1712256841
transform 1 0 1696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1712256841
transform 1 0 1688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1712256841
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1712256841
transform 1 0 1632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1712256841
transform 1 0 1624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1712256841
transform 1 0 1616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1712256841
transform 1 0 1608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1712256841
transform 1 0 1560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1712256841
transform 1 0 1552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1712256841
transform 1 0 1544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1712256841
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1712256841
transform 1 0 1488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1712256841
transform 1 0 1480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1712256841
transform 1 0 1472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1712256841
transform 1 0 1424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1712256841
transform 1 0 1416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1712256841
transform 1 0 1408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1712256841
transform 1 0 1400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1712256841
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1712256841
transform 1 0 1344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1712256841
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1712256841
transform 1 0 1304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1712256841
transform 1 0 1296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1712256841
transform 1 0 1288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1712256841
transform 1 0 1216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1712256841
transform 1 0 1208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1712256841
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1712256841
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1712256841
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1712256841
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1712256841
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1712256841
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1712256841
transform 1 0 1056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1712256841
transform 1 0 1048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1712256841
transform 1 0 1040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1712256841
transform 1 0 992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1712256841
transform 1 0 984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1712256841
transform 1 0 976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1712256841
transform 1 0 968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1712256841
transform 1 0 912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1712256841
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1712256841
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1712256841
transform 1 0 888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1712256841
transform 1 0 840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1712256841
transform 1 0 832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1712256841
transform 1 0 824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1712256841
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1712256841
transform 1 0 808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1712256841
transform 1 0 752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1712256841
transform 1 0 744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1712256841
transform 1 0 736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1712256841
transform 1 0 728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1712256841
transform 1 0 696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1712256841
transform 1 0 688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1712256841
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1712256841
transform 1 0 632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1712256841
transform 1 0 624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1712256841
transform 1 0 616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1712256841
transform 1 0 568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1712256841
transform 1 0 560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1712256841
transform 1 0 552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1712256841
transform 1 0 520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1712256841
transform 1 0 480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1712256841
transform 1 0 472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1712256841
transform 1 0 464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1712256841
transform 1 0 456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1712256841
transform 1 0 408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1712256841
transform 1 0 400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1712256841
transform 1 0 392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1712256841
transform 1 0 384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1712256841
transform 1 0 336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1712256841
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1712256841
transform 1 0 296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1712256841
transform 1 0 288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1712256841
transform 1 0 280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1712256841
transform 1 0 232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1712256841
transform 1 0 224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1712256841
transform 1 0 216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1712256841
transform 1 0 168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1712256841
transform 1 0 160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1712256841
transform 1 0 152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1712256841
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1712256841
transform 1 0 136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1712256841
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1712256841
transform 1 0 3424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1712256841
transform 1 0 3416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1712256841
transform 1 0 3408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1712256841
transform 1 0 3400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1712256841
transform 1 0 3392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1712256841
transform 1 0 3384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1712256841
transform 1 0 3376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1712256841
transform 1 0 3368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1712256841
transform 1 0 3360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1712256841
transform 1 0 3312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1712256841
transform 1 0 3304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1712256841
transform 1 0 3280 0 1 1970
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1712256841
transform 1 0 3272 0 1 1970
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1712256841
transform 1 0 3264 0 1 1970
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1712256841
transform 1 0 3256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1712256841
transform 1 0 3248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1712256841
transform 1 0 3192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1712256841
transform 1 0 3184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1712256841
transform 1 0 3176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1712256841
transform 1 0 3168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1712256841
transform 1 0 3160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1712256841
transform 1 0 3120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1712256841
transform 1 0 3112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1712256841
transform 1 0 3104 0 1 1970
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1712256841
transform 1 0 3056 0 1 1970
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1712256841
transform 1 0 3048 0 1 1970
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1712256841
transform 1 0 3040 0 1 1970
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1712256841
transform 1 0 3032 0 1 1970
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1712256841
transform 1 0 3024 0 1 1970
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1712256841
transform 1 0 2984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1712256841
transform 1 0 2976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1712256841
transform 1 0 2968 0 1 1970
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1712256841
transform 1 0 2960 0 1 1970
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1712256841
transform 1 0 2912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1712256841
transform 1 0 2904 0 1 1970
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1712256841
transform 1 0 2896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1712256841
transform 1 0 2888 0 1 1970
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1712256841
transform 1 0 2848 0 1 1970
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1712256841
transform 1 0 2840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1712256841
transform 1 0 2832 0 1 1970
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1712256841
transform 1 0 2792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1712256841
transform 1 0 2784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1712256841
transform 1 0 2776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1712256841
transform 1 0 2736 0 1 1970
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1712256841
transform 1 0 2728 0 1 1970
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1712256841
transform 1 0 2720 0 1 1970
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1712256841
transform 1 0 2712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1712256841
transform 1 0 2704 0 1 1970
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1712256841
transform 1 0 2640 0 1 1970
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1712256841
transform 1 0 2632 0 1 1970
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1712256841
transform 1 0 2624 0 1 1970
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1712256841
transform 1 0 2616 0 1 1970
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1712256841
transform 1 0 2608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1712256841
transform 1 0 2600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1712256841
transform 1 0 2544 0 1 1970
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1712256841
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1712256841
transform 1 0 2528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1712256841
transform 1 0 2496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1712256841
transform 1 0 2488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1712256841
transform 1 0 2448 0 1 1970
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1712256841
transform 1 0 2440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1712256841
transform 1 0 2432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1712256841
transform 1 0 2392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1712256841
transform 1 0 2384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1712256841
transform 1 0 2376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1712256841
transform 1 0 2368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1712256841
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1712256841
transform 1 0 2304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1712256841
transform 1 0 2296 0 1 1970
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1712256841
transform 1 0 2248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1712256841
transform 1 0 2240 0 1 1970
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1712256841
transform 1 0 2200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1712256841
transform 1 0 2192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1712256841
transform 1 0 2184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1712256841
transform 1 0 2176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1712256841
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1712256841
transform 1 0 2088 0 1 1970
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1712256841
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1712256841
transform 1 0 2072 0 1 1970
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1712256841
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1712256841
transform 1 0 2016 0 1 1970
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1712256841
transform 1 0 2008 0 1 1970
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1712256841
transform 1 0 1968 0 1 1970
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1712256841
transform 1 0 1960 0 1 1970
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1712256841
transform 1 0 1952 0 1 1970
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1712256841
transform 1 0 1912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1712256841
transform 1 0 1904 0 1 1970
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1712256841
transform 1 0 1872 0 1 1970
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1712256841
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1712256841
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1712256841
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1712256841
transform 1 0 1784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1712256841
transform 1 0 1776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1712256841
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1712256841
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1712256841
transform 1 0 1712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1712256841
transform 1 0 1704 0 1 1970
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1712256841
transform 1 0 1664 0 1 1970
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1712256841
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1712256841
transform 1 0 1648 0 1 1970
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1712256841
transform 1 0 1600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1712256841
transform 1 0 1592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1712256841
transform 1 0 1584 0 1 1970
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1712256841
transform 1 0 1528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1712256841
transform 1 0 1520 0 1 1970
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1712256841
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1712256841
transform 1 0 1488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1712256841
transform 1 0 1480 0 1 1970
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1712256841
transform 1 0 1416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1712256841
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1712256841
transform 1 0 1400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1712256841
transform 1 0 1392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1712256841
transform 1 0 1384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1712256841
transform 1 0 1336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1712256841
transform 1 0 1304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1712256841
transform 1 0 1296 0 1 1970
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1712256841
transform 1 0 1288 0 1 1970
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1712256841
transform 1 0 1280 0 1 1970
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1712256841
transform 1 0 1232 0 1 1970
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1712256841
transform 1 0 1224 0 1 1970
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1712256841
transform 1 0 1184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1712256841
transform 1 0 1176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1712256841
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1712256841
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1712256841
transform 1 0 1112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1712256841
transform 1 0 1080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1712256841
transform 1 0 1072 0 1 1970
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1712256841
transform 1 0 1064 0 1 1970
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1712256841
transform 1 0 1016 0 1 1970
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1712256841
transform 1 0 984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1712256841
transform 1 0 976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1712256841
transform 1 0 968 0 1 1970
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1712256841
transform 1 0 960 0 1 1970
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1712256841
transform 1 0 880 0 1 1970
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1712256841
transform 1 0 872 0 1 1970
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1712256841
transform 1 0 864 0 1 1970
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1712256841
transform 1 0 824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1712256841
transform 1 0 816 0 1 1970
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1712256841
transform 1 0 768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1712256841
transform 1 0 760 0 1 1970
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1712256841
transform 1 0 752 0 1 1970
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1712256841
transform 1 0 712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1712256841
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1712256841
transform 1 0 696 0 1 1970
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1712256841
transform 1 0 648 0 1 1970
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1712256841
transform 1 0 640 0 1 1970
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1712256841
transform 1 0 632 0 1 1970
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1712256841
transform 1 0 600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1712256841
transform 1 0 592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1712256841
transform 1 0 584 0 1 1970
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1712256841
transform 1 0 544 0 1 1970
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1712256841
transform 1 0 536 0 1 1970
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1712256841
transform 1 0 504 0 1 1970
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1712256841
transform 1 0 496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1712256841
transform 1 0 488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1712256841
transform 1 0 448 0 1 1970
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1712256841
transform 1 0 440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1712256841
transform 1 0 392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1712256841
transform 1 0 384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1712256841
transform 1 0 376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1712256841
transform 1 0 368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1712256841
transform 1 0 328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1712256841
transform 1 0 320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1712256841
transform 1 0 288 0 1 1970
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1712256841
transform 1 0 280 0 1 1970
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1712256841
transform 1 0 272 0 1 1970
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1712256841
transform 1 0 264 0 1 1970
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1712256841
transform 1 0 224 0 1 1970
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1712256841
transform 1 0 192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1712256841
transform 1 0 184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1712256841
transform 1 0 176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1712256841
transform 1 0 168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1712256841
transform 1 0 136 0 1 1970
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1712256841
transform 1 0 128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1712256841
transform 1 0 80 0 1 1970
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1712256841
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1712256841
transform 1 0 3328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1712256841
transform 1 0 3320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1712256841
transform 1 0 3312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1712256841
transform 1 0 3256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1712256841
transform 1 0 3248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1712256841
transform 1 0 3240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1712256841
transform 1 0 3168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1712256841
transform 1 0 3160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1712256841
transform 1 0 3128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1712256841
transform 1 0 3120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1712256841
transform 1 0 3112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1712256841
transform 1 0 3072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1712256841
transform 1 0 3064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1712256841
transform 1 0 3056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1712256841
transform 1 0 3048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1712256841
transform 1 0 3040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1712256841
transform 1 0 3000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1712256841
transform 1 0 2960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1712256841
transform 1 0 2952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1712256841
transform 1 0 2944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1712256841
transform 1 0 2936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1712256841
transform 1 0 2928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1712256841
transform 1 0 2904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1712256841
transform 1 0 2864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1712256841
transform 1 0 2856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1712256841
transform 1 0 2848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1712256841
transform 1 0 2840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1712256841
transform 1 0 2808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1712256841
transform 1 0 2784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1712256841
transform 1 0 2744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1712256841
transform 1 0 2736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1712256841
transform 1 0 2712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1712256841
transform 1 0 2704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1712256841
transform 1 0 2696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1712256841
transform 1 0 2656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1712256841
transform 1 0 2648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1712256841
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1712256841
transform 1 0 2576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1712256841
transform 1 0 2568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1712256841
transform 1 0 2560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1712256841
transform 1 0 2520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1712256841
transform 1 0 2512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1712256841
transform 1 0 2464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1712256841
transform 1 0 2456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1712256841
transform 1 0 2448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1712256841
transform 1 0 2440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1712256841
transform 1 0 2432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1712256841
transform 1 0 2360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1712256841
transform 1 0 2352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1712256841
transform 1 0 2344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1712256841
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1712256841
transform 1 0 2328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1712256841
transform 1 0 2304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1712256841
transform 1 0 2296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1712256841
transform 1 0 2232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1712256841
transform 1 0 2224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1712256841
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1712256841
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1712256841
transform 1 0 2136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1712256841
transform 1 0 2128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1712256841
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1712256841
transform 1 0 2112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1712256841
transform 1 0 2104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1712256841
transform 1 0 2096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1712256841
transform 1 0 2024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1712256841
transform 1 0 2016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1712256841
transform 1 0 2008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1712256841
transform 1 0 2000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1712256841
transform 1 0 1960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1712256841
transform 1 0 1952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1712256841
transform 1 0 1920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1712256841
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1712256841
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1712256841
transform 1 0 1856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1712256841
transform 1 0 1848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1712256841
transform 1 0 1840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1712256841
transform 1 0 1832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1712256841
transform 1 0 1768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1712256841
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1712256841
transform 1 0 1728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1712256841
transform 1 0 1720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1712256841
transform 1 0 1712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1712256841
transform 1 0 1704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1712256841
transform 1 0 1640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1712256841
transform 1 0 1632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1712256841
transform 1 0 1624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1712256841
transform 1 0 1616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1712256841
transform 1 0 1608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1712256841
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1712256841
transform 1 0 1528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1712256841
transform 1 0 1520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1712256841
transform 1 0 1512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1712256841
transform 1 0 1504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1712256841
transform 1 0 1496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1712256841
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1712256841
transform 1 0 1440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1712256841
transform 1 0 1400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1712256841
transform 1 0 1392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1712256841
transform 1 0 1384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1712256841
transform 1 0 1376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1712256841
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1712256841
transform 1 0 1336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1712256841
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1712256841
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1712256841
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1712256841
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1712256841
transform 1 0 1256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1712256841
transform 1 0 1248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1712256841
transform 1 0 1192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1712256841
transform 1 0 1184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1712256841
transform 1 0 1176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1712256841
transform 1 0 1168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1712256841
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1712256841
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1712256841
transform 1 0 1096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1712256841
transform 1 0 1088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1712256841
transform 1 0 1056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1712256841
transform 1 0 1048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1712256841
transform 1 0 1000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1712256841
transform 1 0 992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1712256841
transform 1 0 984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1712256841
transform 1 0 976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1712256841
transform 1 0 928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1712256841
transform 1 0 920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1712256841
transform 1 0 912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1712256841
transform 1 0 872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1712256841
transform 1 0 864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1712256841
transform 1 0 856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1712256841
transform 1 0 816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1712256841
transform 1 0 808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1712256841
transform 1 0 800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1712256841
transform 1 0 760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1712256841
transform 1 0 752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1712256841
transform 1 0 744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1712256841
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1712256841
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1712256841
transform 1 0 688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1712256841
transform 1 0 664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1712256841
transform 1 0 656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1712256841
transform 1 0 616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1712256841
transform 1 0 608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1712256841
transform 1 0 600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1712256841
transform 1 0 592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1712256841
transform 1 0 544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1712256841
transform 1 0 536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1712256841
transform 1 0 528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1712256841
transform 1 0 496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1712256841
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1712256841
transform 1 0 464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1712256841
transform 1 0 456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1712256841
transform 1 0 448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1712256841
transform 1 0 400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1712256841
transform 1 0 392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1712256841
transform 1 0 384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1712256841
transform 1 0 336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1712256841
transform 1 0 328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1712256841
transform 1 0 320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1712256841
transform 1 0 280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1712256841
transform 1 0 272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1712256841
transform 1 0 264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1712256841
transform 1 0 224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1712256841
transform 1 0 216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1712256841
transform 1 0 208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1712256841
transform 1 0 160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1712256841
transform 1 0 152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1712256841
transform 1 0 144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1712256841
transform 1 0 136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1712256841
transform 1 0 128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1712256841
transform 1 0 80 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1712256841
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1712256841
transform 1 0 3424 0 1 1770
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1712256841
transform 1 0 3416 0 1 1770
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1712256841
transform 1 0 3408 0 1 1770
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1712256841
transform 1 0 3400 0 1 1770
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1712256841
transform 1 0 3392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1712256841
transform 1 0 3384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1712256841
transform 1 0 3376 0 1 1770
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1712256841
transform 1 0 3368 0 1 1770
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1712256841
transform 1 0 3360 0 1 1770
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1712256841
transform 1 0 3352 0 1 1770
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1712256841
transform 1 0 3344 0 1 1770
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1712256841
transform 1 0 3336 0 1 1770
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1712256841
transform 1 0 3328 0 1 1770
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1712256841
transform 1 0 3280 0 1 1770
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1712256841
transform 1 0 3272 0 1 1770
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1712256841
transform 1 0 3264 0 1 1770
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1712256841
transform 1 0 3232 0 1 1770
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1712256841
transform 1 0 3224 0 1 1770
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1712256841
transform 1 0 3216 0 1 1770
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1712256841
transform 1 0 3208 0 1 1770
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1712256841
transform 1 0 3200 0 1 1770
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1712256841
transform 1 0 3168 0 1 1770
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1712256841
transform 1 0 3160 0 1 1770
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1712256841
transform 1 0 3120 0 1 1770
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1712256841
transform 1 0 3112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1712256841
transform 1 0 3104 0 1 1770
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1712256841
transform 1 0 3096 0 1 1770
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1712256841
transform 1 0 3072 0 1 1770
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1712256841
transform 1 0 3064 0 1 1770
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1712256841
transform 1 0 3024 0 1 1770
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1712256841
transform 1 0 3016 0 1 1770
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1712256841
transform 1 0 3008 0 1 1770
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1712256841
transform 1 0 3000 0 1 1770
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1712256841
transform 1 0 2992 0 1 1770
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1712256841
transform 1 0 2944 0 1 1770
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1712256841
transform 1 0 2936 0 1 1770
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1712256841
transform 1 0 2928 0 1 1770
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1712256841
transform 1 0 2920 0 1 1770
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1712256841
transform 1 0 2896 0 1 1770
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1712256841
transform 1 0 2888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1712256841
transform 1 0 2880 0 1 1770
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1712256841
transform 1 0 2872 0 1 1770
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1712256841
transform 1 0 2824 0 1 1770
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1712256841
transform 1 0 2816 0 1 1770
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1712256841
transform 1 0 2808 0 1 1770
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1712256841
transform 1 0 2800 0 1 1770
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1712256841
transform 1 0 2792 0 1 1770
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1712256841
transform 1 0 2744 0 1 1770
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1712256841
transform 1 0 2736 0 1 1770
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1712256841
transform 1 0 2728 0 1 1770
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1712256841
transform 1 0 2720 0 1 1770
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1712256841
transform 1 0 2712 0 1 1770
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1712256841
transform 1 0 2672 0 1 1770
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1712256841
transform 1 0 2664 0 1 1770
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1712256841
transform 1 0 2656 0 1 1770
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1712256841
transform 1 0 2648 0 1 1770
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1712256841
transform 1 0 2640 0 1 1770
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1712256841
transform 1 0 2592 0 1 1770
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1712256841
transform 1 0 2584 0 1 1770
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1712256841
transform 1 0 2576 0 1 1770
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1712256841
transform 1 0 2568 0 1 1770
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1712256841
transform 1 0 2544 0 1 1770
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1712256841
transform 1 0 2512 0 1 1770
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1712256841
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1712256841
transform 1 0 2496 0 1 1770
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1712256841
transform 1 0 2488 0 1 1770
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1712256841
transform 1 0 2480 0 1 1770
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1712256841
transform 1 0 2440 0 1 1770
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1712256841
transform 1 0 2432 0 1 1770
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1712256841
transform 1 0 2400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1712256841
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1712256841
transform 1 0 2384 0 1 1770
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1712256841
transform 1 0 2352 0 1 1770
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1712256841
transform 1 0 2344 0 1 1770
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1712256841
transform 1 0 2336 0 1 1770
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1712256841
transform 1 0 2328 0 1 1770
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1712256841
transform 1 0 2280 0 1 1770
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1712256841
transform 1 0 2272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1712256841
transform 1 0 2264 0 1 1770
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1712256841
transform 1 0 2216 0 1 1770
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1712256841
transform 1 0 2208 0 1 1770
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1712256841
transform 1 0 2200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1712256841
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1712256841
transform 1 0 2184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1712256841
transform 1 0 2136 0 1 1770
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1712256841
transform 1 0 2128 0 1 1770
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1712256841
transform 1 0 2120 0 1 1770
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1712256841
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1712256841
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1712256841
transform 1 0 2056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1712256841
transform 1 0 2048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1712256841
transform 1 0 2016 0 1 1770
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1712256841
transform 1 0 2008 0 1 1770
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1712256841
transform 1 0 2000 0 1 1770
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1712256841
transform 1 0 1992 0 1 1770
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1712256841
transform 1 0 1936 0 1 1770
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1712256841
transform 1 0 1928 0 1 1770
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1712256841
transform 1 0 1920 0 1 1770
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1712256841
transform 1 0 1912 0 1 1770
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1712256841
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1712256841
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1712256841
transform 1 0 1856 0 1 1770
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1712256841
transform 1 0 1808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1712256841
transform 1 0 1800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1712256841
transform 1 0 1792 0 1 1770
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1712256841
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1712256841
transform 1 0 1720 0 1 1770
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1712256841
transform 1 0 1688 0 1 1770
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1712256841
transform 1 0 1640 0 1 1770
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1712256841
transform 1 0 1632 0 1 1770
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1712256841
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1712256841
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1712256841
transform 1 0 1568 0 1 1770
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1712256841
transform 1 0 1560 0 1 1770
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1712256841
transform 1 0 1520 0 1 1770
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1712256841
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1712256841
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1712256841
transform 1 0 1496 0 1 1770
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1712256841
transform 1 0 1416 0 1 1770
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1712256841
transform 1 0 1408 0 1 1770
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1712256841
transform 1 0 1400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1712256841
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1712256841
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1712256841
transform 1 0 1320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1712256841
transform 1 0 1280 0 1 1770
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1712256841
transform 1 0 1272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1712256841
transform 1 0 1264 0 1 1770
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1712256841
transform 1 0 1200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1712256841
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1712256841
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1712256841
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1712256841
transform 1 0 1168 0 1 1770
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1712256841
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1712256841
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1712256841
transform 1 0 1072 0 1 1770
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1712256841
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1712256841
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1712256841
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1712256841
transform 1 0 1000 0 1 1770
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1712256841
transform 1 0 992 0 1 1770
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1712256841
transform 1 0 984 0 1 1770
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1712256841
transform 1 0 944 0 1 1770
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1712256841
transform 1 0 936 0 1 1770
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1712256841
transform 1 0 928 0 1 1770
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1712256841
transform 1 0 920 0 1 1770
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1712256841
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1712256841
transform 1 0 856 0 1 1770
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1712256841
transform 1 0 848 0 1 1770
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1712256841
transform 1 0 824 0 1 1770
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1712256841
transform 1 0 816 0 1 1770
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1712256841
transform 1 0 808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1712256841
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1712256841
transform 1 0 744 0 1 1770
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1712256841
transform 1 0 736 0 1 1770
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1712256841
transform 1 0 728 0 1 1770
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1712256841
transform 1 0 720 0 1 1770
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1712256841
transform 1 0 712 0 1 1770
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1712256841
transform 1 0 664 0 1 1770
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1712256841
transform 1 0 656 0 1 1770
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1712256841
transform 1 0 648 0 1 1770
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1712256841
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1712256841
transform 1 0 600 0 1 1770
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1712256841
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1712256841
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1712256841
transform 1 0 536 0 1 1770
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1712256841
transform 1 0 528 0 1 1770
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1712256841
transform 1 0 520 0 1 1770
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1712256841
transform 1 0 512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1712256841
transform 1 0 504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1712256841
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1712256841
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1712256841
transform 1 0 440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1712256841
transform 1 0 432 0 1 1770
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1712256841
transform 1 0 424 0 1 1770
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1712256841
transform 1 0 376 0 1 1770
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1712256841
transform 1 0 368 0 1 1770
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1712256841
transform 1 0 360 0 1 1770
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1712256841
transform 1 0 352 0 1 1770
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1712256841
transform 1 0 344 0 1 1770
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1712256841
transform 1 0 312 0 1 1770
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1712256841
transform 1 0 304 0 1 1770
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1712256841
transform 1 0 272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1712256841
transform 1 0 264 0 1 1770
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1712256841
transform 1 0 256 0 1 1770
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1712256841
transform 1 0 248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1712256841
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1712256841
transform 1 0 200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1712256841
transform 1 0 192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1712256841
transform 1 0 184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1712256841
transform 1 0 176 0 1 1770
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1712256841
transform 1 0 144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1712256841
transform 1 0 136 0 1 1770
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1712256841
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1712256841
transform 1 0 88 0 1 1770
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1712256841
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1712256841
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1712256841
transform 1 0 3328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1712256841
transform 1 0 3320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1712256841
transform 1 0 3312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1712256841
transform 1 0 3304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1712256841
transform 1 0 3256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1712256841
transform 1 0 3248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1712256841
transform 1 0 3208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1712256841
transform 1 0 3200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1712256841
transform 1 0 3192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1712256841
transform 1 0 3128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1712256841
transform 1 0 3120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1712256841
transform 1 0 3112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1712256841
transform 1 0 3104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1712256841
transform 1 0 3056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1712256841
transform 1 0 3048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1712256841
transform 1 0 3040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1712256841
transform 1 0 3000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1712256841
transform 1 0 2992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1712256841
transform 1 0 2984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1712256841
transform 1 0 2936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1712256841
transform 1 0 2928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1712256841
transform 1 0 2920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1712256841
transform 1 0 2880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1712256841
transform 1 0 2872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1712256841
transform 1 0 2864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1712256841
transform 1 0 2824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1712256841
transform 1 0 2816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1712256841
transform 1 0 2792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1712256841
transform 1 0 2784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1712256841
transform 1 0 2760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1712256841
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1712256841
transform 1 0 2696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1712256841
transform 1 0 2688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1712256841
transform 1 0 2680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1712256841
transform 1 0 2624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1712256841
transform 1 0 2616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1712256841
transform 1 0 2608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1712256841
transform 1 0 2600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1712256841
transform 1 0 2592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1712256841
transform 1 0 2520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1712256841
transform 1 0 2512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1712256841
transform 1 0 2504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1712256841
transform 1 0 2496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1712256841
transform 1 0 2488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1712256841
transform 1 0 2480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1712256841
transform 1 0 2432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1712256841
transform 1 0 2424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1712256841
transform 1 0 2376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1712256841
transform 1 0 2368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1712256841
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1712256841
transform 1 0 2352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1712256841
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1712256841
transform 1 0 2296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1712256841
transform 1 0 2264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1712256841
transform 1 0 2256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1712256841
transform 1 0 2248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1712256841
transform 1 0 2200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1712256841
transform 1 0 2192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1712256841
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1712256841
transform 1 0 2176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1712256841
transform 1 0 2144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1712256841
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1712256841
transform 1 0 2104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1712256841
transform 1 0 2072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1712256841
transform 1 0 2064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1712256841
transform 1 0 2056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1712256841
transform 1 0 2048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1712256841
transform 1 0 2000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1712256841
transform 1 0 1992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1712256841
transform 1 0 1952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1712256841
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1712256841
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1712256841
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1712256841
transform 1 0 1872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1712256841
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1712256841
transform 1 0 1856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1712256841
transform 1 0 1848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1712256841
transform 1 0 1800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1712256841
transform 1 0 1792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1712256841
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1712256841
transform 1 0 1752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1712256841
transform 1 0 1744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1712256841
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1712256841
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1712256841
transform 1 0 1656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1712256841
transform 1 0 1648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1712256841
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1712256841
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1712256841
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1712256841
transform 1 0 1560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1712256841
transform 1 0 1552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1712256841
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1712256841
transform 1 0 1536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1712256841
transform 1 0 1496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1712256841
transform 1 0 1488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1712256841
transform 1 0 1480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1712256841
transform 1 0 1440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1712256841
transform 1 0 1432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1712256841
transform 1 0 1424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1712256841
transform 1 0 1416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1712256841
transform 1 0 1376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1712256841
transform 1 0 1368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1712256841
transform 1 0 1360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1712256841
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1712256841
transform 1 0 1312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1712256841
transform 1 0 1304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1712256841
transform 1 0 1296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1712256841
transform 1 0 1288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1712256841
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1712256841
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1712256841
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1712256841
transform 1 0 1224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1712256841
transform 1 0 1216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1712256841
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1712256841
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1712256841
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1712256841
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1712256841
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1712256841
transform 1 0 1104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1712256841
transform 1 0 1080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1712256841
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1712256841
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1712256841
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1712256841
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1712256841
transform 1 0 1000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1712256841
transform 1 0 992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1712256841
transform 1 0 984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1712256841
transform 1 0 976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1712256841
transform 1 0 968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1712256841
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1712256841
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1712256841
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1712256841
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1712256841
transform 1 0 864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1712256841
transform 1 0 856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1712256841
transform 1 0 848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1712256841
transform 1 0 808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1712256841
transform 1 0 800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1712256841
transform 1 0 792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1712256841
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1712256841
transform 1 0 760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1712256841
transform 1 0 752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1712256841
transform 1 0 744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1712256841
transform 1 0 704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1712256841
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1712256841
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1712256841
transform 1 0 680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1712256841
transform 1 0 648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1712256841
transform 1 0 640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1712256841
transform 1 0 632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1712256841
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1712256841
transform 1 0 584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1712256841
transform 1 0 576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1712256841
transform 1 0 568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1712256841
transform 1 0 536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1712256841
transform 1 0 528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1712256841
transform 1 0 520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1712256841
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1712256841
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1712256841
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1712256841
transform 1 0 440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1712256841
transform 1 0 432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1712256841
transform 1 0 424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1712256841
transform 1 0 416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1712256841
transform 1 0 384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1712256841
transform 1 0 360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1712256841
transform 1 0 352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1712256841
transform 1 0 344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1712256841
transform 1 0 336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1712256841
transform 1 0 328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1712256841
transform 1 0 320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1712256841
transform 1 0 264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1712256841
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1712256841
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1712256841
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1712256841
transform 1 0 232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1712256841
transform 1 0 224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1712256841
transform 1 0 168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1712256841
transform 1 0 160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1712256841
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1712256841
transform 1 0 144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1712256841
transform 1 0 136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1712256841
transform 1 0 128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1712256841
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1712256841
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1712256841
transform 1 0 3328 0 1 1570
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1712256841
transform 1 0 3320 0 1 1570
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1712256841
transform 1 0 3272 0 1 1570
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1712256841
transform 1 0 3264 0 1 1570
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1712256841
transform 1 0 3160 0 1 1570
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1712256841
transform 1 0 3152 0 1 1570
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1712256841
transform 1 0 3120 0 1 1570
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1712256841
transform 1 0 3072 0 1 1570
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1712256841
transform 1 0 3064 0 1 1570
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1712256841
transform 1 0 3040 0 1 1570
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1712256841
transform 1 0 3032 0 1 1570
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1712256841
transform 1 0 3024 0 1 1570
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1712256841
transform 1 0 3016 0 1 1570
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1712256841
transform 1 0 2968 0 1 1570
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1712256841
transform 1 0 2944 0 1 1570
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1712256841
transform 1 0 2936 0 1 1570
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1712256841
transform 1 0 2928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1712256841
transform 1 0 2920 0 1 1570
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1712256841
transform 1 0 2880 0 1 1570
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1712256841
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1712256841
transform 1 0 2840 0 1 1570
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1712256841
transform 1 0 2800 0 1 1570
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1712256841
transform 1 0 2792 0 1 1570
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1712256841
transform 1 0 2784 0 1 1570
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1712256841
transform 1 0 2776 0 1 1570
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1712256841
transform 1 0 2744 0 1 1570
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1712256841
transform 1 0 2712 0 1 1570
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1712256841
transform 1 0 2704 0 1 1570
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1712256841
transform 1 0 2696 0 1 1570
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1712256841
transform 1 0 2656 0 1 1570
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1712256841
transform 1 0 2648 0 1 1570
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1712256841
transform 1 0 2616 0 1 1570
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1712256841
transform 1 0 2608 0 1 1570
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1712256841
transform 1 0 2568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1712256841
transform 1 0 2560 0 1 1570
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1712256841
transform 1 0 2552 0 1 1570
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1712256841
transform 1 0 2544 0 1 1570
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1712256841
transform 1 0 2488 0 1 1570
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1712256841
transform 1 0 2480 0 1 1570
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1712256841
transform 1 0 2472 0 1 1570
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1712256841
transform 1 0 2448 0 1 1570
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1712256841
transform 1 0 2440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1712256841
transform 1 0 2400 0 1 1570
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1712256841
transform 1 0 2392 0 1 1570
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1712256841
transform 1 0 2384 0 1 1570
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1712256841
transform 1 0 2344 0 1 1570
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1712256841
transform 1 0 2336 0 1 1570
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1712256841
transform 1 0 2296 0 1 1570
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1712256841
transform 1 0 2288 0 1 1570
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1712256841
transform 1 0 2280 0 1 1570
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1712256841
transform 1 0 2272 0 1 1570
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1712256841
transform 1 0 2216 0 1 1570
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1712256841
transform 1 0 2208 0 1 1570
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1712256841
transform 1 0 2200 0 1 1570
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1712256841
transform 1 0 2192 0 1 1570
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1712256841
transform 1 0 2184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1712256841
transform 1 0 2128 0 1 1570
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1712256841
transform 1 0 2120 0 1 1570
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1712256841
transform 1 0 2112 0 1 1570
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1712256841
transform 1 0 2104 0 1 1570
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1712256841
transform 1 0 2096 0 1 1570
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1712256841
transform 1 0 2048 0 1 1570
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1712256841
transform 1 0 2040 0 1 1570
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1712256841
transform 1 0 1992 0 1 1570
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1712256841
transform 1 0 1984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1712256841
transform 1 0 1976 0 1 1570
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1712256841
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1712256841
transform 1 0 1928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1712256841
transform 1 0 1920 0 1 1570
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1712256841
transform 1 0 1872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1712256841
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1712256841
transform 1 0 1856 0 1 1570
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1712256841
transform 1 0 1824 0 1 1570
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1712256841
transform 1 0 1816 0 1 1570
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1712256841
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1712256841
transform 1 0 1760 0 1 1570
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1712256841
transform 1 0 1752 0 1 1570
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1712256841
transform 1 0 1744 0 1 1570
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1712256841
transform 1 0 1704 0 1 1570
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1712256841
transform 1 0 1696 0 1 1570
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1712256841
transform 1 0 1656 0 1 1570
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1712256841
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1712256841
transform 1 0 1640 0 1 1570
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1712256841
transform 1 0 1632 0 1 1570
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1712256841
transform 1 0 1584 0 1 1570
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1712256841
transform 1 0 1576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1712256841
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1712256841
transform 1 0 1528 0 1 1570
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1712256841
transform 1 0 1520 0 1 1570
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1712256841
transform 1 0 1512 0 1 1570
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1712256841
transform 1 0 1464 0 1 1570
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1712256841
transform 1 0 1456 0 1 1570
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1712256841
transform 1 0 1448 0 1 1570
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1712256841
transform 1 0 1408 0 1 1570
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1712256841
transform 1 0 1400 0 1 1570
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1712256841
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1712256841
transform 1 0 1384 0 1 1570
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1712256841
transform 1 0 1312 0 1 1570
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1712256841
transform 1 0 1304 0 1 1570
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1712256841
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1712256841
transform 1 0 1288 0 1 1570
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1712256841
transform 1 0 1280 0 1 1570
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1712256841
transform 1 0 1232 0 1 1570
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1712256841
transform 1 0 1224 0 1 1570
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1712256841
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1712256841
transform 1 0 1176 0 1 1570
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1712256841
transform 1 0 1168 0 1 1570
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1712256841
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1712256841
transform 1 0 1128 0 1 1570
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1712256841
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1712256841
transform 1 0 1064 0 1 1570
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1712256841
transform 1 0 1056 0 1 1570
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1712256841
transform 1 0 1048 0 1 1570
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1712256841
transform 1 0 1040 0 1 1570
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1712256841
transform 1 0 1032 0 1 1570
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1712256841
transform 1 0 960 0 1 1570
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1712256841
transform 1 0 952 0 1 1570
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1712256841
transform 1 0 944 0 1 1570
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1712256841
transform 1 0 936 0 1 1570
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1712256841
transform 1 0 928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1712256841
transform 1 0 864 0 1 1570
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1712256841
transform 1 0 856 0 1 1570
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1712256841
transform 1 0 848 0 1 1570
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1712256841
transform 1 0 840 0 1 1570
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1712256841
transform 1 0 808 0 1 1570
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1712256841
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1712256841
transform 1 0 744 0 1 1570
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1712256841
transform 1 0 736 0 1 1570
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1712256841
transform 1 0 728 0 1 1570
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1712256841
transform 1 0 720 0 1 1570
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1712256841
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1712256841
transform 1 0 640 0 1 1570
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1712256841
transform 1 0 632 0 1 1570
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1712256841
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1712256841
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1712256841
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1712256841
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1712256841
transform 1 0 544 0 1 1570
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1712256841
transform 1 0 536 0 1 1570
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1712256841
transform 1 0 528 0 1 1570
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1712256841
transform 1 0 472 0 1 1570
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1712256841
transform 1 0 464 0 1 1570
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1712256841
transform 1 0 456 0 1 1570
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1712256841
transform 1 0 408 0 1 1570
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1712256841
transform 1 0 400 0 1 1570
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1712256841
transform 1 0 360 0 1 1570
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1712256841
transform 1 0 352 0 1 1570
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1712256841
transform 1 0 344 0 1 1570
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1712256841
transform 1 0 336 0 1 1570
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1712256841
transform 1 0 264 0 1 1570
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1712256841
transform 1 0 256 0 1 1570
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1712256841
transform 1 0 248 0 1 1570
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1712256841
transform 1 0 240 0 1 1570
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1712256841
transform 1 0 232 0 1 1570
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1712256841
transform 1 0 184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1712256841
transform 1 0 152 0 1 1570
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1712256841
transform 1 0 144 0 1 1570
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1712256841
transform 1 0 136 0 1 1570
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1712256841
transform 1 0 128 0 1 1570
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1712256841
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1712256841
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1712256841
transform 1 0 3424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1712256841
transform 1 0 3416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1712256841
transform 1 0 3408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1712256841
transform 1 0 3328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1712256841
transform 1 0 3320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1712256841
transform 1 0 3312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1712256841
transform 1 0 3304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1712256841
transform 1 0 3232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1712256841
transform 1 0 3224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1712256841
transform 1 0 3216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1712256841
transform 1 0 3112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1712256841
transform 1 0 3104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1712256841
transform 1 0 3096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1712256841
transform 1 0 3088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1712256841
transform 1 0 3024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1712256841
transform 1 0 3016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1712256841
transform 1 0 3008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1712256841
transform 1 0 3000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1712256841
transform 1 0 2992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1712256841
transform 1 0 2952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1712256841
transform 1 0 2912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1712256841
transform 1 0 2904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1712256841
transform 1 0 2896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1712256841
transform 1 0 2888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1712256841
transform 1 0 2880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1712256841
transform 1 0 2840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1712256841
transform 1 0 2800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1712256841
transform 1 0 2792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1712256841
transform 1 0 2784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1712256841
transform 1 0 2776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1712256841
transform 1 0 2768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1712256841
transform 1 0 2712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1712256841
transform 1 0 2704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1712256841
transform 1 0 2696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1712256841
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1712256841
transform 1 0 2680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1712256841
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1712256841
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1712256841
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1712256841
transform 1 0 2584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1712256841
transform 1 0 2576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1712256841
transform 1 0 2568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1712256841
transform 1 0 2560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1712256841
transform 1 0 2528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1712256841
transform 1 0 2496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1712256841
transform 1 0 2488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1712256841
transform 1 0 2480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1712256841
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1712256841
transform 1 0 2432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1712256841
transform 1 0 2424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1712256841
transform 1 0 2400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1712256841
transform 1 0 2392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1712256841
transform 1 0 2384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1712256841
transform 1 0 2376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1712256841
transform 1 0 2336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1712256841
transform 1 0 2304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1712256841
transform 1 0 2296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1712256841
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1712256841
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1712256841
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1712256841
transform 1 0 2224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1712256841
transform 1 0 2216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1712256841
transform 1 0 2208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1712256841
transform 1 0 2168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1712256841
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1712256841
transform 1 0 2152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1712256841
transform 1 0 2144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1712256841
transform 1 0 2112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1712256841
transform 1 0 2104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1712256841
transform 1 0 2056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1712256841
transform 1 0 2048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1712256841
transform 1 0 2040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1712256841
transform 1 0 2032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1712256841
transform 1 0 2024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1712256841
transform 1 0 1976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1712256841
transform 1 0 1968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1712256841
transform 1 0 1960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1712256841
transform 1 0 1920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1712256841
transform 1 0 1912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1712256841
transform 1 0 1888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1712256841
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1712256841
transform 1 0 1848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1712256841
transform 1 0 1840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1712256841
transform 1 0 1832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1712256841
transform 1 0 1824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1712256841
transform 1 0 1792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1712256841
transform 1 0 1752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1712256841
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1712256841
transform 1 0 1736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1712256841
transform 1 0 1728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1712256841
transform 1 0 1720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1712256841
transform 1 0 1680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1712256841
transform 1 0 1648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1712256841
transform 1 0 1640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1712256841
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1712256841
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1712256841
transform 1 0 1584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1712256841
transform 1 0 1576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1712256841
transform 1 0 1544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1712256841
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1712256841
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1712256841
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1712256841
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1712256841
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1712256841
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1712256841
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1712256841
transform 1 0 1416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1712256841
transform 1 0 1376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1712256841
transform 1 0 1344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1712256841
transform 1 0 1336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1712256841
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1712256841
transform 1 0 1320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1712256841
transform 1 0 1256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1712256841
transform 1 0 1248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1712256841
transform 1 0 1240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1712256841
transform 1 0 1232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1712256841
transform 1 0 1224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1712256841
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1712256841
transform 1 0 1144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1712256841
transform 1 0 1136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1712256841
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1712256841
transform 1 0 1056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1712256841
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1712256841
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1712256841
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1712256841
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1712256841
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1712256841
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1712256841
transform 1 0 944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1712256841
transform 1 0 912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1712256841
transform 1 0 904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1712256841
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1712256841
transform 1 0 840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1712256841
transform 1 0 832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1712256841
transform 1 0 824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1712256841
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1712256841
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1712256841
transform 1 0 768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1712256841
transform 1 0 728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1712256841
transform 1 0 720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1712256841
transform 1 0 712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1712256841
transform 1 0 704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1712256841
transform 1 0 664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1712256841
transform 1 0 656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1712256841
transform 1 0 616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1712256841
transform 1 0 608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1712256841
transform 1 0 600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1712256841
transform 1 0 592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1712256841
transform 1 0 544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1712256841
transform 1 0 536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1712256841
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1712256841
transform 1 0 488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1712256841
transform 1 0 480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1712256841
transform 1 0 440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1712256841
transform 1 0 432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1712256841
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1712256841
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1712256841
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1712256841
transform 1 0 360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1712256841
transform 1 0 312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1712256841
transform 1 0 304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1712256841
transform 1 0 296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1712256841
transform 1 0 288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1712256841
transform 1 0 280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1712256841
transform 1 0 240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1712256841
transform 1 0 200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1712256841
transform 1 0 192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1712256841
transform 1 0 184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1712256841
transform 1 0 176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1712256841
transform 1 0 168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1712256841
transform 1 0 128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1712256841
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1712256841
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1712256841
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1712256841
transform 1 0 3424 0 1 1370
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1712256841
transform 1 0 3416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1712256841
transform 1 0 3408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1712256841
transform 1 0 3400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1712256841
transform 1 0 3336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1712256841
transform 1 0 3328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1712256841
transform 1 0 3320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1712256841
transform 1 0 3312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1712256841
transform 1 0 3304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1712256841
transform 1 0 3296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1712256841
transform 1 0 3240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1712256841
transform 1 0 3232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1712256841
transform 1 0 3224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1712256841
transform 1 0 3216 0 1 1370
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1712256841
transform 1 0 3208 0 1 1370
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1712256841
transform 1 0 3200 0 1 1370
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1712256841
transform 1 0 3168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1712256841
transform 1 0 3160 0 1 1370
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1712256841
transform 1 0 3152 0 1 1370
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1712256841
transform 1 0 3144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1712256841
transform 1 0 3136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1712256841
transform 1 0 3104 0 1 1370
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1712256841
transform 1 0 3064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1712256841
transform 1 0 3056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1712256841
transform 1 0 3048 0 1 1370
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1712256841
transform 1 0 3040 0 1 1370
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1712256841
transform 1 0 3032 0 1 1370
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1712256841
transform 1 0 3024 0 1 1370
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1712256841
transform 1 0 3016 0 1 1370
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1712256841
transform 1 0 2952 0 1 1370
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1712256841
transform 1 0 2944 0 1 1370
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1712256841
transform 1 0 2936 0 1 1370
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1712256841
transform 1 0 2928 0 1 1370
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1712256841
transform 1 0 2920 0 1 1370
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1712256841
transform 1 0 2912 0 1 1370
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1712256841
transform 1 0 2872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1712256841
transform 1 0 2832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1712256841
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1712256841
transform 1 0 2816 0 1 1370
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1712256841
transform 1 0 2808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1712256841
transform 1 0 2800 0 1 1370
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1712256841
transform 1 0 2792 0 1 1370
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1712256841
transform 1 0 2744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1712256841
transform 1 0 2736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1712256841
transform 1 0 2712 0 1 1370
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1712256841
transform 1 0 2704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1712256841
transform 1 0 2696 0 1 1370
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1712256841
transform 1 0 2688 0 1 1370
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1712256841
transform 1 0 2640 0 1 1370
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1712256841
transform 1 0 2632 0 1 1370
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1712256841
transform 1 0 2624 0 1 1370
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1712256841
transform 1 0 2616 0 1 1370
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1712256841
transform 1 0 2576 0 1 1370
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1712256841
transform 1 0 2568 0 1 1370
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1712256841
transform 1 0 2528 0 1 1370
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1712256841
transform 1 0 2520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1712256841
transform 1 0 2512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1712256841
transform 1 0 2504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1712256841
transform 1 0 2496 0 1 1370
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1712256841
transform 1 0 2488 0 1 1370
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1712256841
transform 1 0 2440 0 1 1370
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1712256841
transform 1 0 2432 0 1 1370
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1712256841
transform 1 0 2424 0 1 1370
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1712256841
transform 1 0 2384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1712256841
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1712256841
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1712256841
transform 1 0 2344 0 1 1370
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1712256841
transform 1 0 2336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1712256841
transform 1 0 2328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1712256841
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1712256841
transform 1 0 2264 0 1 1370
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1712256841
transform 1 0 2256 0 1 1370
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1712256841
transform 1 0 2248 0 1 1370
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1712256841
transform 1 0 2240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1712256841
transform 1 0 2232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1712256841
transform 1 0 2192 0 1 1370
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1712256841
transform 1 0 2152 0 1 1370
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1712256841
transform 1 0 2144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1712256841
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1712256841
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1712256841
transform 1 0 2088 0 1 1370
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1712256841
transform 1 0 2080 0 1 1370
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1712256841
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1712256841
transform 1 0 2032 0 1 1370
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1712256841
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1712256841
transform 1 0 2000 0 1 1370
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1712256841
transform 1 0 1992 0 1 1370
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1712256841
transform 1 0 1984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1712256841
transform 1 0 1944 0 1 1370
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1712256841
transform 1 0 1936 0 1 1370
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1712256841
transform 1 0 1896 0 1 1370
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1712256841
transform 1 0 1888 0 1 1370
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1712256841
transform 1 0 1880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1712256841
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1712256841
transform 1 0 1864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1712256841
transform 1 0 1808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1712256841
transform 1 0 1800 0 1 1370
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1712256841
transform 1 0 1792 0 1 1370
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1712256841
transform 1 0 1784 0 1 1370
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1712256841
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1712256841
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1712256841
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1712256841
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1712256841
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1712256841
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1712256841
transform 1 0 1672 0 1 1370
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1712256841
transform 1 0 1616 0 1 1370
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1712256841
transform 1 0 1608 0 1 1370
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1712256841
transform 1 0 1600 0 1 1370
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1712256841
transform 1 0 1592 0 1 1370
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1712256841
transform 1 0 1584 0 1 1370
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1712256841
transform 1 0 1576 0 1 1370
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1712256841
transform 1 0 1520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1712256841
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1712256841
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1712256841
transform 1 0 1496 0 1 1370
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1712256841
transform 1 0 1488 0 1 1370
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1712256841
transform 1 0 1480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1712256841
transform 1 0 1416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1712256841
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1712256841
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1712256841
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1712256841
transform 1 0 1384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1712256841
transform 1 0 1376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1712256841
transform 1 0 1344 0 1 1370
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1712256841
transform 1 0 1336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1712256841
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1712256841
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1712256841
transform 1 0 1272 0 1 1370
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1712256841
transform 1 0 1264 0 1 1370
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1712256841
transform 1 0 1232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1712256841
transform 1 0 1224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1712256841
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1712256841
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1712256841
transform 1 0 1168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1712256841
transform 1 0 1160 0 1 1370
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1712256841
transform 1 0 1120 0 1 1370
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1712256841
transform 1 0 1112 0 1 1370
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1712256841
transform 1 0 1104 0 1 1370
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1712256841
transform 1 0 1056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1712256841
transform 1 0 1048 0 1 1370
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1712256841
transform 1 0 1024 0 1 1370
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1712256841
transform 1 0 1016 0 1 1370
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1712256841
transform 1 0 1008 0 1 1370
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1712256841
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1712256841
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1712256841
transform 1 0 944 0 1 1370
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1712256841
transform 1 0 904 0 1 1370
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1712256841
transform 1 0 896 0 1 1370
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1712256841
transform 1 0 888 0 1 1370
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1712256841
transform 1 0 880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1712256841
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1712256841
transform 1 0 808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1712256841
transform 1 0 800 0 1 1370
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1712256841
transform 1 0 792 0 1 1370
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1712256841
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1712256841
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1712256841
transform 1 0 704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1712256841
transform 1 0 696 0 1 1370
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1712256841
transform 1 0 688 0 1 1370
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1712256841
transform 1 0 680 0 1 1370
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1712256841
transform 1 0 672 0 1 1370
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1712256841
transform 1 0 616 0 1 1370
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1712256841
transform 1 0 608 0 1 1370
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1712256841
transform 1 0 600 0 1 1370
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1712256841
transform 1 0 592 0 1 1370
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1712256841
transform 1 0 544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1712256841
transform 1 0 536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1712256841
transform 1 0 488 0 1 1370
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1712256841
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1712256841
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1712256841
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1712256841
transform 1 0 456 0 1 1370
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1712256841
transform 1 0 384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1712256841
transform 1 0 376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1712256841
transform 1 0 368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1712256841
transform 1 0 360 0 1 1370
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1712256841
transform 1 0 352 0 1 1370
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1712256841
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1712256841
transform 1 0 264 0 1 1370
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1712256841
transform 1 0 256 0 1 1370
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1712256841
transform 1 0 248 0 1 1370
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1712256841
transform 1 0 240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1712256841
transform 1 0 232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1712256841
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1712256841
transform 1 0 144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1712256841
transform 1 0 136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1712256841
transform 1 0 128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1712256841
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1712256841
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1712256841
transform 1 0 3424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1712256841
transform 1 0 3416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1712256841
transform 1 0 3408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1712256841
transform 1 0 3384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1712256841
transform 1 0 3328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1712256841
transform 1 0 3320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1712256841
transform 1 0 3312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1712256841
transform 1 0 3304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1712256841
transform 1 0 3296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1712256841
transform 1 0 3232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1712256841
transform 1 0 3224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1712256841
transform 1 0 3216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1712256841
transform 1 0 3112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1712256841
transform 1 0 3104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1712256841
transform 1 0 3096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1712256841
transform 1 0 3088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1712256841
transform 1 0 3080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1712256841
transform 1 0 3024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1712256841
transform 1 0 3016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1712256841
transform 1 0 3008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1712256841
transform 1 0 3000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1712256841
transform 1 0 2960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1712256841
transform 1 0 2952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1712256841
transform 1 0 2904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1712256841
transform 1 0 2896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1712256841
transform 1 0 2888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1712256841
transform 1 0 2880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1712256841
transform 1 0 2872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1712256841
transform 1 0 2824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1712256841
transform 1 0 2816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1712256841
transform 1 0 2808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1712256841
transform 1 0 2800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1712256841
transform 1 0 2744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1712256841
transform 1 0 2736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1712256841
transform 1 0 2728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1712256841
transform 1 0 2720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1712256841
transform 1 0 2712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1712256841
transform 1 0 2704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1712256841
transform 1 0 2696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1712256841
transform 1 0 2632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1712256841
transform 1 0 2624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1712256841
transform 1 0 2616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1712256841
transform 1 0 2576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1712256841
transform 1 0 2568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1712256841
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1712256841
transform 1 0 2552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1712256841
transform 1 0 2544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1712256841
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1712256841
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1712256841
transform 1 0 2480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1712256841
transform 1 0 2448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1712256841
transform 1 0 2440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1712256841
transform 1 0 2432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1712256841
transform 1 0 2424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1712256841
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1712256841
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1712256841
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1712256841
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1712256841
transform 1 0 2312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1712256841
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1712256841
transform 1 0 2296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1712256841
transform 1 0 2288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1712256841
transform 1 0 2248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1712256841
transform 1 0 2240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1712256841
transform 1 0 2232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1712256841
transform 1 0 2224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1712256841
transform 1 0 2184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1712256841
transform 1 0 2176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1712256841
transform 1 0 2168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1712256841
transform 1 0 2160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1712256841
transform 1 0 2112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1712256841
transform 1 0 2104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1712256841
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1712256841
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1712256841
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1712256841
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1712256841
transform 1 0 2048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1712256841
transform 1 0 2016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1712256841
transform 1 0 2008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1712256841
transform 1 0 2000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1712256841
transform 1 0 1992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1712256841
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1712256841
transform 1 0 1952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1712256841
transform 1 0 1944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1712256841
transform 1 0 1912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1712256841
transform 1 0 1904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1712256841
transform 1 0 1896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1712256841
transform 1 0 1888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1712256841
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1712256841
transform 1 0 1832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1712256841
transform 1 0 1824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1712256841
transform 1 0 1816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1712256841
transform 1 0 1808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1712256841
transform 1 0 1800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1712256841
transform 1 0 1760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1712256841
transform 1 0 1752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1712256841
transform 1 0 1744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1712256841
transform 1 0 1736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1712256841
transform 1 0 1696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1712256841
transform 1 0 1688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1712256841
transform 1 0 1680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1712256841
transform 1 0 1672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1712256841
transform 1 0 1664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1712256841
transform 1 0 1656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1712256841
transform 1 0 1616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1712256841
transform 1 0 1608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1712256841
transform 1 0 1600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1712256841
transform 1 0 1592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1712256841
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1712256841
transform 1 0 1536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1712256841
transform 1 0 1528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1712256841
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1712256841
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1712256841
transform 1 0 1504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1712256841
transform 1 0 1496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1712256841
transform 1 0 1488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1712256841
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1712256841
transform 1 0 1432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1712256841
transform 1 0 1424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1712256841
transform 1 0 1416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1712256841
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1712256841
transform 1 0 1376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1712256841
transform 1 0 1368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1712256841
transform 1 0 1360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1712256841
transform 1 0 1336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1712256841
transform 1 0 1312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1712256841
transform 1 0 1304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1712256841
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1712256841
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1712256841
transform 1 0 1280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1712256841
transform 1 0 1272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1712256841
transform 1 0 1224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1712256841
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1712256841
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1712256841
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1712256841
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1712256841
transform 1 0 1144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1712256841
transform 1 0 1136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1712256841
transform 1 0 1128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1712256841
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1712256841
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1712256841
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1712256841
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1712256841
transform 1 0 1048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1712256841
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1712256841
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1712256841
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1712256841
transform 1 0 1016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1712256841
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1712256841
transform 1 0 960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1712256841
transform 1 0 952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1712256841
transform 1 0 944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1712256841
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1712256841
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1712256841
transform 1 0 904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1712256841
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1712256841
transform 1 0 864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1712256841
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1712256841
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1712256841
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1712256841
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1712256841
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1712256841
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1712256841
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1712256841
transform 1 0 752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1712256841
transform 1 0 712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1712256841
transform 1 0 704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1712256841
transform 1 0 696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1712256841
transform 1 0 688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1712256841
transform 1 0 680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1712256841
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1712256841
transform 1 0 632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1712256841
transform 1 0 624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1712256841
transform 1 0 616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1712256841
transform 1 0 608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1712256841
transform 1 0 560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1712256841
transform 1 0 552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1712256841
transform 1 0 544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1712256841
transform 1 0 536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1712256841
transform 1 0 528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1712256841
transform 1 0 520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1712256841
transform 1 0 472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1712256841
transform 1 0 464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1712256841
transform 1 0 456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1712256841
transform 1 0 448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1712256841
transform 1 0 440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1712256841
transform 1 0 432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1712256841
transform 1 0 424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1712256841
transform 1 0 368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1712256841
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1712256841
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1712256841
transform 1 0 344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1712256841
transform 1 0 336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1712256841
transform 1 0 312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1712256841
transform 1 0 304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1712256841
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1712256841
transform 1 0 256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1712256841
transform 1 0 248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1712256841
transform 1 0 240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1712256841
transform 1 0 216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1712256841
transform 1 0 208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1712256841
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1712256841
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1712256841
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1712256841
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1712256841
transform 1 0 128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1712256841
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1712256841
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1712256841
transform 1 0 104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1712256841
transform 1 0 96 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1712256841
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1712256841
transform 1 0 3424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1712256841
transform 1 0 3416 0 1 1170
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1712256841
transform 1 0 3376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1712256841
transform 1 0 3368 0 1 1170
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1712256841
transform 1 0 3360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1712256841
transform 1 0 3352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1712256841
transform 1 0 3304 0 1 1170
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1712256841
transform 1 0 3296 0 1 1170
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1712256841
transform 1 0 3288 0 1 1170
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1712256841
transform 1 0 3280 0 1 1170
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1712256841
transform 1 0 3240 0 1 1170
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1712256841
transform 1 0 3232 0 1 1170
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1712256841
transform 1 0 3224 0 1 1170
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1712256841
transform 1 0 3216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1712256841
transform 1 0 3176 0 1 1170
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1712256841
transform 1 0 3168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1712256841
transform 1 0 3160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1712256841
transform 1 0 3120 0 1 1170
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1712256841
transform 1 0 3112 0 1 1170
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1712256841
transform 1 0 3104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1712256841
transform 1 0 3096 0 1 1170
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1712256841
transform 1 0 3088 0 1 1170
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1712256841
transform 1 0 3048 0 1 1170
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1712256841
transform 1 0 3040 0 1 1170
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1712256841
transform 1 0 3000 0 1 1170
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1712256841
transform 1 0 2992 0 1 1170
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1712256841
transform 1 0 2984 0 1 1170
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1712256841
transform 1 0 2976 0 1 1170
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1712256841
transform 1 0 2944 0 1 1170
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1712256841
transform 1 0 2936 0 1 1170
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1712256841
transform 1 0 2888 0 1 1170
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1712256841
transform 1 0 2880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1712256841
transform 1 0 2872 0 1 1170
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1712256841
transform 1 0 2864 0 1 1170
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1712256841
transform 1 0 2856 0 1 1170
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1712256841
transform 1 0 2848 0 1 1170
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1712256841
transform 1 0 2792 0 1 1170
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1712256841
transform 1 0 2784 0 1 1170
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1712256841
transform 1 0 2776 0 1 1170
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1712256841
transform 1 0 2744 0 1 1170
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1712256841
transform 1 0 2736 0 1 1170
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1712256841
transform 1 0 2728 0 1 1170
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1712256841
transform 1 0 2720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1712256841
transform 1 0 2696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1712256841
transform 1 0 2664 0 1 1170
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1712256841
transform 1 0 2640 0 1 1170
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1712256841
transform 1 0 2632 0 1 1170
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1712256841
transform 1 0 2624 0 1 1170
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1712256841
transform 1 0 2616 0 1 1170
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1712256841
transform 1 0 2608 0 1 1170
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1712256841
transform 1 0 2600 0 1 1170
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1712256841
transform 1 0 2552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1712256841
transform 1 0 2544 0 1 1170
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1712256841
transform 1 0 2536 0 1 1170
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1712256841
transform 1 0 2528 0 1 1170
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1712256841
transform 1 0 2496 0 1 1170
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1712256841
transform 1 0 2464 0 1 1170
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1712256841
transform 1 0 2456 0 1 1170
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1712256841
transform 1 0 2448 0 1 1170
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1712256841
transform 1 0 2440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1712256841
transform 1 0 2432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1712256841
transform 1 0 2400 0 1 1170
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1712256841
transform 1 0 2376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1712256841
transform 1 0 2368 0 1 1170
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1712256841
transform 1 0 2360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1712256841
transform 1 0 2320 0 1 1170
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1712256841
transform 1 0 2312 0 1 1170
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1712256841
transform 1 0 2304 0 1 1170
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1712256841
transform 1 0 2296 0 1 1170
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1712256841
transform 1 0 2288 0 1 1170
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1712256841
transform 1 0 2240 0 1 1170
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1712256841
transform 1 0 2232 0 1 1170
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1712256841
transform 1 0 2224 0 1 1170
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1712256841
transform 1 0 2192 0 1 1170
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1712256841
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1712256841
transform 1 0 2176 0 1 1170
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1712256841
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1712256841
transform 1 0 2120 0 1 1170
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1712256841
transform 1 0 2112 0 1 1170
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1712256841
transform 1 0 2104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1712256841
transform 1 0 2096 0 1 1170
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1712256841
transform 1 0 2088 0 1 1170
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1712256841
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_3130
timestamp 1712256841
transform 1 0 2040 0 1 1170
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1712256841
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1712256841
transform 1 0 2000 0 1 1170
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1712256841
transform 1 0 1992 0 1 1170
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1712256841
transform 1 0 1984 0 1 1170
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1712256841
transform 1 0 1944 0 1 1170
box -8 -3 16 105
use FILL  FILL_3136
timestamp 1712256841
transform 1 0 1936 0 1 1170
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1712256841
transform 1 0 1928 0 1 1170
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1712256841
transform 1 0 1920 0 1 1170
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1712256841
transform 1 0 1880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1712256841
transform 1 0 1872 0 1 1170
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1712256841
transform 1 0 1864 0 1 1170
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1712256841
transform 1 0 1824 0 1 1170
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1712256841
transform 1 0 1816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1712256841
transform 1 0 1808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1712256841
transform 1 0 1800 0 1 1170
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1712256841
transform 1 0 1760 0 1 1170
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1712256841
transform 1 0 1752 0 1 1170
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1712256841
transform 1 0 1744 0 1 1170
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1712256841
transform 1 0 1736 0 1 1170
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1712256841
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1712256841
transform 1 0 1672 0 1 1170
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1712256841
transform 1 0 1664 0 1 1170
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1712256841
transform 1 0 1656 0 1 1170
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1712256841
transform 1 0 1648 0 1 1170
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1712256841
transform 1 0 1640 0 1 1170
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1712256841
transform 1 0 1592 0 1 1170
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1712256841
transform 1 0 1584 0 1 1170
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1712256841
transform 1 0 1576 0 1 1170
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1712256841
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1712256841
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1712256841
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1712256841
transform 1 0 1512 0 1 1170
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1712256841
transform 1 0 1504 0 1 1170
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1712256841
transform 1 0 1456 0 1 1170
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1712256841
transform 1 0 1448 0 1 1170
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1712256841
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1712256841
transform 1 0 1432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1712256841
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1712256841
transform 1 0 1384 0 1 1170
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1712256841
transform 1 0 1376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1712256841
transform 1 0 1368 0 1 1170
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1712256841
transform 1 0 1328 0 1 1170
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1712256841
transform 1 0 1320 0 1 1170
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1712256841
transform 1 0 1312 0 1 1170
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1712256841
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1712256841
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1712256841
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1712256841
transform 1 0 1240 0 1 1170
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1712256841
transform 1 0 1232 0 1 1170
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1712256841
transform 1 0 1224 0 1 1170
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1712256841
transform 1 0 1216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1712256841
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1712256841
transform 1 0 1160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1712256841
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1712256841
transform 1 0 1144 0 1 1170
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1712256841
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1712256841
transform 1 0 1104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1712256841
transform 1 0 1096 0 1 1170
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1712256841
transform 1 0 1064 0 1 1170
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1712256841
transform 1 0 1056 0 1 1170
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1712256841
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1712256841
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1712256841
transform 1 0 1000 0 1 1170
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1712256841
transform 1 0 992 0 1 1170
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1712256841
transform 1 0 944 0 1 1170
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1712256841
transform 1 0 936 0 1 1170
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1712256841
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1712256841
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1712256841
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1712256841
transform 1 0 872 0 1 1170
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1712256841
transform 1 0 864 0 1 1170
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1712256841
transform 1 0 856 0 1 1170
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1712256841
transform 1 0 816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1712256841
transform 1 0 808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1712256841
transform 1 0 800 0 1 1170
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1712256841
transform 1 0 792 0 1 1170
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1712256841
transform 1 0 784 0 1 1170
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1712256841
transform 1 0 776 0 1 1170
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1712256841
transform 1 0 728 0 1 1170
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1712256841
transform 1 0 720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1712256841
transform 1 0 712 0 1 1170
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1712256841
transform 1 0 704 0 1 1170
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1712256841
transform 1 0 696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1712256841
transform 1 0 688 0 1 1170
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1712256841
transform 1 0 632 0 1 1170
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1712256841
transform 1 0 624 0 1 1170
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1712256841
transform 1 0 616 0 1 1170
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1712256841
transform 1 0 608 0 1 1170
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1712256841
transform 1 0 568 0 1 1170
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1712256841
transform 1 0 560 0 1 1170
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1712256841
transform 1 0 552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1712256841
transform 1 0 544 0 1 1170
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1712256841
transform 1 0 536 0 1 1170
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1712256841
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1712256841
transform 1 0 480 0 1 1170
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1712256841
transform 1 0 472 0 1 1170
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1712256841
transform 1 0 440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1712256841
transform 1 0 432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1712256841
transform 1 0 424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1712256841
transform 1 0 416 0 1 1170
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1712256841
transform 1 0 408 0 1 1170
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1712256841
transform 1 0 360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1712256841
transform 1 0 352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1712256841
transform 1 0 344 0 1 1170
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1712256841
transform 1 0 336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1712256841
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1712256841
transform 1 0 288 0 1 1170
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1712256841
transform 1 0 280 0 1 1170
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1712256841
transform 1 0 272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1712256841
transform 1 0 264 0 1 1170
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1712256841
transform 1 0 256 0 1 1170
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1712256841
transform 1 0 216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1712256841
transform 1 0 208 0 1 1170
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1712256841
transform 1 0 200 0 1 1170
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1712256841
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1712256841
transform 1 0 184 0 1 1170
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1712256841
transform 1 0 152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1712256841
transform 1 0 144 0 1 1170
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1712256841
transform 1 0 136 0 1 1170
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1712256841
transform 1 0 128 0 1 1170
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1712256841
transform 1 0 88 0 1 1170
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1712256841
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1712256841
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1712256841
transform 1 0 3424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1712256841
transform 1 0 3416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1712256841
transform 1 0 3376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1712256841
transform 1 0 3368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1712256841
transform 1 0 3360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1712256841
transform 1 0 3336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1712256841
transform 1 0 3328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1712256841
transform 1 0 3320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1712256841
transform 1 0 3312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1712256841
transform 1 0 3264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1712256841
transform 1 0 3256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1712256841
transform 1 0 3248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1712256841
transform 1 0 3240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1712256841
transform 1 0 3232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1712256841
transform 1 0 3224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1712256841
transform 1 0 3216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1712256841
transform 1 0 3168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1712256841
transform 1 0 3160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1712256841
transform 1 0 3120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1712256841
transform 1 0 3112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1712256841
transform 1 0 3104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1712256841
transform 1 0 3096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1712256841
transform 1 0 3088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1712256841
transform 1 0 3080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1712256841
transform 1 0 3072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1712256841
transform 1 0 3064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1712256841
transform 1 0 3056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1712256841
transform 1 0 3048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1712256841
transform 1 0 3040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1712256841
transform 1 0 3032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1712256841
transform 1 0 3024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1712256841
transform 1 0 3016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1712256841
transform 1 0 3008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1712256841
transform 1 0 3000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1712256841
transform 1 0 2976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1712256841
transform 1 0 2968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1712256841
transform 1 0 2960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1712256841
transform 1 0 2952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1712256841
transform 1 0 2944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1712256841
transform 1 0 2912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1712256841
transform 1 0 2904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1712256841
transform 1 0 2896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1712256841
transform 1 0 2856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1712256841
transform 1 0 2848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1712256841
transform 1 0 2840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1712256841
transform 1 0 2816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1712256841
transform 1 0 2808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1712256841
transform 1 0 2800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1712256841
transform 1 0 2792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1712256841
transform 1 0 2760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1712256841
transform 1 0 2752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1712256841
transform 1 0 2744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1712256841
transform 1 0 2736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1712256841
transform 1 0 2704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1712256841
transform 1 0 2696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1712256841
transform 1 0 2656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1712256841
transform 1 0 2648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1712256841
transform 1 0 2640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1712256841
transform 1 0 2632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1712256841
transform 1 0 2584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1712256841
transform 1 0 2576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1712256841
transform 1 0 2568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1712256841
transform 1 0 2560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1712256841
transform 1 0 2552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1712256841
transform 1 0 2544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1712256841
transform 1 0 2512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1712256841
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1712256841
transform 1 0 2472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1712256841
transform 1 0 2464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1712256841
transform 1 0 2456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1712256841
transform 1 0 2448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1712256841
transform 1 0 2440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1712256841
transform 1 0 2392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1712256841
transform 1 0 2384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1712256841
transform 1 0 2376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3329
timestamp 1712256841
transform 1 0 2368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1712256841
transform 1 0 2360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1712256841
transform 1 0 2320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1712256841
transform 1 0 2312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1712256841
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1712256841
transform 1 0 2296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1712256841
transform 1 0 2264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1712256841
transform 1 0 2256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1712256841
transform 1 0 2248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1712256841
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1712256841
transform 1 0 2208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1712256841
transform 1 0 2200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1712256841
transform 1 0 2176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1712256841
transform 1 0 2168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1712256841
transform 1 0 2160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1712256841
transform 1 0 2152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1712256841
transform 1 0 2112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1712256841
transform 1 0 2104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1712256841
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1712256841
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1712256841
transform 1 0 2056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1712256841
transform 1 0 2048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1712256841
transform 1 0 2040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1712256841
transform 1 0 2032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1712256841
transform 1 0 2008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1712256841
transform 1 0 2000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1712256841
transform 1 0 1960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1712256841
transform 1 0 1952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1712256841
transform 1 0 1944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1712256841
transform 1 0 1936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1712256841
transform 1 0 1928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1712256841
transform 1 0 1920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1712256841
transform 1 0 1888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1712256841
transform 1 0 1856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1712256841
transform 1 0 1848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1712256841
transform 1 0 1840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1712256841
transform 1 0 1832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1712256841
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1712256841
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1712256841
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1712256841
transform 1 0 1760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1712256841
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1712256841
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1712256841
transform 1 0 1736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1712256841
transform 1 0 1712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1712256841
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1712256841
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1712256841
transform 1 0 1688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1712256841
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1712256841
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1712256841
transform 1 0 1632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3380
timestamp 1712256841
transform 1 0 1624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1712256841
transform 1 0 1600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1712256841
transform 1 0 1592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1712256841
transform 1 0 1568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1712256841
transform 1 0 1560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1712256841
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1712256841
transform 1 0 1544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1712256841
transform 1 0 1504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1712256841
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1712256841
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1712256841
transform 1 0 1480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1712256841
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1712256841
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1712256841
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1712256841
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1712256841
transform 1 0 1392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1712256841
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1712256841
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1712256841
transform 1 0 1336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3399
timestamp 1712256841
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1712256841
transform 1 0 1320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1712256841
transform 1 0 1288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1712256841
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1712256841
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1712256841
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1712256841
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1712256841
transform 1 0 1224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1712256841
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1712256841
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1712256841
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1712256841
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1712256841
transform 1 0 1160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1712256841
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1712256841
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1712256841
transform 1 0 1112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1712256841
transform 1 0 1104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1712256841
transform 1 0 1056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1712256841
transform 1 0 1048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1712256841
transform 1 0 1040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1712256841
transform 1 0 1032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1712256841
transform 1 0 1024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1712256841
transform 1 0 1016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1712256841
transform 1 0 984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1712256841
transform 1 0 976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1712256841
transform 1 0 944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1712256841
transform 1 0 936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1712256841
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1712256841
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1712256841
transform 1 0 888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1712256841
transform 1 0 880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1712256841
transform 1 0 872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1712256841
transform 1 0 832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1712256841
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1712256841
transform 1 0 816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1712256841
transform 1 0 808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1712256841
transform 1 0 784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1712256841
transform 1 0 744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1712256841
transform 1 0 736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1712256841
transform 1 0 728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1712256841
transform 1 0 720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1712256841
transform 1 0 712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1712256841
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1712256841
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1712256841
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1712256841
transform 1 0 632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1712256841
transform 1 0 624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1712256841
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1712256841
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3448
timestamp 1712256841
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1712256841
transform 1 0 528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1712256841
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1712256841
transform 1 0 512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1712256841
transform 1 0 504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1712256841
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1712256841
transform 1 0 448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1712256841
transform 1 0 440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1712256841
transform 1 0 432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1712256841
transform 1 0 384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3458
timestamp 1712256841
transform 1 0 376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1712256841
transform 1 0 368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1712256841
transform 1 0 360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1712256841
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1712256841
transform 1 0 288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1712256841
transform 1 0 280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3464
timestamp 1712256841
transform 1 0 272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1712256841
transform 1 0 264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1712256841
transform 1 0 256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1712256841
transform 1 0 248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1712256841
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3469
timestamp 1712256841
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1712256841
transform 1 0 168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1712256841
transform 1 0 160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1712256841
transform 1 0 152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1712256841
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1712256841
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1712256841
transform 1 0 3424 0 1 970
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1712256841
transform 1 0 3384 0 1 970
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1712256841
transform 1 0 3376 0 1 970
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1712256841
transform 1 0 3344 0 1 970
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1712256841
transform 1 0 3336 0 1 970
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1712256841
transform 1 0 3328 0 1 970
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1712256841
transform 1 0 3280 0 1 970
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1712256841
transform 1 0 3272 0 1 970
box -8 -3 16 105
use FILL  FILL_3483
timestamp 1712256841
transform 1 0 3224 0 1 970
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1712256841
transform 1 0 3216 0 1 970
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1712256841
transform 1 0 3208 0 1 970
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1712256841
transform 1 0 3200 0 1 970
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1712256841
transform 1 0 3192 0 1 970
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1712256841
transform 1 0 3128 0 1 970
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1712256841
transform 1 0 3120 0 1 970
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1712256841
transform 1 0 3016 0 1 970
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1712256841
transform 1 0 3008 0 1 970
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1712256841
transform 1 0 3000 0 1 970
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1712256841
transform 1 0 2944 0 1 970
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1712256841
transform 1 0 2936 0 1 970
box -8 -3 16 105
use FILL  FILL_3495
timestamp 1712256841
transform 1 0 2928 0 1 970
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1712256841
transform 1 0 2920 0 1 970
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1712256841
transform 1 0 2912 0 1 970
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1712256841
transform 1 0 2872 0 1 970
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1712256841
transform 1 0 2864 0 1 970
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1712256841
transform 1 0 2856 0 1 970
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1712256841
transform 1 0 2816 0 1 970
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1712256841
transform 1 0 2808 0 1 970
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1712256841
transform 1 0 2800 0 1 970
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1712256841
transform 1 0 2792 0 1 970
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1712256841
transform 1 0 2752 0 1 970
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1712256841
transform 1 0 2744 0 1 970
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1712256841
transform 1 0 2736 0 1 970
box -8 -3 16 105
use FILL  FILL_3508
timestamp 1712256841
transform 1 0 2688 0 1 970
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1712256841
transform 1 0 2680 0 1 970
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1712256841
transform 1 0 2672 0 1 970
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1712256841
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1712256841
transform 1 0 2656 0 1 970
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1712256841
transform 1 0 2648 0 1 970
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1712256841
transform 1 0 2592 0 1 970
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1712256841
transform 1 0 2584 0 1 970
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1712256841
transform 1 0 2576 0 1 970
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1712256841
transform 1 0 2568 0 1 970
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1712256841
transform 1 0 2544 0 1 970
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1712256841
transform 1 0 2536 0 1 970
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1712256841
transform 1 0 2504 0 1 970
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1712256841
transform 1 0 2496 0 1 970
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1712256841
transform 1 0 2488 0 1 970
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1712256841
transform 1 0 2480 0 1 970
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1712256841
transform 1 0 2432 0 1 970
box -8 -3 16 105
use FILL  FILL_3525
timestamp 1712256841
transform 1 0 2424 0 1 970
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1712256841
transform 1 0 2416 0 1 970
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1712256841
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1712256841
transform 1 0 2360 0 1 970
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1712256841
transform 1 0 2352 0 1 970
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1712256841
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1712256841
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1712256841
transform 1 0 2296 0 1 970
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1712256841
transform 1 0 2288 0 1 970
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1712256841
transform 1 0 2280 0 1 970
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1712256841
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1712256841
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1712256841
transform 1 0 2224 0 1 970
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1712256841
transform 1 0 2216 0 1 970
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1712256841
transform 1 0 2176 0 1 970
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1712256841
transform 1 0 2168 0 1 970
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1712256841
transform 1 0 2160 0 1 970
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1712256841
transform 1 0 2128 0 1 970
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1712256841
transform 1 0 2120 0 1 970
box -8 -3 16 105
use FILL  FILL_3544
timestamp 1712256841
transform 1 0 2112 0 1 970
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1712256841
transform 1 0 2104 0 1 970
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1712256841
transform 1 0 2064 0 1 970
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1712256841
transform 1 0 2056 0 1 970
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1712256841
transform 1 0 2048 0 1 970
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1712256841
transform 1 0 2008 0 1 970
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1712256841
transform 1 0 2000 0 1 970
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1712256841
transform 1 0 1992 0 1 970
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1712256841
transform 1 0 1984 0 1 970
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1712256841
transform 1 0 1976 0 1 970
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1712256841
transform 1 0 1952 0 1 970
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1712256841
transform 1 0 1912 0 1 970
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1712256841
transform 1 0 1904 0 1 970
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1712256841
transform 1 0 1896 0 1 970
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1712256841
transform 1 0 1888 0 1 970
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1712256841
transform 1 0 1880 0 1 970
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1712256841
transform 1 0 1856 0 1 970
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1712256841
transform 1 0 1824 0 1 970
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1712256841
transform 1 0 1816 0 1 970
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1712256841
transform 1 0 1808 0 1 970
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1712256841
transform 1 0 1800 0 1 970
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1712256841
transform 1 0 1760 0 1 970
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1712256841
transform 1 0 1752 0 1 970
box -8 -3 16 105
use FILL  FILL_3567
timestamp 1712256841
transform 1 0 1744 0 1 970
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1712256841
transform 1 0 1712 0 1 970
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1712256841
transform 1 0 1704 0 1 970
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1712256841
transform 1 0 1696 0 1 970
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1712256841
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1712256841
transform 1 0 1648 0 1 970
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1712256841
transform 1 0 1640 0 1 970
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1712256841
transform 1 0 1632 0 1 970
box -8 -3 16 105
use FILL  FILL_3575
timestamp 1712256841
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1712256841
transform 1 0 1576 0 1 970
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1712256841
transform 1 0 1568 0 1 970
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1712256841
transform 1 0 1560 0 1 970
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1712256841
transform 1 0 1552 0 1 970
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1712256841
transform 1 0 1544 0 1 970
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1712256841
transform 1 0 1536 0 1 970
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1712256841
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1712256841
transform 1 0 1480 0 1 970
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1712256841
transform 1 0 1472 0 1 970
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1712256841
transform 1 0 1432 0 1 970
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1712256841
transform 1 0 1424 0 1 970
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1712256841
transform 1 0 1416 0 1 970
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1712256841
transform 1 0 1384 0 1 970
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1712256841
transform 1 0 1376 0 1 970
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1712256841
transform 1 0 1368 0 1 970
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1712256841
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1712256841
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1712256841
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1712256841
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1712256841
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1712256841
transform 1 0 1256 0 1 970
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1712256841
transform 1 0 1248 0 1 970
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1712256841
transform 1 0 1240 0 1 970
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1712256841
transform 1 0 1232 0 1 970
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1712256841
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1712256841
transform 1 0 1192 0 1 970
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1712256841
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1712256841
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1712256841
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1712256841
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1712256841
transform 1 0 1120 0 1 970
box -8 -3 16 105
use FILL  FILL_3607
timestamp 1712256841
transform 1 0 1080 0 1 970
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1712256841
transform 1 0 1072 0 1 970
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1712256841
transform 1 0 1064 0 1 970
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1712256841
transform 1 0 1056 0 1 970
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1712256841
transform 1 0 1016 0 1 970
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1712256841
transform 1 0 1008 0 1 970
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1712256841
transform 1 0 1000 0 1 970
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1712256841
transform 1 0 960 0 1 970
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1712256841
transform 1 0 952 0 1 970
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1712256841
transform 1 0 944 0 1 970
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1712256841
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1712256841
transform 1 0 928 0 1 970
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1712256841
transform 1 0 904 0 1 970
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1712256841
transform 1 0 872 0 1 970
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1712256841
transform 1 0 864 0 1 970
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1712256841
transform 1 0 856 0 1 970
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1712256841
transform 1 0 848 0 1 970
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1712256841
transform 1 0 808 0 1 970
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1712256841
transform 1 0 800 0 1 970
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1712256841
transform 1 0 792 0 1 970
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1712256841
transform 1 0 784 0 1 970
box -8 -3 16 105
use FILL  FILL_3628
timestamp 1712256841
transform 1 0 776 0 1 970
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1712256841
transform 1 0 736 0 1 970
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1712256841
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1712256841
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1712256841
transform 1 0 712 0 1 970
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1712256841
transform 1 0 704 0 1 970
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1712256841
transform 1 0 664 0 1 970
box -8 -3 16 105
use FILL  FILL_3635
timestamp 1712256841
transform 1 0 656 0 1 970
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1712256841
transform 1 0 648 0 1 970
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1712256841
transform 1 0 624 0 1 970
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1712256841
transform 1 0 592 0 1 970
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1712256841
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1712256841
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1712256841
transform 1 0 568 0 1 970
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1712256841
transform 1 0 560 0 1 970
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1712256841
transform 1 0 552 0 1 970
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1712256841
transform 1 0 496 0 1 970
box -8 -3 16 105
use FILL  FILL_3645
timestamp 1712256841
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1712256841
transform 1 0 480 0 1 970
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1712256841
transform 1 0 472 0 1 970
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1712256841
transform 1 0 464 0 1 970
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1712256841
transform 1 0 416 0 1 970
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1712256841
transform 1 0 408 0 1 970
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1712256841
transform 1 0 400 0 1 970
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1712256841
transform 1 0 392 0 1 970
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1712256841
transform 1 0 384 0 1 970
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1712256841
transform 1 0 376 0 1 970
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1712256841
transform 1 0 344 0 1 970
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1712256841
transform 1 0 336 0 1 970
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1712256841
transform 1 0 328 0 1 970
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1712256841
transform 1 0 288 0 1 970
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1712256841
transform 1 0 280 0 1 970
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1712256841
transform 1 0 272 0 1 970
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1712256841
transform 1 0 264 0 1 970
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1712256841
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1712256841
transform 1 0 248 0 1 970
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1712256841
transform 1 0 240 0 1 970
box -8 -3 16 105
use FILL  FILL_3665
timestamp 1712256841
transform 1 0 192 0 1 970
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1712256841
transform 1 0 184 0 1 970
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1712256841
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1712256841
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1712256841
transform 1 0 160 0 1 970
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1712256841
transform 1 0 152 0 1 970
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1712256841
transform 1 0 120 0 1 970
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1712256841
transform 1 0 112 0 1 970
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1712256841
transform 1 0 88 0 1 970
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1712256841
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1712256841
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1712256841
transform 1 0 3424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3677
timestamp 1712256841
transform 1 0 3416 0 -1 970
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1712256841
transform 1 0 3360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1712256841
transform 1 0 3352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1712256841
transform 1 0 3312 0 -1 970
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1712256841
transform 1 0 3304 0 -1 970
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1712256841
transform 1 0 3296 0 -1 970
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1712256841
transform 1 0 3288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1712256841
transform 1 0 3232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1712256841
transform 1 0 3224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1712256841
transform 1 0 3216 0 -1 970
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1712256841
transform 1 0 3152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1712256841
transform 1 0 3144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1712256841
transform 1 0 3136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1712256841
transform 1 0 3032 0 -1 970
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1712256841
transform 1 0 3024 0 -1 970
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1712256841
transform 1 0 3016 0 -1 970
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1712256841
transform 1 0 2960 0 -1 970
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1712256841
transform 1 0 2952 0 -1 970
box -8 -3 16 105
use FILL  FILL_3695
timestamp 1712256841
transform 1 0 2944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1712256841
transform 1 0 2936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1712256841
transform 1 0 2896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1712256841
transform 1 0 2888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1712256841
transform 1 0 2880 0 -1 970
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1712256841
transform 1 0 2840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1712256841
transform 1 0 2832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1712256841
transform 1 0 2792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1712256841
transform 1 0 2784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1712256841
transform 1 0 2776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1712256841
transform 1 0 2736 0 -1 970
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1712256841
transform 1 0 2728 0 -1 970
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1712256841
transform 1 0 2720 0 -1 970
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1712256841
transform 1 0 2712 0 -1 970
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1712256841
transform 1 0 2688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1712256841
transform 1 0 2648 0 -1 970
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1712256841
transform 1 0 2640 0 -1 970
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1712256841
transform 1 0 2632 0 -1 970
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1712256841
transform 1 0 2584 0 -1 970
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1712256841
transform 1 0 2576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3715
timestamp 1712256841
transform 1 0 2568 0 -1 970
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1712256841
transform 1 0 2560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1712256841
transform 1 0 2512 0 -1 970
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1712256841
transform 1 0 2504 0 -1 970
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1712256841
transform 1 0 2496 0 -1 970
box -8 -3 16 105
use FILL  FILL_3720
timestamp 1712256841
transform 1 0 2448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1712256841
transform 1 0 2440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1712256841
transform 1 0 2432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1712256841
transform 1 0 2424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1712256841
transform 1 0 2376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1712256841
transform 1 0 2368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1712256841
transform 1 0 2360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1712256841
transform 1 0 2352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1712256841
transform 1 0 2320 0 -1 970
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1712256841
transform 1 0 2312 0 -1 970
box -8 -3 16 105
use FILL  FILL_3730
timestamp 1712256841
transform 1 0 2304 0 -1 970
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1712256841
transform 1 0 2272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1712256841
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1712256841
transform 1 0 2224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1712256841
transform 1 0 2216 0 -1 970
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1712256841
transform 1 0 2208 0 -1 970
box -8 -3 16 105
use FILL  FILL_3736
timestamp 1712256841
transform 1 0 2200 0 -1 970
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1712256841
transform 1 0 2152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1712256841
transform 1 0 2144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1712256841
transform 1 0 2136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1712256841
transform 1 0 2128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1712256841
transform 1 0 2120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1712256841
transform 1 0 2072 0 -1 970
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1712256841
transform 1 0 2064 0 -1 970
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1712256841
transform 1 0 2056 0 -1 970
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1712256841
transform 1 0 2024 0 -1 970
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1712256841
transform 1 0 2016 0 -1 970
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1712256841
transform 1 0 2008 0 -1 970
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1712256841
transform 1 0 1968 0 -1 970
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1712256841
transform 1 0 1960 0 -1 970
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1712256841
transform 1 0 1952 0 -1 970
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1712256841
transform 1 0 1944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1712256841
transform 1 0 1904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1712256841
transform 1 0 1896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1712256841
transform 1 0 1888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1712256841
transform 1 0 1880 0 -1 970
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1712256841
transform 1 0 1848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3757
timestamp 1712256841
transform 1 0 1840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1712256841
transform 1 0 1832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1712256841
transform 1 0 1792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1712256841
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1712256841
transform 1 0 1776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1712256841
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1712256841
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1712256841
transform 1 0 1728 0 -1 970
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1712256841
transform 1 0 1720 0 -1 970
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1712256841
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1712256841
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3768
timestamp 1712256841
transform 1 0 1672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1712256841
transform 1 0 1664 0 -1 970
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1712256841
transform 1 0 1640 0 -1 970
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1712256841
transform 1 0 1632 0 -1 970
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1712256841
transform 1 0 1600 0 -1 970
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1712256841
transform 1 0 1592 0 -1 970
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1712256841
transform 1 0 1584 0 -1 970
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1712256841
transform 1 0 1576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1712256841
transform 1 0 1536 0 -1 970
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1712256841
transform 1 0 1528 0 -1 970
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1712256841
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1712256841
transform 1 0 1512 0 -1 970
box -8 -3 16 105
use FILL  FILL_3780
timestamp 1712256841
transform 1 0 1504 0 -1 970
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1712256841
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1712256841
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1712256841
transform 1 0 1448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1712256841
transform 1 0 1440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3785
timestamp 1712256841
transform 1 0 1400 0 -1 970
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1712256841
transform 1 0 1392 0 -1 970
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1712256841
transform 1 0 1384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1712256841
transform 1 0 1376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3789
timestamp 1712256841
transform 1 0 1344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1712256841
transform 1 0 1336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1712256841
transform 1 0 1328 0 -1 970
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1712256841
transform 1 0 1320 0 -1 970
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1712256841
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1712256841
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1712256841
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1712256841
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1712256841
transform 1 0 1232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1712256841
transform 1 0 1224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1712256841
transform 1 0 1216 0 -1 970
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1712256841
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1712256841
transform 1 0 1168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1712256841
transform 1 0 1160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1712256841
transform 1 0 1120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1712256841
transform 1 0 1112 0 -1 970
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1712256841
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use FILL  FILL_3806
timestamp 1712256841
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1712256841
transform 1 0 1088 0 -1 970
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1712256841
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1712256841
transform 1 0 1032 0 -1 970
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1712256841
transform 1 0 1024 0 -1 970
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1712256841
transform 1 0 1016 0 -1 970
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1712256841
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1712256841
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1712256841
transform 1 0 976 0 -1 970
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1712256841
transform 1 0 968 0 -1 970
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1712256841
transform 1 0 928 0 -1 970
box -8 -3 16 105
use FILL  FILL_3817
timestamp 1712256841
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1712256841
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1712256841
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1712256841
transform 1 0 872 0 -1 970
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1712256841
transform 1 0 864 0 -1 970
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1712256841
transform 1 0 856 0 -1 970
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1712256841
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1712256841
transform 1 0 808 0 -1 970
box -8 -3 16 105
use FILL  FILL_3825
timestamp 1712256841
transform 1 0 800 0 -1 970
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1712256841
transform 1 0 792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1712256841
transform 1 0 752 0 -1 970
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1712256841
transform 1 0 744 0 -1 970
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1712256841
transform 1 0 736 0 -1 970
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1712256841
transform 1 0 728 0 -1 970
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1712256841
transform 1 0 688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1712256841
transform 1 0 680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1712256841
transform 1 0 672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1712256841
transform 1 0 664 0 -1 970
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1712256841
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1712256841
transform 1 0 616 0 -1 970
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1712256841
transform 1 0 608 0 -1 970
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1712256841
transform 1 0 600 0 -1 970
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1712256841
transform 1 0 560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1712256841
transform 1 0 552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3841
timestamp 1712256841
transform 1 0 544 0 -1 970
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1712256841
transform 1 0 536 0 -1 970
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1712256841
transform 1 0 488 0 -1 970
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1712256841
transform 1 0 480 0 -1 970
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1712256841
transform 1 0 440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1712256841
transform 1 0 432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1712256841
transform 1 0 424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1712256841
transform 1 0 392 0 -1 970
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1712256841
transform 1 0 384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1712256841
transform 1 0 376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1712256841
transform 1 0 336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1712256841
transform 1 0 328 0 -1 970
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1712256841
transform 1 0 320 0 -1 970
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1712256841
transform 1 0 312 0 -1 970
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1712256841
transform 1 0 304 0 -1 970
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1712256841
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3857
timestamp 1712256841
transform 1 0 264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1712256841
transform 1 0 240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1712256841
transform 1 0 232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1712256841
transform 1 0 224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1712256841
transform 1 0 200 0 -1 970
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1712256841
transform 1 0 192 0 -1 970
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1712256841
transform 1 0 184 0 -1 970
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1712256841
transform 1 0 152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1712256841
transform 1 0 144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1712256841
transform 1 0 136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1712256841
transform 1 0 128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1712256841
transform 1 0 120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1712256841
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1712256841
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1712256841
transform 1 0 3424 0 1 770
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1712256841
transform 1 0 3416 0 1 770
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1712256841
transform 1 0 3408 0 1 770
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1712256841
transform 1 0 3352 0 1 770
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1712256841
transform 1 0 3320 0 1 770
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1712256841
transform 1 0 3312 0 1 770
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1712256841
transform 1 0 3304 0 1 770
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1712256841
transform 1 0 3256 0 1 770
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1712256841
transform 1 0 3248 0 1 770
box -8 -3 16 105
use FILL  FILL_3880
timestamp 1712256841
transform 1 0 3240 0 1 770
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1712256841
transform 1 0 3232 0 1 770
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1712256841
transform 1 0 3224 0 1 770
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1712256841
transform 1 0 3192 0 1 770
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1712256841
transform 1 0 3104 0 1 770
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1712256841
transform 1 0 3096 0 1 770
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1712256841
transform 1 0 3088 0 1 770
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1712256841
transform 1 0 2984 0 1 770
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1712256841
transform 1 0 2976 0 1 770
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1712256841
transform 1 0 2832 0 1 770
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1712256841
transform 1 0 2824 0 1 770
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1712256841
transform 1 0 2816 0 1 770
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1712256841
transform 1 0 2712 0 1 770
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1712256841
transform 1 0 2704 0 1 770
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1712256841
transform 1 0 2696 0 1 770
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1712256841
transform 1 0 2688 0 1 770
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1712256841
transform 1 0 2656 0 1 770
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1712256841
transform 1 0 2632 0 1 770
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1712256841
transform 1 0 2624 0 1 770
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1712256841
transform 1 0 2592 0 1 770
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1712256841
transform 1 0 2584 0 1 770
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1712256841
transform 1 0 2576 0 1 770
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1712256841
transform 1 0 2568 0 1 770
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1712256841
transform 1 0 2560 0 1 770
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1712256841
transform 1 0 2552 0 1 770
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1712256841
transform 1 0 2544 0 1 770
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1712256841
transform 1 0 2496 0 1 770
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1712256841
transform 1 0 2488 0 1 770
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1712256841
transform 1 0 2480 0 1 770
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1712256841
transform 1 0 2472 0 1 770
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1712256841
transform 1 0 2448 0 1 770
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1712256841
transform 1 0 2440 0 1 770
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1712256841
transform 1 0 2432 0 1 770
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1712256841
transform 1 0 2400 0 1 770
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1712256841
transform 1 0 2392 0 1 770
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1712256841
transform 1 0 2368 0 1 770
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1712256841
transform 1 0 2360 0 1 770
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1712256841
transform 1 0 2352 0 1 770
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1712256841
transform 1 0 2344 0 1 770
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1712256841
transform 1 0 2336 0 1 770
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1712256841
transform 1 0 2296 0 1 770
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1712256841
transform 1 0 2288 0 1 770
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1712256841
transform 1 0 2280 0 1 770
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1712256841
transform 1 0 2272 0 1 770
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1712256841
transform 1 0 2264 0 1 770
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1712256841
transform 1 0 2224 0 1 770
box -8 -3 16 105
use FILL  FILL_3926
timestamp 1712256841
transform 1 0 2216 0 1 770
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1712256841
transform 1 0 2208 0 1 770
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1712256841
transform 1 0 2200 0 1 770
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1712256841
transform 1 0 2192 0 1 770
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1712256841
transform 1 0 2160 0 1 770
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1712256841
transform 1 0 2152 0 1 770
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1712256841
transform 1 0 2144 0 1 770
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1712256841
transform 1 0 2112 0 1 770
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1712256841
transform 1 0 2104 0 1 770
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1712256841
transform 1 0 2096 0 1 770
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1712256841
transform 1 0 2088 0 1 770
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1712256841
transform 1 0 2080 0 1 770
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1712256841
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1712256841
transform 1 0 2024 0 1 770
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1712256841
transform 1 0 2016 0 1 770
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1712256841
transform 1 0 2008 0 1 770
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1712256841
transform 1 0 2000 0 1 770
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1712256841
transform 1 0 1992 0 1 770
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1712256841
transform 1 0 1952 0 1 770
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1712256841
transform 1 0 1944 0 1 770
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1712256841
transform 1 0 1936 0 1 770
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1712256841
transform 1 0 1928 0 1 770
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1712256841
transform 1 0 1920 0 1 770
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1712256841
transform 1 0 1880 0 1 770
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1712256841
transform 1 0 1872 0 1 770
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1712256841
transform 1 0 1864 0 1 770
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1712256841
transform 1 0 1856 0 1 770
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1712256841
transform 1 0 1848 0 1 770
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1712256841
transform 1 0 1808 0 1 770
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1712256841
transform 1 0 1800 0 1 770
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1712256841
transform 1 0 1792 0 1 770
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1712256841
transform 1 0 1784 0 1 770
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1712256841
transform 1 0 1776 0 1 770
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1712256841
transform 1 0 1744 0 1 770
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1712256841
transform 1 0 1736 0 1 770
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1712256841
transform 1 0 1728 0 1 770
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1712256841
transform 1 0 1696 0 1 770
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1712256841
transform 1 0 1688 0 1 770
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1712256841
transform 1 0 1680 0 1 770
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1712256841
transform 1 0 1672 0 1 770
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1712256841
transform 1 0 1664 0 1 770
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1712256841
transform 1 0 1624 0 1 770
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1712256841
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1712256841
transform 1 0 1608 0 1 770
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1712256841
transform 1 0 1600 0 1 770
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1712256841
transform 1 0 1592 0 1 770
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1712256841
transform 1 0 1584 0 1 770
box -8 -3 16 105
use FILL  FILL_3973
timestamp 1712256841
transform 1 0 1536 0 1 770
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1712256841
transform 1 0 1528 0 1 770
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1712256841
transform 1 0 1520 0 1 770
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1712256841
transform 1 0 1512 0 1 770
box -8 -3 16 105
use FILL  FILL_3977
timestamp 1712256841
transform 1 0 1504 0 1 770
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1712256841
transform 1 0 1496 0 1 770
box -8 -3 16 105
use FILL  FILL_3979
timestamp 1712256841
transform 1 0 1456 0 1 770
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1712256841
transform 1 0 1448 0 1 770
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1712256841
transform 1 0 1424 0 1 770
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1712256841
transform 1 0 1416 0 1 770
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1712256841
transform 1 0 1408 0 1 770
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1712256841
transform 1 0 1400 0 1 770
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1712256841
transform 1 0 1392 0 1 770
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1712256841
transform 1 0 1344 0 1 770
box -8 -3 16 105
use FILL  FILL_3987
timestamp 1712256841
transform 1 0 1336 0 1 770
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1712256841
transform 1 0 1328 0 1 770
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1712256841
transform 1 0 1320 0 1 770
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1712256841
transform 1 0 1312 0 1 770
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1712256841
transform 1 0 1264 0 1 770
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1712256841
transform 1 0 1256 0 1 770
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1712256841
transform 1 0 1248 0 1 770
box -8 -3 16 105
use FILL  FILL_3994
timestamp 1712256841
transform 1 0 1240 0 1 770
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1712256841
transform 1 0 1208 0 1 770
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1712256841
transform 1 0 1200 0 1 770
box -8 -3 16 105
use FILL  FILL_3997
timestamp 1712256841
transform 1 0 1192 0 1 770
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1712256841
transform 1 0 1184 0 1 770
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1712256841
transform 1 0 1176 0 1 770
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1712256841
transform 1 0 1128 0 1 770
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1712256841
transform 1 0 1120 0 1 770
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1712256841
transform 1 0 1112 0 1 770
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1712256841
transform 1 0 1088 0 1 770
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1712256841
transform 1 0 1080 0 1 770
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1712256841
transform 1 0 1072 0 1 770
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1712256841
transform 1 0 1064 0 1 770
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1712256841
transform 1 0 1024 0 1 770
box -8 -3 16 105
use FILL  FILL_4008
timestamp 1712256841
transform 1 0 1016 0 1 770
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1712256841
transform 1 0 1008 0 1 770
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1712256841
transform 1 0 968 0 1 770
box -8 -3 16 105
use FILL  FILL_4011
timestamp 1712256841
transform 1 0 960 0 1 770
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1712256841
transform 1 0 952 0 1 770
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1712256841
transform 1 0 944 0 1 770
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1712256841
transform 1 0 936 0 1 770
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1712256841
transform 1 0 896 0 1 770
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1712256841
transform 1 0 888 0 1 770
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1712256841
transform 1 0 848 0 1 770
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1712256841
transform 1 0 840 0 1 770
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1712256841
transform 1 0 832 0 1 770
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1712256841
transform 1 0 824 0 1 770
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1712256841
transform 1 0 816 0 1 770
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1712256841
transform 1 0 808 0 1 770
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1712256841
transform 1 0 800 0 1 770
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1712256841
transform 1 0 736 0 1 770
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1712256841
transform 1 0 728 0 1 770
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1712256841
transform 1 0 720 0 1 770
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1712256841
transform 1 0 712 0 1 770
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1712256841
transform 1 0 704 0 1 770
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1712256841
transform 1 0 696 0 1 770
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1712256841
transform 1 0 656 0 1 770
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1712256841
transform 1 0 648 0 1 770
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1712256841
transform 1 0 640 0 1 770
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1712256841
transform 1 0 592 0 1 770
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1712256841
transform 1 0 584 0 1 770
box -8 -3 16 105
use FILL  FILL_4035
timestamp 1712256841
transform 1 0 576 0 1 770
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1712256841
transform 1 0 568 0 1 770
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1712256841
transform 1 0 560 0 1 770
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1712256841
transform 1 0 552 0 1 770
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1712256841
transform 1 0 504 0 1 770
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1712256841
transform 1 0 496 0 1 770
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1712256841
transform 1 0 488 0 1 770
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1712256841
transform 1 0 480 0 1 770
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1712256841
transform 1 0 472 0 1 770
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1712256841
transform 1 0 424 0 1 770
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1712256841
transform 1 0 416 0 1 770
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1712256841
transform 1 0 408 0 1 770
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1712256841
transform 1 0 400 0 1 770
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1712256841
transform 1 0 392 0 1 770
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1712256841
transform 1 0 344 0 1 770
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1712256841
transform 1 0 336 0 1 770
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1712256841
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1712256841
transform 1 0 320 0 1 770
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1712256841
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1712256841
transform 1 0 272 0 1 770
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1712256841
transform 1 0 264 0 1 770
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1712256841
transform 1 0 256 0 1 770
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1712256841
transform 1 0 216 0 1 770
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1712256841
transform 1 0 208 0 1 770
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1712256841
transform 1 0 200 0 1 770
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1712256841
transform 1 0 192 0 1 770
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1712256841
transform 1 0 184 0 1 770
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1712256841
transform 1 0 136 0 1 770
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1712256841
transform 1 0 128 0 1 770
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1712256841
transform 1 0 120 0 1 770
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1712256841
transform 1 0 112 0 1 770
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1712256841
transform 1 0 80 0 1 770
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1712256841
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1712256841
transform 1 0 3424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1712256841
transform 1 0 3400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1712256841
transform 1 0 3392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1712256841
transform 1 0 3384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4072
timestamp 1712256841
transform 1 0 3376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1712256841
transform 1 0 3312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1712256841
transform 1 0 3224 0 -1 770
box -8 -3 16 105
use FILL  FILL_4075
timestamp 1712256841
transform 1 0 3184 0 -1 770
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1712256841
transform 1 0 3176 0 -1 770
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1712256841
transform 1 0 3168 0 -1 770
box -8 -3 16 105
use FILL  FILL_4078
timestamp 1712256841
transform 1 0 3160 0 -1 770
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1712256841
transform 1 0 3120 0 -1 770
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1712256841
transform 1 0 3088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1712256841
transform 1 0 3080 0 -1 770
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1712256841
transform 1 0 3072 0 -1 770
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1712256841
transform 1 0 3008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1712256841
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1712256841
transform 1 0 2952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1712256841
transform 1 0 2944 0 -1 770
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1712256841
transform 1 0 2896 0 -1 770
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1712256841
transform 1 0 2888 0 -1 770
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1712256841
transform 1 0 2880 0 -1 770
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1712256841
transform 1 0 2872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4091
timestamp 1712256841
transform 1 0 2864 0 -1 770
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1712256841
transform 1 0 2776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1712256841
transform 1 0 2672 0 -1 770
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1712256841
transform 1 0 2664 0 -1 770
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1712256841
transform 1 0 2656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1712256841
transform 1 0 2600 0 -1 770
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1712256841
transform 1 0 2592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1712256841
transform 1 0 2560 0 -1 770
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1712256841
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1712256841
transform 1 0 2528 0 -1 770
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1712256841
transform 1 0 2520 0 -1 770
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1712256841
transform 1 0 2480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4103
timestamp 1712256841
transform 1 0 2472 0 -1 770
box -8 -3 16 105
use FILL  FILL_4104
timestamp 1712256841
transform 1 0 2464 0 -1 770
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1712256841
transform 1 0 2456 0 -1 770
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1712256841
transform 1 0 2408 0 -1 770
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1712256841
transform 1 0 2400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1712256841
transform 1 0 2392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1712256841
transform 1 0 2384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4110
timestamp 1712256841
transform 1 0 2336 0 -1 770
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1712256841
transform 1 0 2328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1712256841
transform 1 0 2320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4113
timestamp 1712256841
transform 1 0 2272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1712256841
transform 1 0 2264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1712256841
transform 1 0 2256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1712256841
transform 1 0 2248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1712256841
transform 1 0 2200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1712256841
transform 1 0 2192 0 -1 770
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1712256841
transform 1 0 2184 0 -1 770
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1712256841
transform 1 0 2176 0 -1 770
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1712256841
transform 1 0 2128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4122
timestamp 1712256841
transform 1 0 2120 0 -1 770
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1712256841
transform 1 0 2112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1712256841
transform 1 0 2072 0 -1 770
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1712256841
transform 1 0 2064 0 -1 770
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1712256841
transform 1 0 2056 0 -1 770
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1712256841
transform 1 0 2048 0 -1 770
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1712256841
transform 1 0 2008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1712256841
transform 1 0 2000 0 -1 770
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1712256841
transform 1 0 1992 0 -1 770
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1712256841
transform 1 0 1952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1712256841
transform 1 0 1944 0 -1 770
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1712256841
transform 1 0 1936 0 -1 770
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1712256841
transform 1 0 1912 0 -1 770
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1712256841
transform 1 0 1904 0 -1 770
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1712256841
transform 1 0 1864 0 -1 770
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1712256841
transform 1 0 1856 0 -1 770
box -8 -3 16 105
use FILL  FILL_4138
timestamp 1712256841
transform 1 0 1848 0 -1 770
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1712256841
transform 1 0 1816 0 -1 770
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1712256841
transform 1 0 1808 0 -1 770
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1712256841
transform 1 0 1800 0 -1 770
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1712256841
transform 1 0 1776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1712256841
transform 1 0 1736 0 -1 770
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1712256841
transform 1 0 1728 0 -1 770
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1712256841
transform 1 0 1720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1712256841
transform 1 0 1712 0 -1 770
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1712256841
transform 1 0 1704 0 -1 770
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1712256841
transform 1 0 1664 0 -1 770
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1712256841
transform 1 0 1656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1712256841
transform 1 0 1648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1712256841
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1712256841
transform 1 0 1600 0 -1 770
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1712256841
transform 1 0 1592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4154
timestamp 1712256841
transform 1 0 1552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1712256841
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1712256841
transform 1 0 1520 0 -1 770
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1712256841
transform 1 0 1488 0 -1 770
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1712256841
transform 1 0 1480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1712256841
transform 1 0 1472 0 -1 770
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1712256841
transform 1 0 1432 0 -1 770
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1712256841
transform 1 0 1424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1712256841
transform 1 0 1416 0 -1 770
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1712256841
transform 1 0 1376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1712256841
transform 1 0 1368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4165
timestamp 1712256841
transform 1 0 1360 0 -1 770
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1712256841
transform 1 0 1352 0 -1 770
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1712256841
transform 1 0 1312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1712256841
transform 1 0 1304 0 -1 770
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1712256841
transform 1 0 1264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1712256841
transform 1 0 1256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1712256841
transform 1 0 1248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1712256841
transform 1 0 1240 0 -1 770
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1712256841
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1712256841
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1712256841
transform 1 0 1152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1712256841
transform 1 0 1144 0 -1 770
box -8 -3 16 105
use FILL  FILL_4177
timestamp 1712256841
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1712256841
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1712256841
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1712256841
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1712256841
transform 1 0 1048 0 -1 770
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1712256841
transform 1 0 1040 0 -1 770
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1712256841
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1712256841
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1712256841
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use FILL  FILL_4186
timestamp 1712256841
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1712256841
transform 1 0 944 0 -1 770
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1712256841
transform 1 0 936 0 -1 770
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1712256841
transform 1 0 928 0 -1 770
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1712256841
transform 1 0 920 0 -1 770
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1712256841
transform 1 0 912 0 -1 770
box -8 -3 16 105
use FILL  FILL_4192
timestamp 1712256841
transform 1 0 904 0 -1 770
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1712256841
transform 1 0 840 0 -1 770
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1712256841
transform 1 0 832 0 -1 770
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1712256841
transform 1 0 824 0 -1 770
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1712256841
transform 1 0 816 0 -1 770
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1712256841
transform 1 0 792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1712256841
transform 1 0 784 0 -1 770
box -8 -3 16 105
use FILL  FILL_4199
timestamp 1712256841
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1712256841
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1712256841
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1712256841
transform 1 0 688 0 -1 770
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1712256841
transform 1 0 680 0 -1 770
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1712256841
transform 1 0 672 0 -1 770
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1712256841
transform 1 0 664 0 -1 770
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1712256841
transform 1 0 616 0 -1 770
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1712256841
transform 1 0 608 0 -1 770
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1712256841
transform 1 0 600 0 -1 770
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1712256841
transform 1 0 592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1712256841
transform 1 0 544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4211
timestamp 1712256841
transform 1 0 536 0 -1 770
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1712256841
transform 1 0 528 0 -1 770
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1712256841
transform 1 0 488 0 -1 770
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1712256841
transform 1 0 480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1712256841
transform 1 0 472 0 -1 770
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1712256841
transform 1 0 464 0 -1 770
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1712256841
transform 1 0 432 0 -1 770
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1712256841
transform 1 0 384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1712256841
transform 1 0 376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1712256841
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4221
timestamp 1712256841
transform 1 0 360 0 -1 770
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1712256841
transform 1 0 352 0 -1 770
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1712256841
transform 1 0 344 0 -1 770
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1712256841
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1712256841
transform 1 0 280 0 -1 770
box -8 -3 16 105
use FILL  FILL_4226
timestamp 1712256841
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1712256841
transform 1 0 264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1712256841
transform 1 0 256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1712256841
transform 1 0 192 0 -1 770
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1712256841
transform 1 0 184 0 -1 770
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1712256841
transform 1 0 176 0 -1 770
box -8 -3 16 105
use FILL  FILL_4232
timestamp 1712256841
transform 1 0 168 0 -1 770
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1712256841
transform 1 0 160 0 -1 770
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1712256841
transform 1 0 152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1712256841
transform 1 0 144 0 -1 770
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1712256841
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1712256841
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1712256841
transform 1 0 3424 0 1 570
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1712256841
transform 1 0 3416 0 1 570
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1712256841
transform 1 0 3408 0 1 570
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1712256841
transform 1 0 3360 0 1 570
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1712256841
transform 1 0 3352 0 1 570
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1712256841
transform 1 0 3344 0 1 570
box -8 -3 16 105
use FILL  FILL_4244
timestamp 1712256841
transform 1 0 3336 0 1 570
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1712256841
transform 1 0 3328 0 1 570
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1712256841
transform 1 0 3288 0 1 570
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1712256841
transform 1 0 3280 0 1 570
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1712256841
transform 1 0 3240 0 1 570
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1712256841
transform 1 0 3232 0 1 570
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1712256841
transform 1 0 3224 0 1 570
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1712256841
transform 1 0 3216 0 1 570
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1712256841
transform 1 0 3208 0 1 570
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1712256841
transform 1 0 3200 0 1 570
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1712256841
transform 1 0 3192 0 1 570
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1712256841
transform 1 0 3144 0 1 570
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1712256841
transform 1 0 3136 0 1 570
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1712256841
transform 1 0 3128 0 1 570
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1712256841
transform 1 0 3104 0 1 570
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1712256841
transform 1 0 3096 0 1 570
box -8 -3 16 105
use FILL  FILL_4260
timestamp 1712256841
transform 1 0 3088 0 1 570
box -8 -3 16 105
use FILL  FILL_4261
timestamp 1712256841
transform 1 0 3080 0 1 570
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1712256841
transform 1 0 3072 0 1 570
box -8 -3 16 105
use FILL  FILL_4263
timestamp 1712256841
transform 1 0 3064 0 1 570
box -8 -3 16 105
use FILL  FILL_4264
timestamp 1712256841
transform 1 0 3008 0 1 570
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1712256841
transform 1 0 3000 0 1 570
box -8 -3 16 105
use FILL  FILL_4266
timestamp 1712256841
transform 1 0 2992 0 1 570
box -8 -3 16 105
use FILL  FILL_4267
timestamp 1712256841
transform 1 0 2984 0 1 570
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1712256841
transform 1 0 2976 0 1 570
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1712256841
transform 1 0 2968 0 1 570
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1712256841
transform 1 0 2928 0 1 570
box -8 -3 16 105
use FILL  FILL_4271
timestamp 1712256841
transform 1 0 2904 0 1 570
box -8 -3 16 105
use FILL  FILL_4272
timestamp 1712256841
transform 1 0 2896 0 1 570
box -8 -3 16 105
use FILL  FILL_4273
timestamp 1712256841
transform 1 0 2888 0 1 570
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1712256841
transform 1 0 2880 0 1 570
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1712256841
transform 1 0 2872 0 1 570
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1712256841
transform 1 0 2824 0 1 570
box -8 -3 16 105
use FILL  FILL_4277
timestamp 1712256841
transform 1 0 2816 0 1 570
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1712256841
transform 1 0 2808 0 1 570
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1712256841
transform 1 0 2800 0 1 570
box -8 -3 16 105
use FILL  FILL_4280
timestamp 1712256841
transform 1 0 2768 0 1 570
box -8 -3 16 105
use FILL  FILL_4281
timestamp 1712256841
transform 1 0 2760 0 1 570
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1712256841
transform 1 0 2752 0 1 570
box -8 -3 16 105
use FILL  FILL_4283
timestamp 1712256841
transform 1 0 2720 0 1 570
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1712256841
transform 1 0 2680 0 1 570
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1712256841
transform 1 0 2672 0 1 570
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1712256841
transform 1 0 2664 0 1 570
box -8 -3 16 105
use FILL  FILL_4287
timestamp 1712256841
transform 1 0 2656 0 1 570
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1712256841
transform 1 0 2608 0 1 570
box -8 -3 16 105
use FILL  FILL_4289
timestamp 1712256841
transform 1 0 2600 0 1 570
box -8 -3 16 105
use FILL  FILL_4290
timestamp 1712256841
transform 1 0 2592 0 1 570
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1712256841
transform 1 0 2560 0 1 570
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1712256841
transform 1 0 2552 0 1 570
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1712256841
transform 1 0 2544 0 1 570
box -8 -3 16 105
use FILL  FILL_4294
timestamp 1712256841
transform 1 0 2496 0 1 570
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1712256841
transform 1 0 2488 0 1 570
box -8 -3 16 105
use FILL  FILL_4296
timestamp 1712256841
transform 1 0 2480 0 1 570
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1712256841
transform 1 0 2472 0 1 570
box -8 -3 16 105
use FILL  FILL_4298
timestamp 1712256841
transform 1 0 2440 0 1 570
box -8 -3 16 105
use FILL  FILL_4299
timestamp 1712256841
transform 1 0 2432 0 1 570
box -8 -3 16 105
use FILL  FILL_4300
timestamp 1712256841
transform 1 0 2392 0 1 570
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1712256841
transform 1 0 2384 0 1 570
box -8 -3 16 105
use FILL  FILL_4302
timestamp 1712256841
transform 1 0 2376 0 1 570
box -8 -3 16 105
use FILL  FILL_4303
timestamp 1712256841
transform 1 0 2368 0 1 570
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1712256841
transform 1 0 2328 0 1 570
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1712256841
transform 1 0 2320 0 1 570
box -8 -3 16 105
use FILL  FILL_4306
timestamp 1712256841
transform 1 0 2280 0 1 570
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1712256841
transform 1 0 2272 0 1 570
box -8 -3 16 105
use FILL  FILL_4308
timestamp 1712256841
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_4309
timestamp 1712256841
transform 1 0 2256 0 1 570
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1712256841
transform 1 0 2208 0 1 570
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1712256841
transform 1 0 2200 0 1 570
box -8 -3 16 105
use FILL  FILL_4312
timestamp 1712256841
transform 1 0 2192 0 1 570
box -8 -3 16 105
use FILL  FILL_4313
timestamp 1712256841
transform 1 0 2160 0 1 570
box -8 -3 16 105
use FILL  FILL_4314
timestamp 1712256841
transform 1 0 2152 0 1 570
box -8 -3 16 105
use FILL  FILL_4315
timestamp 1712256841
transform 1 0 2120 0 1 570
box -8 -3 16 105
use FILL  FILL_4316
timestamp 1712256841
transform 1 0 2112 0 1 570
box -8 -3 16 105
use FILL  FILL_4317
timestamp 1712256841
transform 1 0 2072 0 1 570
box -8 -3 16 105
use FILL  FILL_4318
timestamp 1712256841
transform 1 0 2064 0 1 570
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1712256841
transform 1 0 2056 0 1 570
box -8 -3 16 105
use FILL  FILL_4320
timestamp 1712256841
transform 1 0 2048 0 1 570
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1712256841
transform 1 0 2008 0 1 570
box -8 -3 16 105
use FILL  FILL_4322
timestamp 1712256841
transform 1 0 2000 0 1 570
box -8 -3 16 105
use FILL  FILL_4323
timestamp 1712256841
transform 1 0 1992 0 1 570
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1712256841
transform 1 0 1960 0 1 570
box -8 -3 16 105
use FILL  FILL_4325
timestamp 1712256841
transform 1 0 1952 0 1 570
box -8 -3 16 105
use FILL  FILL_4326
timestamp 1712256841
transform 1 0 1920 0 1 570
box -8 -3 16 105
use FILL  FILL_4327
timestamp 1712256841
transform 1 0 1912 0 1 570
box -8 -3 16 105
use FILL  FILL_4328
timestamp 1712256841
transform 1 0 1904 0 1 570
box -8 -3 16 105
use FILL  FILL_4329
timestamp 1712256841
transform 1 0 1848 0 1 570
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1712256841
transform 1 0 1840 0 1 570
box -8 -3 16 105
use FILL  FILL_4331
timestamp 1712256841
transform 1 0 1832 0 1 570
box -8 -3 16 105
use FILL  FILL_4332
timestamp 1712256841
transform 1 0 1824 0 1 570
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1712256841
transform 1 0 1816 0 1 570
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1712256841
transform 1 0 1808 0 1 570
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1712256841
transform 1 0 1752 0 1 570
box -8 -3 16 105
use FILL  FILL_4336
timestamp 1712256841
transform 1 0 1744 0 1 570
box -8 -3 16 105
use FILL  FILL_4337
timestamp 1712256841
transform 1 0 1736 0 1 570
box -8 -3 16 105
use FILL  FILL_4338
timestamp 1712256841
transform 1 0 1712 0 1 570
box -8 -3 16 105
use FILL  FILL_4339
timestamp 1712256841
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1712256841
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_4341
timestamp 1712256841
transform 1 0 1656 0 1 570
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1712256841
transform 1 0 1648 0 1 570
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1712256841
transform 1 0 1608 0 1 570
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1712256841
transform 1 0 1576 0 1 570
box -8 -3 16 105
use FILL  FILL_4345
timestamp 1712256841
transform 1 0 1568 0 1 570
box -8 -3 16 105
use FILL  FILL_4346
timestamp 1712256841
transform 1 0 1560 0 1 570
box -8 -3 16 105
use FILL  FILL_4347
timestamp 1712256841
transform 1 0 1552 0 1 570
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1712256841
transform 1 0 1544 0 1 570
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1712256841
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1712256841
transform 1 0 1480 0 1 570
box -8 -3 16 105
use FILL  FILL_4351
timestamp 1712256841
transform 1 0 1472 0 1 570
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1712256841
transform 1 0 1464 0 1 570
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1712256841
transform 1 0 1456 0 1 570
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1712256841
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_4355
timestamp 1712256841
transform 1 0 1392 0 1 570
box -8 -3 16 105
use FILL  FILL_4356
timestamp 1712256841
transform 1 0 1384 0 1 570
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1712256841
transform 1 0 1376 0 1 570
box -8 -3 16 105
use FILL  FILL_4358
timestamp 1712256841
transform 1 0 1336 0 1 570
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1712256841
transform 1 0 1328 0 1 570
box -8 -3 16 105
use FILL  FILL_4360
timestamp 1712256841
transform 1 0 1288 0 1 570
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1712256841
transform 1 0 1280 0 1 570
box -8 -3 16 105
use FILL  FILL_4362
timestamp 1712256841
transform 1 0 1272 0 1 570
box -8 -3 16 105
use FILL  FILL_4363
timestamp 1712256841
transform 1 0 1264 0 1 570
box -8 -3 16 105
use FILL  FILL_4364
timestamp 1712256841
transform 1 0 1256 0 1 570
box -8 -3 16 105
use FILL  FILL_4365
timestamp 1712256841
transform 1 0 1216 0 1 570
box -8 -3 16 105
use FILL  FILL_4366
timestamp 1712256841
transform 1 0 1208 0 1 570
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1712256841
transform 1 0 1168 0 1 570
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1712256841
transform 1 0 1160 0 1 570
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1712256841
transform 1 0 1152 0 1 570
box -8 -3 16 105
use FILL  FILL_4370
timestamp 1712256841
transform 1 0 1144 0 1 570
box -8 -3 16 105
use FILL  FILL_4371
timestamp 1712256841
transform 1 0 1136 0 1 570
box -8 -3 16 105
use FILL  FILL_4372
timestamp 1712256841
transform 1 0 1088 0 1 570
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1712256841
transform 1 0 1080 0 1 570
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1712256841
transform 1 0 1072 0 1 570
box -8 -3 16 105
use FILL  FILL_4375
timestamp 1712256841
transform 1 0 1064 0 1 570
box -8 -3 16 105
use FILL  FILL_4376
timestamp 1712256841
transform 1 0 992 0 1 570
box -8 -3 16 105
use FILL  FILL_4377
timestamp 1712256841
transform 1 0 984 0 1 570
box -8 -3 16 105
use FILL  FILL_4378
timestamp 1712256841
transform 1 0 976 0 1 570
box -8 -3 16 105
use FILL  FILL_4379
timestamp 1712256841
transform 1 0 936 0 1 570
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1712256841
transform 1 0 928 0 1 570
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1712256841
transform 1 0 920 0 1 570
box -8 -3 16 105
use FILL  FILL_4382
timestamp 1712256841
transform 1 0 912 0 1 570
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1712256841
transform 1 0 872 0 1 570
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1712256841
transform 1 0 864 0 1 570
box -8 -3 16 105
use FILL  FILL_4385
timestamp 1712256841
transform 1 0 856 0 1 570
box -8 -3 16 105
use FILL  FILL_4386
timestamp 1712256841
transform 1 0 816 0 1 570
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1712256841
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1712256841
transform 1 0 800 0 1 570
box -8 -3 16 105
use FILL  FILL_4389
timestamp 1712256841
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_4390
timestamp 1712256841
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_4391
timestamp 1712256841
transform 1 0 744 0 1 570
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1712256841
transform 1 0 720 0 1 570
box -8 -3 16 105
use FILL  FILL_4393
timestamp 1712256841
transform 1 0 712 0 1 570
box -8 -3 16 105
use FILL  FILL_4394
timestamp 1712256841
transform 1 0 704 0 1 570
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1712256841
transform 1 0 696 0 1 570
box -8 -3 16 105
use FILL  FILL_4396
timestamp 1712256841
transform 1 0 656 0 1 570
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1712256841
transform 1 0 648 0 1 570
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1712256841
transform 1 0 640 0 1 570
box -8 -3 16 105
use FILL  FILL_4399
timestamp 1712256841
transform 1 0 600 0 1 570
box -8 -3 16 105
use FILL  FILL_4400
timestamp 1712256841
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1712256841
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1712256841
transform 1 0 576 0 1 570
box -8 -3 16 105
use FILL  FILL_4403
timestamp 1712256841
transform 1 0 568 0 1 570
box -8 -3 16 105
use FILL  FILL_4404
timestamp 1712256841
transform 1 0 528 0 1 570
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1712256841
transform 1 0 520 0 1 570
box -8 -3 16 105
use FILL  FILL_4406
timestamp 1712256841
transform 1 0 512 0 1 570
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1712256841
transform 1 0 504 0 1 570
box -8 -3 16 105
use FILL  FILL_4408
timestamp 1712256841
transform 1 0 480 0 1 570
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1712256841
transform 1 0 472 0 1 570
box -8 -3 16 105
use FILL  FILL_4410
timestamp 1712256841
transform 1 0 424 0 1 570
box -8 -3 16 105
use FILL  FILL_4411
timestamp 1712256841
transform 1 0 416 0 1 570
box -8 -3 16 105
use FILL  FILL_4412
timestamp 1712256841
transform 1 0 408 0 1 570
box -8 -3 16 105
use FILL  FILL_4413
timestamp 1712256841
transform 1 0 400 0 1 570
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1712256841
transform 1 0 392 0 1 570
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1712256841
transform 1 0 384 0 1 570
box -8 -3 16 105
use FILL  FILL_4416
timestamp 1712256841
transform 1 0 336 0 1 570
box -8 -3 16 105
use FILL  FILL_4417
timestamp 1712256841
transform 1 0 328 0 1 570
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1712256841
transform 1 0 320 0 1 570
box -8 -3 16 105
use FILL  FILL_4419
timestamp 1712256841
transform 1 0 312 0 1 570
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1712256841
transform 1 0 272 0 1 570
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1712256841
transform 1 0 264 0 1 570
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1712256841
transform 1 0 256 0 1 570
box -8 -3 16 105
use FILL  FILL_4423
timestamp 1712256841
transform 1 0 248 0 1 570
box -8 -3 16 105
use FILL  FILL_4424
timestamp 1712256841
transform 1 0 240 0 1 570
box -8 -3 16 105
use FILL  FILL_4425
timestamp 1712256841
transform 1 0 192 0 1 570
box -8 -3 16 105
use FILL  FILL_4426
timestamp 1712256841
transform 1 0 184 0 1 570
box -8 -3 16 105
use FILL  FILL_4427
timestamp 1712256841
transform 1 0 176 0 1 570
box -8 -3 16 105
use FILL  FILL_4428
timestamp 1712256841
transform 1 0 168 0 1 570
box -8 -3 16 105
use FILL  FILL_4429
timestamp 1712256841
transform 1 0 160 0 1 570
box -8 -3 16 105
use FILL  FILL_4430
timestamp 1712256841
transform 1 0 128 0 1 570
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1712256841
transform 1 0 120 0 1 570
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1712256841
transform 1 0 88 0 1 570
box -8 -3 16 105
use FILL  FILL_4433
timestamp 1712256841
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1712256841
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_4435
timestamp 1712256841
transform 1 0 3424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4436
timestamp 1712256841
transform 1 0 3384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4437
timestamp 1712256841
transform 1 0 3376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1712256841
transform 1 0 3368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4439
timestamp 1712256841
transform 1 0 3360 0 -1 570
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1712256841
transform 1 0 3320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4441
timestamp 1712256841
transform 1 0 3312 0 -1 570
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1712256841
transform 1 0 3272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1712256841
transform 1 0 3264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1712256841
transform 1 0 3256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4445
timestamp 1712256841
transform 1 0 3248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4446
timestamp 1712256841
transform 1 0 3208 0 -1 570
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1712256841
transform 1 0 3200 0 -1 570
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1712256841
transform 1 0 3160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4449
timestamp 1712256841
transform 1 0 3152 0 -1 570
box -8 -3 16 105
use FILL  FILL_4450
timestamp 1712256841
transform 1 0 3144 0 -1 570
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1712256841
transform 1 0 3136 0 -1 570
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1712256841
transform 1 0 3128 0 -1 570
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1712256841
transform 1 0 3088 0 -1 570
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1712256841
transform 1 0 3048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4455
timestamp 1712256841
transform 1 0 3040 0 -1 570
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1712256841
transform 1 0 3032 0 -1 570
box -8 -3 16 105
use FILL  FILL_4457
timestamp 1712256841
transform 1 0 3024 0 -1 570
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1712256841
transform 1 0 2976 0 -1 570
box -8 -3 16 105
use FILL  FILL_4459
timestamp 1712256841
transform 1 0 2968 0 -1 570
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1712256841
transform 1 0 2960 0 -1 570
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1712256841
transform 1 0 2920 0 -1 570
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1712256841
transform 1 0 2912 0 -1 570
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1712256841
transform 1 0 2904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4464
timestamp 1712256841
transform 1 0 2848 0 -1 570
box -8 -3 16 105
use FILL  FILL_4465
timestamp 1712256841
transform 1 0 2840 0 -1 570
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1712256841
transform 1 0 2832 0 -1 570
box -8 -3 16 105
use FILL  FILL_4467
timestamp 1712256841
transform 1 0 2824 0 -1 570
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1712256841
transform 1 0 2816 0 -1 570
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1712256841
transform 1 0 2768 0 -1 570
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1712256841
transform 1 0 2760 0 -1 570
box -8 -3 16 105
use FILL  FILL_4471
timestamp 1712256841
transform 1 0 2752 0 -1 570
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1712256841
transform 1 0 2744 0 -1 570
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1712256841
transform 1 0 2712 0 -1 570
box -8 -3 16 105
use FILL  FILL_4474
timestamp 1712256841
transform 1 0 2672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4475
timestamp 1712256841
transform 1 0 2664 0 -1 570
box -8 -3 16 105
use FILL  FILL_4476
timestamp 1712256841
transform 1 0 2656 0 -1 570
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1712256841
transform 1 0 2648 0 -1 570
box -8 -3 16 105
use FILL  FILL_4478
timestamp 1712256841
transform 1 0 2640 0 -1 570
box -8 -3 16 105
use FILL  FILL_4479
timestamp 1712256841
transform 1 0 2608 0 -1 570
box -8 -3 16 105
use FILL  FILL_4480
timestamp 1712256841
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1712256841
transform 1 0 2568 0 -1 570
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1712256841
transform 1 0 2560 0 -1 570
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1712256841
transform 1 0 2552 0 -1 570
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1712256841
transform 1 0 2528 0 -1 570
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1712256841
transform 1 0 2520 0 -1 570
box -8 -3 16 105
use FILL  FILL_4486
timestamp 1712256841
transform 1 0 2488 0 -1 570
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1712256841
transform 1 0 2480 0 -1 570
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1712256841
transform 1 0 2448 0 -1 570
box -8 -3 16 105
use FILL  FILL_4489
timestamp 1712256841
transform 1 0 2440 0 -1 570
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1712256841
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4491
timestamp 1712256841
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4492
timestamp 1712256841
transform 1 0 2376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1712256841
transform 1 0 2368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4494
timestamp 1712256841
transform 1 0 2336 0 -1 570
box -8 -3 16 105
use FILL  FILL_4495
timestamp 1712256841
transform 1 0 2328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4496
timestamp 1712256841
transform 1 0 2320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1712256841
transform 1 0 2312 0 -1 570
box -8 -3 16 105
use FILL  FILL_4498
timestamp 1712256841
transform 1 0 2264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1712256841
transform 1 0 2256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4500
timestamp 1712256841
transform 1 0 2248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4501
timestamp 1712256841
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1712256841
transform 1 0 2192 0 -1 570
box -8 -3 16 105
use FILL  FILL_4503
timestamp 1712256841
transform 1 0 2184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1712256841
transform 1 0 2176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4505
timestamp 1712256841
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1712256841
transform 1 0 2128 0 -1 570
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1712256841
transform 1 0 2120 0 -1 570
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1712256841
transform 1 0 2112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1712256841
transform 1 0 2064 0 -1 570
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1712256841
transform 1 0 2056 0 -1 570
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1712256841
transform 1 0 2048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4512
timestamp 1712256841
transform 1 0 2040 0 -1 570
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1712256841
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use FILL  FILL_4514
timestamp 1712256841
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use FILL  FILL_4515
timestamp 1712256841
transform 1 0 1976 0 -1 570
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1712256841
transform 1 0 1968 0 -1 570
box -8 -3 16 105
use FILL  FILL_4517
timestamp 1712256841
transform 1 0 1920 0 -1 570
box -8 -3 16 105
use FILL  FILL_4518
timestamp 1712256841
transform 1 0 1912 0 -1 570
box -8 -3 16 105
use FILL  FILL_4519
timestamp 1712256841
transform 1 0 1904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1712256841
transform 1 0 1864 0 -1 570
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1712256841
transform 1 0 1856 0 -1 570
box -8 -3 16 105
use FILL  FILL_4522
timestamp 1712256841
transform 1 0 1848 0 -1 570
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1712256841
transform 1 0 1800 0 -1 570
box -8 -3 16 105
use FILL  FILL_4524
timestamp 1712256841
transform 1 0 1792 0 -1 570
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1712256841
transform 1 0 1784 0 -1 570
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1712256841
transform 1 0 1744 0 -1 570
box -8 -3 16 105
use FILL  FILL_4527
timestamp 1712256841
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1712256841
transform 1 0 1728 0 -1 570
box -8 -3 16 105
use FILL  FILL_4529
timestamp 1712256841
transform 1 0 1688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1712256841
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4531
timestamp 1712256841
transform 1 0 1640 0 -1 570
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1712256841
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1712256841
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_4534
timestamp 1712256841
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1712256841
transform 1 0 1576 0 -1 570
box -8 -3 16 105
use FILL  FILL_4536
timestamp 1712256841
transform 1 0 1552 0 -1 570
box -8 -3 16 105
use FILL  FILL_4537
timestamp 1712256841
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_4538
timestamp 1712256841
transform 1 0 1504 0 -1 570
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1712256841
transform 1 0 1496 0 -1 570
box -8 -3 16 105
use FILL  FILL_4540
timestamp 1712256841
transform 1 0 1488 0 -1 570
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1712256841
transform 1 0 1440 0 -1 570
box -8 -3 16 105
use FILL  FILL_4542
timestamp 1712256841
transform 1 0 1432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1712256841
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1712256841
transform 1 0 1376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1712256841
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1712256841
transform 1 0 1360 0 -1 570
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1712256841
transform 1 0 1320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1712256841
transform 1 0 1288 0 -1 570
box -8 -3 16 105
use FILL  FILL_4549
timestamp 1712256841
transform 1 0 1280 0 -1 570
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1712256841
transform 1 0 1272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4551
timestamp 1712256841
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4552
timestamp 1712256841
transform 1 0 1208 0 -1 570
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1712256841
transform 1 0 1200 0 -1 570
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1712256841
transform 1 0 1192 0 -1 570
box -8 -3 16 105
use FILL  FILL_4555
timestamp 1712256841
transform 1 0 1184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4556
timestamp 1712256841
transform 1 0 1152 0 -1 570
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1712256841
transform 1 0 1144 0 -1 570
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1712256841
transform 1 0 1136 0 -1 570
box -8 -3 16 105
use FILL  FILL_4559
timestamp 1712256841
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use FILL  FILL_4560
timestamp 1712256841
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_4561
timestamp 1712256841
transform 1 0 1048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4562
timestamp 1712256841
transform 1 0 1040 0 -1 570
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1712256841
transform 1 0 1032 0 -1 570
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1712256841
transform 1 0 1024 0 -1 570
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1712256841
transform 1 0 976 0 -1 570
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1712256841
transform 1 0 968 0 -1 570
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1712256841
transform 1 0 960 0 -1 570
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1712256841
transform 1 0 912 0 -1 570
box -8 -3 16 105
use FILL  FILL_4569
timestamp 1712256841
transform 1 0 904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4570
timestamp 1712256841
transform 1 0 864 0 -1 570
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1712256841
transform 1 0 856 0 -1 570
box -8 -3 16 105
use FILL  FILL_4572
timestamp 1712256841
transform 1 0 848 0 -1 570
box -8 -3 16 105
use FILL  FILL_4573
timestamp 1712256841
transform 1 0 800 0 -1 570
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1712256841
transform 1 0 792 0 -1 570
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1712256841
transform 1 0 784 0 -1 570
box -8 -3 16 105
use FILL  FILL_4576
timestamp 1712256841
transform 1 0 744 0 -1 570
box -8 -3 16 105
use FILL  FILL_4577
timestamp 1712256841
transform 1 0 736 0 -1 570
box -8 -3 16 105
use FILL  FILL_4578
timestamp 1712256841
transform 1 0 728 0 -1 570
box -8 -3 16 105
use FILL  FILL_4579
timestamp 1712256841
transform 1 0 688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1712256841
transform 1 0 680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1712256841
transform 1 0 672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4582
timestamp 1712256841
transform 1 0 640 0 -1 570
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1712256841
transform 1 0 632 0 -1 570
box -8 -3 16 105
use FILL  FILL_4584
timestamp 1712256841
transform 1 0 600 0 -1 570
box -8 -3 16 105
use FILL  FILL_4585
timestamp 1712256841
transform 1 0 592 0 -1 570
box -8 -3 16 105
use FILL  FILL_4586
timestamp 1712256841
transform 1 0 584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1712256841
transform 1 0 536 0 -1 570
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1712256841
transform 1 0 528 0 -1 570
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1712256841
transform 1 0 520 0 -1 570
box -8 -3 16 105
use FILL  FILL_4590
timestamp 1712256841
transform 1 0 512 0 -1 570
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1712256841
transform 1 0 472 0 -1 570
box -8 -3 16 105
use FILL  FILL_4592
timestamp 1712256841
transform 1 0 464 0 -1 570
box -8 -3 16 105
use FILL  FILL_4593
timestamp 1712256841
transform 1 0 456 0 -1 570
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1712256841
transform 1 0 416 0 -1 570
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1712256841
transform 1 0 408 0 -1 570
box -8 -3 16 105
use FILL  FILL_4596
timestamp 1712256841
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1712256841
transform 1 0 392 0 -1 570
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1712256841
transform 1 0 368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4599
timestamp 1712256841
transform 1 0 320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1712256841
transform 1 0 312 0 -1 570
box -8 -3 16 105
use FILL  FILL_4601
timestamp 1712256841
transform 1 0 304 0 -1 570
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1712256841
transform 1 0 296 0 -1 570
box -8 -3 16 105
use FILL  FILL_4603
timestamp 1712256841
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_4604
timestamp 1712256841
transform 1 0 248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4605
timestamp 1712256841
transform 1 0 240 0 -1 570
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1712256841
transform 1 0 192 0 -1 570
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1712256841
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1712256841
transform 1 0 176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1712256841
transform 1 0 168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1712256841
transform 1 0 160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1712256841
transform 1 0 128 0 -1 570
box -8 -3 16 105
use FILL  FILL_4612
timestamp 1712256841
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_4613
timestamp 1712256841
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1712256841
transform 1 0 3424 0 1 370
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1712256841
transform 1 0 3320 0 1 370
box -8 -3 16 105
use FILL  FILL_4616
timestamp 1712256841
transform 1 0 3216 0 1 370
box -8 -3 16 105
use FILL  FILL_4617
timestamp 1712256841
transform 1 0 3208 0 1 370
box -8 -3 16 105
use FILL  FILL_4618
timestamp 1712256841
transform 1 0 3104 0 1 370
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1712256841
transform 1 0 3096 0 1 370
box -8 -3 16 105
use FILL  FILL_4620
timestamp 1712256841
transform 1 0 3088 0 1 370
box -8 -3 16 105
use FILL  FILL_4621
timestamp 1712256841
transform 1 0 3080 0 1 370
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1712256841
transform 1 0 3032 0 1 370
box -8 -3 16 105
use FILL  FILL_4623
timestamp 1712256841
transform 1 0 3024 0 1 370
box -8 -3 16 105
use FILL  FILL_4624
timestamp 1712256841
transform 1 0 3016 0 1 370
box -8 -3 16 105
use FILL  FILL_4625
timestamp 1712256841
transform 1 0 2912 0 1 370
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1712256841
transform 1 0 2904 0 1 370
box -8 -3 16 105
use FILL  FILL_4627
timestamp 1712256841
transform 1 0 2896 0 1 370
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1712256841
transform 1 0 2792 0 1 370
box -8 -3 16 105
use FILL  FILL_4629
timestamp 1712256841
transform 1 0 2784 0 1 370
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1712256841
transform 1 0 2776 0 1 370
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1712256841
transform 1 0 2768 0 1 370
box -8 -3 16 105
use FILL  FILL_4632
timestamp 1712256841
transform 1 0 2760 0 1 370
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1712256841
transform 1 0 2752 0 1 370
box -8 -3 16 105
use FILL  FILL_4634
timestamp 1712256841
transform 1 0 2696 0 1 370
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1712256841
transform 1 0 2688 0 1 370
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1712256841
transform 1 0 2680 0 1 370
box -8 -3 16 105
use FILL  FILL_4637
timestamp 1712256841
transform 1 0 2672 0 1 370
box -8 -3 16 105
use FILL  FILL_4638
timestamp 1712256841
transform 1 0 2664 0 1 370
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1712256841
transform 1 0 2656 0 1 370
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1712256841
transform 1 0 2632 0 1 370
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1712256841
transform 1 0 2592 0 1 370
box -8 -3 16 105
use FILL  FILL_4642
timestamp 1712256841
transform 1 0 2584 0 1 370
box -8 -3 16 105
use FILL  FILL_4643
timestamp 1712256841
transform 1 0 2576 0 1 370
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1712256841
transform 1 0 2568 0 1 370
box -8 -3 16 105
use FILL  FILL_4645
timestamp 1712256841
transform 1 0 2560 0 1 370
box -8 -3 16 105
use FILL  FILL_4646
timestamp 1712256841
transform 1 0 2552 0 1 370
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1712256841
transform 1 0 2504 0 1 370
box -8 -3 16 105
use FILL  FILL_4648
timestamp 1712256841
transform 1 0 2496 0 1 370
box -8 -3 16 105
use FILL  FILL_4649
timestamp 1712256841
transform 1 0 2488 0 1 370
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1712256841
transform 1 0 2480 0 1 370
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1712256841
transform 1 0 2472 0 1 370
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1712256841
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_4653
timestamp 1712256841
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_4654
timestamp 1712256841
transform 1 0 2408 0 1 370
box -8 -3 16 105
use FILL  FILL_4655
timestamp 1712256841
transform 1 0 2400 0 1 370
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1712256841
transform 1 0 2368 0 1 370
box -8 -3 16 105
use FILL  FILL_4657
timestamp 1712256841
transform 1 0 2360 0 1 370
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1712256841
transform 1 0 2352 0 1 370
box -8 -3 16 105
use FILL  FILL_4659
timestamp 1712256841
transform 1 0 2344 0 1 370
box -8 -3 16 105
use FILL  FILL_4660
timestamp 1712256841
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1712256841
transform 1 0 2272 0 1 370
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1712256841
transform 1 0 2264 0 1 370
box -8 -3 16 105
use FILL  FILL_4663
timestamp 1712256841
transform 1 0 2256 0 1 370
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1712256841
transform 1 0 2248 0 1 370
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1712256841
transform 1 0 2240 0 1 370
box -8 -3 16 105
use FILL  FILL_4666
timestamp 1712256841
transform 1 0 2192 0 1 370
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1712256841
transform 1 0 2184 0 1 370
box -8 -3 16 105
use FILL  FILL_4668
timestamp 1712256841
transform 1 0 2176 0 1 370
box -8 -3 16 105
use FILL  FILL_4669
timestamp 1712256841
transform 1 0 2168 0 1 370
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1712256841
transform 1 0 2160 0 1 370
box -8 -3 16 105
use FILL  FILL_4671
timestamp 1712256841
transform 1 0 2112 0 1 370
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1712256841
transform 1 0 2104 0 1 370
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1712256841
transform 1 0 2096 0 1 370
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1712256841
transform 1 0 2088 0 1 370
box -8 -3 16 105
use FILL  FILL_4675
timestamp 1712256841
transform 1 0 2080 0 1 370
box -8 -3 16 105
use FILL  FILL_4676
timestamp 1712256841
transform 1 0 2032 0 1 370
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1712256841
transform 1 0 2024 0 1 370
box -8 -3 16 105
use FILL  FILL_4678
timestamp 1712256841
transform 1 0 2000 0 1 370
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1712256841
transform 1 0 1992 0 1 370
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1712256841
transform 1 0 1984 0 1 370
box -8 -3 16 105
use FILL  FILL_4681
timestamp 1712256841
transform 1 0 1976 0 1 370
box -8 -3 16 105
use FILL  FILL_4682
timestamp 1712256841
transform 1 0 1928 0 1 370
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1712256841
transform 1 0 1920 0 1 370
box -8 -3 16 105
use FILL  FILL_4684
timestamp 1712256841
transform 1 0 1912 0 1 370
box -8 -3 16 105
use FILL  FILL_4685
timestamp 1712256841
transform 1 0 1904 0 1 370
box -8 -3 16 105
use FILL  FILL_4686
timestamp 1712256841
transform 1 0 1864 0 1 370
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1712256841
transform 1 0 1856 0 1 370
box -8 -3 16 105
use FILL  FILL_4688
timestamp 1712256841
transform 1 0 1848 0 1 370
box -8 -3 16 105
use FILL  FILL_4689
timestamp 1712256841
transform 1 0 1816 0 1 370
box -8 -3 16 105
use FILL  FILL_4690
timestamp 1712256841
transform 1 0 1808 0 1 370
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1712256841
transform 1 0 1800 0 1 370
box -8 -3 16 105
use FILL  FILL_4692
timestamp 1712256841
transform 1 0 1760 0 1 370
box -8 -3 16 105
use FILL  FILL_4693
timestamp 1712256841
transform 1 0 1752 0 1 370
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1712256841
transform 1 0 1744 0 1 370
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1712256841
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_4696
timestamp 1712256841
transform 1 0 1688 0 1 370
box -8 -3 16 105
use FILL  FILL_4697
timestamp 1712256841
transform 1 0 1680 0 1 370
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1712256841
transform 1 0 1672 0 1 370
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1712256841
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1712256841
transform 1 0 1624 0 1 370
box -8 -3 16 105
use FILL  FILL_4701
timestamp 1712256841
transform 1 0 1616 0 1 370
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1712256841
transform 1 0 1576 0 1 370
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1712256841
transform 1 0 1568 0 1 370
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1712256841
transform 1 0 1536 0 1 370
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1712256841
transform 1 0 1528 0 1 370
box -8 -3 16 105
use FILL  FILL_4706
timestamp 1712256841
transform 1 0 1488 0 1 370
box -8 -3 16 105
use FILL  FILL_4707
timestamp 1712256841
transform 1 0 1480 0 1 370
box -8 -3 16 105
use FILL  FILL_4708
timestamp 1712256841
transform 1 0 1472 0 1 370
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1712256841
transform 1 0 1464 0 1 370
box -8 -3 16 105
use FILL  FILL_4710
timestamp 1712256841
transform 1 0 1432 0 1 370
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1712256841
transform 1 0 1392 0 1 370
box -8 -3 16 105
use FILL  FILL_4712
timestamp 1712256841
transform 1 0 1384 0 1 370
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1712256841
transform 1 0 1352 0 1 370
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1712256841
transform 1 0 1344 0 1 370
box -8 -3 16 105
use FILL  FILL_4715
timestamp 1712256841
transform 1 0 1336 0 1 370
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1712256841
transform 1 0 1288 0 1 370
box -8 -3 16 105
use FILL  FILL_4717
timestamp 1712256841
transform 1 0 1280 0 1 370
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1712256841
transform 1 0 1272 0 1 370
box -8 -3 16 105
use FILL  FILL_4719
timestamp 1712256841
transform 1 0 1264 0 1 370
box -8 -3 16 105
use FILL  FILL_4720
timestamp 1712256841
transform 1 0 1240 0 1 370
box -8 -3 16 105
use FILL  FILL_4721
timestamp 1712256841
transform 1 0 1232 0 1 370
box -8 -3 16 105
use FILL  FILL_4722
timestamp 1712256841
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_4723
timestamp 1712256841
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_4724
timestamp 1712256841
transform 1 0 1160 0 1 370
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1712256841
transform 1 0 1152 0 1 370
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1712256841
transform 1 0 1144 0 1 370
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1712256841
transform 1 0 1136 0 1 370
box -8 -3 16 105
use FILL  FILL_4728
timestamp 1712256841
transform 1 0 1104 0 1 370
box -8 -3 16 105
use FILL  FILL_4729
timestamp 1712256841
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1712256841
transform 1 0 1064 0 1 370
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1712256841
transform 1 0 1056 0 1 370
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1712256841
transform 1 0 1024 0 1 370
box -8 -3 16 105
use FILL  FILL_4733
timestamp 1712256841
transform 1 0 1016 0 1 370
box -8 -3 16 105
use FILL  FILL_4734
timestamp 1712256841
transform 1 0 1008 0 1 370
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1712256841
transform 1 0 1000 0 1 370
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1712256841
transform 1 0 952 0 1 370
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1712256841
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_4738
timestamp 1712256841
transform 1 0 936 0 1 370
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1712256841
transform 1 0 928 0 1 370
box -8 -3 16 105
use FILL  FILL_4740
timestamp 1712256841
transform 1 0 920 0 1 370
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1712256841
transform 1 0 856 0 1 370
box -8 -3 16 105
use FILL  FILL_4742
timestamp 1712256841
transform 1 0 848 0 1 370
box -8 -3 16 105
use FILL  FILL_4743
timestamp 1712256841
transform 1 0 840 0 1 370
box -8 -3 16 105
use FILL  FILL_4744
timestamp 1712256841
transform 1 0 832 0 1 370
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1712256841
transform 1 0 824 0 1 370
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1712256841
transform 1 0 816 0 1 370
box -8 -3 16 105
use FILL  FILL_4747
timestamp 1712256841
transform 1 0 808 0 1 370
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1712256841
transform 1 0 760 0 1 370
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1712256841
transform 1 0 752 0 1 370
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1712256841
transform 1 0 744 0 1 370
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1712256841
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_4752
timestamp 1712256841
transform 1 0 688 0 1 370
box -8 -3 16 105
use FILL  FILL_4753
timestamp 1712256841
transform 1 0 680 0 1 370
box -8 -3 16 105
use FILL  FILL_4754
timestamp 1712256841
transform 1 0 672 0 1 370
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1712256841
transform 1 0 664 0 1 370
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1712256841
transform 1 0 656 0 1 370
box -8 -3 16 105
use FILL  FILL_4757
timestamp 1712256841
transform 1 0 608 0 1 370
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1712256841
transform 1 0 600 0 1 370
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1712256841
transform 1 0 592 0 1 370
box -8 -3 16 105
use FILL  FILL_4760
timestamp 1712256841
transform 1 0 584 0 1 370
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1712256841
transform 1 0 552 0 1 370
box -8 -3 16 105
use FILL  FILL_4762
timestamp 1712256841
transform 1 0 544 0 1 370
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1712256841
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_4764
timestamp 1712256841
transform 1 0 496 0 1 370
box -8 -3 16 105
use FILL  FILL_4765
timestamp 1712256841
transform 1 0 488 0 1 370
box -8 -3 16 105
use FILL  FILL_4766
timestamp 1712256841
transform 1 0 480 0 1 370
box -8 -3 16 105
use FILL  FILL_4767
timestamp 1712256841
transform 1 0 472 0 1 370
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1712256841
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1712256841
transform 1 0 416 0 1 370
box -8 -3 16 105
use FILL  FILL_4770
timestamp 1712256841
transform 1 0 408 0 1 370
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1712256841
transform 1 0 400 0 1 370
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1712256841
transform 1 0 392 0 1 370
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1712256841
transform 1 0 360 0 1 370
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1712256841
transform 1 0 352 0 1 370
box -8 -3 16 105
use FILL  FILL_4775
timestamp 1712256841
transform 1 0 344 0 1 370
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1712256841
transform 1 0 336 0 1 370
box -8 -3 16 105
use FILL  FILL_4777
timestamp 1712256841
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_4778
timestamp 1712256841
transform 1 0 288 0 1 370
box -8 -3 16 105
use FILL  FILL_4779
timestamp 1712256841
transform 1 0 280 0 1 370
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1712256841
transform 1 0 248 0 1 370
box -8 -3 16 105
use FILL  FILL_4781
timestamp 1712256841
transform 1 0 240 0 1 370
box -8 -3 16 105
use FILL  FILL_4782
timestamp 1712256841
transform 1 0 232 0 1 370
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1712256841
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_4784
timestamp 1712256841
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1712256841
transform 1 0 168 0 1 370
box -8 -3 16 105
use FILL  FILL_4786
timestamp 1712256841
transform 1 0 160 0 1 370
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1712256841
transform 1 0 152 0 1 370
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1712256841
transform 1 0 144 0 1 370
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1712256841
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_4790
timestamp 1712256841
transform 1 0 104 0 1 370
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1712256841
transform 1 0 96 0 1 370
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1712256841
transform 1 0 88 0 1 370
box -8 -3 16 105
use FILL  FILL_4793
timestamp 1712256841
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1712256841
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_4795
timestamp 1712256841
transform 1 0 3424 0 -1 370
box -8 -3 16 105
use FILL  FILL_4796
timestamp 1712256841
transform 1 0 3320 0 -1 370
box -8 -3 16 105
use FILL  FILL_4797
timestamp 1712256841
transform 1 0 3312 0 -1 370
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1712256841
transform 1 0 3208 0 -1 370
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1712256841
transform 1 0 3200 0 -1 370
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1712256841
transform 1 0 3192 0 -1 370
box -8 -3 16 105
use FILL  FILL_4801
timestamp 1712256841
transform 1 0 3184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4802
timestamp 1712256841
transform 1 0 3080 0 -1 370
box -8 -3 16 105
use FILL  FILL_4803
timestamp 1712256841
transform 1 0 3072 0 -1 370
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1712256841
transform 1 0 2968 0 -1 370
box -8 -3 16 105
use FILL  FILL_4805
timestamp 1712256841
transform 1 0 2960 0 -1 370
box -8 -3 16 105
use FILL  FILL_4806
timestamp 1712256841
transform 1 0 2952 0 -1 370
box -8 -3 16 105
use FILL  FILL_4807
timestamp 1712256841
transform 1 0 2944 0 -1 370
box -8 -3 16 105
use FILL  FILL_4808
timestamp 1712256841
transform 1 0 2840 0 -1 370
box -8 -3 16 105
use FILL  FILL_4809
timestamp 1712256841
transform 1 0 2832 0 -1 370
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1712256841
transform 1 0 2824 0 -1 370
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1712256841
transform 1 0 2816 0 -1 370
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1712256841
transform 1 0 2808 0 -1 370
box -8 -3 16 105
use FILL  FILL_4813
timestamp 1712256841
transform 1 0 2800 0 -1 370
box -8 -3 16 105
use FILL  FILL_4814
timestamp 1712256841
transform 1 0 2744 0 -1 370
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1712256841
transform 1 0 2736 0 -1 370
box -8 -3 16 105
use FILL  FILL_4816
timestamp 1712256841
transform 1 0 2728 0 -1 370
box -8 -3 16 105
use FILL  FILL_4817
timestamp 1712256841
transform 1 0 2720 0 -1 370
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1712256841
transform 1 0 2680 0 -1 370
box -8 -3 16 105
use FILL  FILL_4819
timestamp 1712256841
transform 1 0 2672 0 -1 370
box -8 -3 16 105
use FILL  FILL_4820
timestamp 1712256841
transform 1 0 2664 0 -1 370
box -8 -3 16 105
use FILL  FILL_4821
timestamp 1712256841
transform 1 0 2656 0 -1 370
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1712256841
transform 1 0 2616 0 -1 370
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1712256841
transform 1 0 2608 0 -1 370
box -8 -3 16 105
use FILL  FILL_4824
timestamp 1712256841
transform 1 0 2600 0 -1 370
box -8 -3 16 105
use FILL  FILL_4825
timestamp 1712256841
transform 1 0 2592 0 -1 370
box -8 -3 16 105
use FILL  FILL_4826
timestamp 1712256841
transform 1 0 2552 0 -1 370
box -8 -3 16 105
use FILL  FILL_4827
timestamp 1712256841
transform 1 0 2544 0 -1 370
box -8 -3 16 105
use FILL  FILL_4828
timestamp 1712256841
transform 1 0 2536 0 -1 370
box -8 -3 16 105
use FILL  FILL_4829
timestamp 1712256841
transform 1 0 2528 0 -1 370
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1712256841
transform 1 0 2520 0 -1 370
box -8 -3 16 105
use FILL  FILL_4831
timestamp 1712256841
transform 1 0 2472 0 -1 370
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1712256841
transform 1 0 2464 0 -1 370
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1712256841
transform 1 0 2456 0 -1 370
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1712256841
transform 1 0 2448 0 -1 370
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1712256841
transform 1 0 2440 0 -1 370
box -8 -3 16 105
use FILL  FILL_4836
timestamp 1712256841
transform 1 0 2432 0 -1 370
box -8 -3 16 105
use FILL  FILL_4837
timestamp 1712256841
transform 1 0 2376 0 -1 370
box -8 -3 16 105
use FILL  FILL_4838
timestamp 1712256841
transform 1 0 2368 0 -1 370
box -8 -3 16 105
use FILL  FILL_4839
timestamp 1712256841
transform 1 0 2360 0 -1 370
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1712256841
transform 1 0 2352 0 -1 370
box -8 -3 16 105
use FILL  FILL_4841
timestamp 1712256841
transform 1 0 2344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1712256841
transform 1 0 2336 0 -1 370
box -8 -3 16 105
use FILL  FILL_4843
timestamp 1712256841
transform 1 0 2328 0 -1 370
box -8 -3 16 105
use FILL  FILL_4844
timestamp 1712256841
transform 1 0 2264 0 -1 370
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1712256841
transform 1 0 2256 0 -1 370
box -8 -3 16 105
use FILL  FILL_4846
timestamp 1712256841
transform 1 0 2248 0 -1 370
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1712256841
transform 1 0 2240 0 -1 370
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1712256841
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use FILL  FILL_4849
timestamp 1712256841
transform 1 0 2224 0 -1 370
box -8 -3 16 105
use FILL  FILL_4850
timestamp 1712256841
transform 1 0 2192 0 -1 370
box -8 -3 16 105
use FILL  FILL_4851
timestamp 1712256841
transform 1 0 2184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4852
timestamp 1712256841
transform 1 0 2136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1712256841
transform 1 0 2128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4854
timestamp 1712256841
transform 1 0 2120 0 -1 370
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1712256841
transform 1 0 2112 0 -1 370
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1712256841
transform 1 0 2104 0 -1 370
box -8 -3 16 105
use FILL  FILL_4857
timestamp 1712256841
transform 1 0 2072 0 -1 370
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1712256841
transform 1 0 2064 0 -1 370
box -8 -3 16 105
use FILL  FILL_4859
timestamp 1712256841
transform 1 0 2024 0 -1 370
box -8 -3 16 105
use FILL  FILL_4860
timestamp 1712256841
transform 1 0 2016 0 -1 370
box -8 -3 16 105
use FILL  FILL_4861
timestamp 1712256841
transform 1 0 2008 0 -1 370
box -8 -3 16 105
use FILL  FILL_4862
timestamp 1712256841
transform 1 0 2000 0 -1 370
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1712256841
transform 1 0 1992 0 -1 370
box -8 -3 16 105
use FILL  FILL_4864
timestamp 1712256841
transform 1 0 1960 0 -1 370
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1712256841
transform 1 0 1952 0 -1 370
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1712256841
transform 1 0 1944 0 -1 370
box -8 -3 16 105
use FILL  FILL_4867
timestamp 1712256841
transform 1 0 1896 0 -1 370
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1712256841
transform 1 0 1888 0 -1 370
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1712256841
transform 1 0 1880 0 -1 370
box -8 -3 16 105
use FILL  FILL_4870
timestamp 1712256841
transform 1 0 1872 0 -1 370
box -8 -3 16 105
use FILL  FILL_4871
timestamp 1712256841
transform 1 0 1864 0 -1 370
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1712256841
transform 1 0 1824 0 -1 370
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1712256841
transform 1 0 1816 0 -1 370
box -8 -3 16 105
use FILL  FILL_4874
timestamp 1712256841
transform 1 0 1808 0 -1 370
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1712256841
transform 1 0 1776 0 -1 370
box -8 -3 16 105
use FILL  FILL_4876
timestamp 1712256841
transform 1 0 1768 0 -1 370
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1712256841
transform 1 0 1760 0 -1 370
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1712256841
transform 1 0 1712 0 -1 370
box -8 -3 16 105
use FILL  FILL_4879
timestamp 1712256841
transform 1 0 1704 0 -1 370
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1712256841
transform 1 0 1696 0 -1 370
box -8 -3 16 105
use FILL  FILL_4881
timestamp 1712256841
transform 1 0 1688 0 -1 370
box -8 -3 16 105
use FILL  FILL_4882
timestamp 1712256841
transform 1 0 1680 0 -1 370
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1712256841
transform 1 0 1648 0 -1 370
box -8 -3 16 105
use FILL  FILL_4884
timestamp 1712256841
transform 1 0 1640 0 -1 370
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1712256841
transform 1 0 1592 0 -1 370
box -8 -3 16 105
use FILL  FILL_4886
timestamp 1712256841
transform 1 0 1584 0 -1 370
box -8 -3 16 105
use FILL  FILL_4887
timestamp 1712256841
transform 1 0 1576 0 -1 370
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1712256841
transform 1 0 1568 0 -1 370
box -8 -3 16 105
use FILL  FILL_4889
timestamp 1712256841
transform 1 0 1560 0 -1 370
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1712256841
transform 1 0 1552 0 -1 370
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1712256841
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_4892
timestamp 1712256841
transform 1 0 1480 0 -1 370
box -8 -3 16 105
use FILL  FILL_4893
timestamp 1712256841
transform 1 0 1472 0 -1 370
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1712256841
transform 1 0 1464 0 -1 370
box -8 -3 16 105
use FILL  FILL_4895
timestamp 1712256841
transform 1 0 1456 0 -1 370
box -8 -3 16 105
use FILL  FILL_4896
timestamp 1712256841
transform 1 0 1448 0 -1 370
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1712256841
transform 1 0 1416 0 -1 370
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1712256841
transform 1 0 1392 0 -1 370
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1712256841
transform 1 0 1368 0 -1 370
box -8 -3 16 105
use FILL  FILL_4900
timestamp 1712256841
transform 1 0 1360 0 -1 370
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1712256841
transform 1 0 1352 0 -1 370
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1712256841
transform 1 0 1344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4903
timestamp 1712256841
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use FILL  FILL_4904
timestamp 1712256841
transform 1 0 1288 0 -1 370
box -8 -3 16 105
use FILL  FILL_4905
timestamp 1712256841
transform 1 0 1280 0 -1 370
box -8 -3 16 105
use FILL  FILL_4906
timestamp 1712256841
transform 1 0 1272 0 -1 370
box -8 -3 16 105
use FILL  FILL_4907
timestamp 1712256841
transform 1 0 1264 0 -1 370
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1712256841
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_4909
timestamp 1712256841
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4910
timestamp 1712256841
transform 1 0 1208 0 -1 370
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1712256841
transform 1 0 1168 0 -1 370
box -8 -3 16 105
use FILL  FILL_4912
timestamp 1712256841
transform 1 0 1160 0 -1 370
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1712256841
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use FILL  FILL_4914
timestamp 1712256841
transform 1 0 1144 0 -1 370
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1712256841
transform 1 0 1136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4916
timestamp 1712256841
transform 1 0 1088 0 -1 370
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1712256841
transform 1 0 1080 0 -1 370
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1712256841
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1712256841
transform 1 0 1032 0 -1 370
box -8 -3 16 105
use FILL  FILL_4920
timestamp 1712256841
transform 1 0 1024 0 -1 370
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1712256841
transform 1 0 1016 0 -1 370
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1712256841
transform 1 0 1008 0 -1 370
box -8 -3 16 105
use FILL  FILL_4923
timestamp 1712256841
transform 1 0 1000 0 -1 370
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1712256841
transform 1 0 952 0 -1 370
box -8 -3 16 105
use FILL  FILL_4925
timestamp 1712256841
transform 1 0 944 0 -1 370
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1712256841
transform 1 0 936 0 -1 370
box -8 -3 16 105
use FILL  FILL_4927
timestamp 1712256841
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_4928
timestamp 1712256841
transform 1 0 896 0 -1 370
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1712256841
transform 1 0 888 0 -1 370
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1712256841
transform 1 0 880 0 -1 370
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1712256841
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1712256841
transform 1 0 840 0 -1 370
box -8 -3 16 105
use FILL  FILL_4933
timestamp 1712256841
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_4934
timestamp 1712256841
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1712256841
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1712256841
transform 1 0 776 0 -1 370
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1712256841
transform 1 0 768 0 -1 370
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1712256841
transform 1 0 760 0 -1 370
box -8 -3 16 105
use FILL  FILL_4939
timestamp 1712256841
transform 1 0 696 0 -1 370
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1712256841
transform 1 0 688 0 -1 370
box -8 -3 16 105
use FILL  FILL_4941
timestamp 1712256841
transform 1 0 680 0 -1 370
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1712256841
transform 1 0 672 0 -1 370
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1712256841
transform 1 0 664 0 -1 370
box -8 -3 16 105
use FILL  FILL_4944
timestamp 1712256841
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1712256841
transform 1 0 648 0 -1 370
box -8 -3 16 105
use FILL  FILL_4946
timestamp 1712256841
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1712256841
transform 1 0 576 0 -1 370
box -8 -3 16 105
use FILL  FILL_4948
timestamp 1712256841
transform 1 0 568 0 -1 370
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1712256841
transform 1 0 560 0 -1 370
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1712256841
transform 1 0 552 0 -1 370
box -8 -3 16 105
use FILL  FILL_4951
timestamp 1712256841
transform 1 0 544 0 -1 370
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1712256841
transform 1 0 512 0 -1 370
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1712256841
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1712256841
transform 1 0 456 0 -1 370
box -8 -3 16 105
use FILL  FILL_4955
timestamp 1712256841
transform 1 0 448 0 -1 370
box -8 -3 16 105
use FILL  FILL_4956
timestamp 1712256841
transform 1 0 440 0 -1 370
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1712256841
transform 1 0 432 0 -1 370
box -8 -3 16 105
use FILL  FILL_4958
timestamp 1712256841
transform 1 0 384 0 -1 370
box -8 -3 16 105
use FILL  FILL_4959
timestamp 1712256841
transform 1 0 376 0 -1 370
box -8 -3 16 105
use FILL  FILL_4960
timestamp 1712256841
transform 1 0 368 0 -1 370
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1712256841
transform 1 0 320 0 -1 370
box -8 -3 16 105
use FILL  FILL_4962
timestamp 1712256841
transform 1 0 312 0 -1 370
box -8 -3 16 105
use FILL  FILL_4963
timestamp 1712256841
transform 1 0 304 0 -1 370
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1712256841
transform 1 0 296 0 -1 370
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1712256841
transform 1 0 288 0 -1 370
box -8 -3 16 105
use FILL  FILL_4966
timestamp 1712256841
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_4967
timestamp 1712256841
transform 1 0 216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1712256841
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1712256841
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1712256841
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_4971
timestamp 1712256841
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4972
timestamp 1712256841
transform 1 0 136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4973
timestamp 1712256841
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1712256841
transform 1 0 120 0 -1 370
box -8 -3 16 105
use FILL  FILL_4975
timestamp 1712256841
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1712256841
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1712256841
transform 1 0 3368 0 1 170
box -8 -3 16 105
use FILL  FILL_4978
timestamp 1712256841
transform 1 0 3360 0 1 170
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1712256841
transform 1 0 3352 0 1 170
box -8 -3 16 105
use FILL  FILL_4980
timestamp 1712256841
transform 1 0 3344 0 1 170
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1712256841
transform 1 0 3256 0 1 170
box -8 -3 16 105
use FILL  FILL_4982
timestamp 1712256841
transform 1 0 3248 0 1 170
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1712256841
transform 1 0 3240 0 1 170
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1712256841
transform 1 0 3232 0 1 170
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1712256841
transform 1 0 3224 0 1 170
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1712256841
transform 1 0 3168 0 1 170
box -8 -3 16 105
use FILL  FILL_4987
timestamp 1712256841
transform 1 0 3160 0 1 170
box -8 -3 16 105
use FILL  FILL_4988
timestamp 1712256841
transform 1 0 3152 0 1 170
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1712256841
transform 1 0 3088 0 1 170
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1712256841
transform 1 0 3080 0 1 170
box -8 -3 16 105
use FILL  FILL_4991
timestamp 1712256841
transform 1 0 3048 0 1 170
box -8 -3 16 105
use FILL  FILL_4992
timestamp 1712256841
transform 1 0 3040 0 1 170
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1712256841
transform 1 0 3032 0 1 170
box -8 -3 16 105
use FILL  FILL_4994
timestamp 1712256841
transform 1 0 2952 0 1 170
box -8 -3 16 105
use FILL  FILL_4995
timestamp 1712256841
transform 1 0 2944 0 1 170
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1712256841
transform 1 0 2936 0 1 170
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1712256841
transform 1 0 2928 0 1 170
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1712256841
transform 1 0 2888 0 1 170
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1712256841
transform 1 0 2880 0 1 170
box -8 -3 16 105
use FILL  FILL_5000
timestamp 1712256841
transform 1 0 2816 0 1 170
box -8 -3 16 105
use FILL  FILL_5001
timestamp 1712256841
transform 1 0 2808 0 1 170
box -8 -3 16 105
use FILL  FILL_5002
timestamp 1712256841
transform 1 0 2800 0 1 170
box -8 -3 16 105
use FILL  FILL_5003
timestamp 1712256841
transform 1 0 2776 0 1 170
box -8 -3 16 105
use FILL  FILL_5004
timestamp 1712256841
transform 1 0 2736 0 1 170
box -8 -3 16 105
use FILL  FILL_5005
timestamp 1712256841
transform 1 0 2728 0 1 170
box -8 -3 16 105
use FILL  FILL_5006
timestamp 1712256841
transform 1 0 2720 0 1 170
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1712256841
transform 1 0 2712 0 1 170
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1712256841
transform 1 0 2704 0 1 170
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1712256841
transform 1 0 2648 0 1 170
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1712256841
transform 1 0 2640 0 1 170
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1712256841
transform 1 0 2632 0 1 170
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1712256841
transform 1 0 2624 0 1 170
box -8 -3 16 105
use FILL  FILL_5013
timestamp 1712256841
transform 1 0 2584 0 1 170
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1712256841
transform 1 0 2576 0 1 170
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1712256841
transform 1 0 2568 0 1 170
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1712256841
transform 1 0 2560 0 1 170
box -8 -3 16 105
use FILL  FILL_5017
timestamp 1712256841
transform 1 0 2520 0 1 170
box -8 -3 16 105
use FILL  FILL_5018
timestamp 1712256841
transform 1 0 2512 0 1 170
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1712256841
transform 1 0 2504 0 1 170
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1712256841
transform 1 0 2480 0 1 170
box -8 -3 16 105
use FILL  FILL_5021
timestamp 1712256841
transform 1 0 2472 0 1 170
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1712256841
transform 1 0 2464 0 1 170
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1712256841
transform 1 0 2424 0 1 170
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1712256841
transform 1 0 2416 0 1 170
box -8 -3 16 105
use FILL  FILL_5025
timestamp 1712256841
transform 1 0 2408 0 1 170
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1712256841
transform 1 0 2400 0 1 170
box -8 -3 16 105
use FILL  FILL_5027
timestamp 1712256841
transform 1 0 2360 0 1 170
box -8 -3 16 105
use FILL  FILL_5028
timestamp 1712256841
transform 1 0 2352 0 1 170
box -8 -3 16 105
use FILL  FILL_5029
timestamp 1712256841
transform 1 0 2344 0 1 170
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1712256841
transform 1 0 2336 0 1 170
box -8 -3 16 105
use FILL  FILL_5031
timestamp 1712256841
transform 1 0 2328 0 1 170
box -8 -3 16 105
use FILL  FILL_5032
timestamp 1712256841
transform 1 0 2280 0 1 170
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1712256841
transform 1 0 2272 0 1 170
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1712256841
transform 1 0 2264 0 1 170
box -8 -3 16 105
use FILL  FILL_5035
timestamp 1712256841
transform 1 0 2256 0 1 170
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1712256841
transform 1 0 2248 0 1 170
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1712256841
transform 1 0 2200 0 1 170
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1712256841
transform 1 0 2192 0 1 170
box -8 -3 16 105
use FILL  FILL_5039
timestamp 1712256841
transform 1 0 2184 0 1 170
box -8 -3 16 105
use FILL  FILL_5040
timestamp 1712256841
transform 1 0 2176 0 1 170
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1712256841
transform 1 0 2168 0 1 170
box -8 -3 16 105
use FILL  FILL_5042
timestamp 1712256841
transform 1 0 2160 0 1 170
box -8 -3 16 105
use FILL  FILL_5043
timestamp 1712256841
transform 1 0 2112 0 1 170
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1712256841
transform 1 0 2104 0 1 170
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1712256841
transform 1 0 2096 0 1 170
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1712256841
transform 1 0 2088 0 1 170
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1712256841
transform 1 0 2056 0 1 170
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1712256841
transform 1 0 2048 0 1 170
box -8 -3 16 105
use FILL  FILL_5049
timestamp 1712256841
transform 1 0 2040 0 1 170
box -8 -3 16 105
use FILL  FILL_5050
timestamp 1712256841
transform 1 0 2032 0 1 170
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1712256841
transform 1 0 2008 0 1 170
box -8 -3 16 105
use FILL  FILL_5052
timestamp 1712256841
transform 1 0 2000 0 1 170
box -8 -3 16 105
use FILL  FILL_5053
timestamp 1712256841
transform 1 0 1952 0 1 170
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1712256841
transform 1 0 1944 0 1 170
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1712256841
transform 1 0 1936 0 1 170
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1712256841
transform 1 0 1928 0 1 170
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1712256841
transform 1 0 1920 0 1 170
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1712256841
transform 1 0 1912 0 1 170
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1712256841
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1712256841
transform 1 0 1840 0 1 170
box -8 -3 16 105
use FILL  FILL_5061
timestamp 1712256841
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_5062
timestamp 1712256841
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_5063
timestamp 1712256841
transform 1 0 1816 0 1 170
box -8 -3 16 105
use FILL  FILL_5064
timestamp 1712256841
transform 1 0 1808 0 1 170
box -8 -3 16 105
use FILL  FILL_5065
timestamp 1712256841
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1712256841
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1712256841
transform 1 0 1736 0 1 170
box -8 -3 16 105
use FILL  FILL_5068
timestamp 1712256841
transform 1 0 1728 0 1 170
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1712256841
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_5070
timestamp 1712256841
transform 1 0 1712 0 1 170
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1712256841
transform 1 0 1704 0 1 170
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1712256841
transform 1 0 1656 0 1 170
box -8 -3 16 105
use FILL  FILL_5073
timestamp 1712256841
transform 1 0 1648 0 1 170
box -8 -3 16 105
use FILL  FILL_5074
timestamp 1712256841
transform 1 0 1640 0 1 170
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1712256841
transform 1 0 1632 0 1 170
box -8 -3 16 105
use FILL  FILL_5076
timestamp 1712256841
transform 1 0 1584 0 1 170
box -8 -3 16 105
use FILL  FILL_5077
timestamp 1712256841
transform 1 0 1576 0 1 170
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1712256841
transform 1 0 1568 0 1 170
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1712256841
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1712256841
transform 1 0 1536 0 1 170
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1712256841
transform 1 0 1504 0 1 170
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1712256841
transform 1 0 1496 0 1 170
box -8 -3 16 105
use FILL  FILL_5083
timestamp 1712256841
transform 1 0 1488 0 1 170
box -8 -3 16 105
use FILL  FILL_5084
timestamp 1712256841
transform 1 0 1480 0 1 170
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1712256841
transform 1 0 1432 0 1 170
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1712256841
transform 1 0 1424 0 1 170
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1712256841
transform 1 0 1416 0 1 170
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1712256841
transform 1 0 1376 0 1 170
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1712256841
transform 1 0 1368 0 1 170
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1712256841
transform 1 0 1360 0 1 170
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1712256841
transform 1 0 1352 0 1 170
box -8 -3 16 105
use FILL  FILL_5092
timestamp 1712256841
transform 1 0 1304 0 1 170
box -8 -3 16 105
use FILL  FILL_5093
timestamp 1712256841
transform 1 0 1296 0 1 170
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1712256841
transform 1 0 1288 0 1 170
box -8 -3 16 105
use FILL  FILL_5095
timestamp 1712256841
transform 1 0 1280 0 1 170
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1712256841
transform 1 0 1232 0 1 170
box -8 -3 16 105
use FILL  FILL_5097
timestamp 1712256841
transform 1 0 1224 0 1 170
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1712256841
transform 1 0 1216 0 1 170
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1712256841
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_5100
timestamp 1712256841
transform 1 0 1176 0 1 170
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1712256841
transform 1 0 1168 0 1 170
box -8 -3 16 105
use FILL  FILL_5102
timestamp 1712256841
transform 1 0 1160 0 1 170
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1712256841
transform 1 0 1112 0 1 170
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1712256841
transform 1 0 1104 0 1 170
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1712256841
transform 1 0 1096 0 1 170
box -8 -3 16 105
use FILL  FILL_5106
timestamp 1712256841
transform 1 0 1064 0 1 170
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1712256841
transform 1 0 1056 0 1 170
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1712256841
transform 1 0 1024 0 1 170
box -8 -3 16 105
use FILL  FILL_5109
timestamp 1712256841
transform 1 0 1016 0 1 170
box -8 -3 16 105
use FILL  FILL_5110
timestamp 1712256841
transform 1 0 1008 0 1 170
box -8 -3 16 105
use FILL  FILL_5111
timestamp 1712256841
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_5112
timestamp 1712256841
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1712256841
transform 1 0 952 0 1 170
box -8 -3 16 105
use FILL  FILL_5114
timestamp 1712256841
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1712256841
transform 1 0 904 0 1 170
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1712256841
transform 1 0 872 0 1 170
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1712256841
transform 1 0 864 0 1 170
box -8 -3 16 105
use FILL  FILL_5118
timestamp 1712256841
transform 1 0 856 0 1 170
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1712256841
transform 1 0 848 0 1 170
box -8 -3 16 105
use FILL  FILL_5120
timestamp 1712256841
transform 1 0 816 0 1 170
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1712256841
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_5122
timestamp 1712256841
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_5123
timestamp 1712256841
transform 1 0 752 0 1 170
box -8 -3 16 105
use FILL  FILL_5124
timestamp 1712256841
transform 1 0 744 0 1 170
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1712256841
transform 1 0 736 0 1 170
box -8 -3 16 105
use FILL  FILL_5126
timestamp 1712256841
transform 1 0 728 0 1 170
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1712256841
transform 1 0 680 0 1 170
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1712256841
transform 1 0 672 0 1 170
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1712256841
transform 1 0 632 0 1 170
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1712256841
transform 1 0 624 0 1 170
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1712256841
transform 1 0 616 0 1 170
box -8 -3 16 105
use FILL  FILL_5132
timestamp 1712256841
transform 1 0 608 0 1 170
box -8 -3 16 105
use FILL  FILL_5133
timestamp 1712256841
transform 1 0 600 0 1 170
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1712256841
transform 1 0 552 0 1 170
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1712256841
transform 1 0 544 0 1 170
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1712256841
transform 1 0 536 0 1 170
box -8 -3 16 105
use FILL  FILL_5137
timestamp 1712256841
transform 1 0 504 0 1 170
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1712256841
transform 1 0 496 0 1 170
box -8 -3 16 105
use FILL  FILL_5139
timestamp 1712256841
transform 1 0 488 0 1 170
box -8 -3 16 105
use FILL  FILL_5140
timestamp 1712256841
transform 1 0 456 0 1 170
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1712256841
transform 1 0 448 0 1 170
box -8 -3 16 105
use FILL  FILL_5142
timestamp 1712256841
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_5143
timestamp 1712256841
transform 1 0 400 0 1 170
box -8 -3 16 105
use FILL  FILL_5144
timestamp 1712256841
transform 1 0 392 0 1 170
box -8 -3 16 105
use FILL  FILL_5145
timestamp 1712256841
transform 1 0 384 0 1 170
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1712256841
transform 1 0 344 0 1 170
box -8 -3 16 105
use FILL  FILL_5147
timestamp 1712256841
transform 1 0 336 0 1 170
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1712256841
transform 1 0 328 0 1 170
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1712256841
transform 1 0 320 0 1 170
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1712256841
transform 1 0 272 0 1 170
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1712256841
transform 1 0 264 0 1 170
box -8 -3 16 105
use FILL  FILL_5152
timestamp 1712256841
transform 1 0 256 0 1 170
box -8 -3 16 105
use FILL  FILL_5153
timestamp 1712256841
transform 1 0 248 0 1 170
box -8 -3 16 105
use FILL  FILL_5154
timestamp 1712256841
transform 1 0 208 0 1 170
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1712256841
transform 1 0 200 0 1 170
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1712256841
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1712256841
transform 1 0 184 0 1 170
box -8 -3 16 105
use FILL  FILL_5158
timestamp 1712256841
transform 1 0 176 0 1 170
box -8 -3 16 105
use FILL  FILL_5159
timestamp 1712256841
transform 1 0 128 0 1 170
box -8 -3 16 105
use FILL  FILL_5160
timestamp 1712256841
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_5161
timestamp 1712256841
transform 1 0 112 0 1 170
box -8 -3 16 105
use FILL  FILL_5162
timestamp 1712256841
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_5163
timestamp 1712256841
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1712256841
transform 1 0 3424 0 -1 170
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1712256841
transform 1 0 3400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5166
timestamp 1712256841
transform 1 0 3392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1712256841
transform 1 0 3384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1712256841
transform 1 0 3376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1712256841
transform 1 0 3312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5170
timestamp 1712256841
transform 1 0 3304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1712256841
transform 1 0 3296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5172
timestamp 1712256841
transform 1 0 3288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1712256841
transform 1 0 3280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5174
timestamp 1712256841
transform 1 0 3272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5175
timestamp 1712256841
transform 1 0 3264 0 -1 170
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1712256841
transform 1 0 3216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5177
timestamp 1712256841
transform 1 0 3208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1712256841
transform 1 0 3200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1712256841
transform 1 0 3160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1712256841
transform 1 0 3152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1712256841
transform 1 0 3144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5182
timestamp 1712256841
transform 1 0 3136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1712256841
transform 1 0 3128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5184
timestamp 1712256841
transform 1 0 3120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1712256841
transform 1 0 3112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1712256841
transform 1 0 3048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1712256841
transform 1 0 3040 0 -1 170
box -8 -3 16 105
use FILL  FILL_5188
timestamp 1712256841
transform 1 0 3032 0 -1 170
box -8 -3 16 105
use FILL  FILL_5189
timestamp 1712256841
transform 1 0 3024 0 -1 170
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1712256841
transform 1 0 3016 0 -1 170
box -8 -3 16 105
use FILL  FILL_5191
timestamp 1712256841
transform 1 0 2992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5192
timestamp 1712256841
transform 1 0 2928 0 -1 170
box -8 -3 16 105
use FILL  FILL_5193
timestamp 1712256841
transform 1 0 2920 0 -1 170
box -8 -3 16 105
use FILL  FILL_5194
timestamp 1712256841
transform 1 0 2912 0 -1 170
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1712256841
transform 1 0 2904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1712256841
transform 1 0 2896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1712256841
transform 1 0 2832 0 -1 170
box -8 -3 16 105
use FILL  FILL_5198
timestamp 1712256841
transform 1 0 2824 0 -1 170
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1712256841
transform 1 0 2816 0 -1 170
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1712256841
transform 1 0 2808 0 -1 170
box -8 -3 16 105
use FILL  FILL_5201
timestamp 1712256841
transform 1 0 2744 0 -1 170
box -8 -3 16 105
use FILL  FILL_5202
timestamp 1712256841
transform 1 0 2712 0 -1 170
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1712256841
transform 1 0 2704 0 -1 170
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1712256841
transform 1 0 2696 0 -1 170
box -8 -3 16 105
use FILL  FILL_5205
timestamp 1712256841
transform 1 0 2688 0 -1 170
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1712256841
transform 1 0 2680 0 -1 170
box -8 -3 16 105
use FILL  FILL_5207
timestamp 1712256841
transform 1 0 2672 0 -1 170
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1712256841
transform 1 0 2664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5209
timestamp 1712256841
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5210
timestamp 1712256841
transform 1 0 2632 0 -1 170
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1712256841
transform 1 0 2624 0 -1 170
box -8 -3 16 105
use FILL  FILL_5212
timestamp 1712256841
transform 1 0 2616 0 -1 170
box -8 -3 16 105
use FILL  FILL_5213
timestamp 1712256841
transform 1 0 2576 0 -1 170
box -8 -3 16 105
use FILL  FILL_5214
timestamp 1712256841
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1712256841
transform 1 0 2560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1712256841
transform 1 0 2552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1712256841
transform 1 0 2544 0 -1 170
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1712256841
transform 1 0 2536 0 -1 170
box -8 -3 16 105
use FILL  FILL_5219
timestamp 1712256841
transform 1 0 2528 0 -1 170
box -8 -3 16 105
use FILL  FILL_5220
timestamp 1712256841
transform 1 0 2520 0 -1 170
box -8 -3 16 105
use FILL  FILL_5221
timestamp 1712256841
transform 1 0 2512 0 -1 170
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1712256841
transform 1 0 2464 0 -1 170
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1712256841
transform 1 0 2456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5224
timestamp 1712256841
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1712256841
transform 1 0 2440 0 -1 170
box -8 -3 16 105
use FILL  FILL_5226
timestamp 1712256841
transform 1 0 2432 0 -1 170
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1712256841
transform 1 0 2384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5228
timestamp 1712256841
transform 1 0 2376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5229
timestamp 1712256841
transform 1 0 2368 0 -1 170
box -8 -3 16 105
use FILL  FILL_5230
timestamp 1712256841
transform 1 0 2360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5231
timestamp 1712256841
transform 1 0 2352 0 -1 170
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1712256841
transform 1 0 2304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1712256841
transform 1 0 2296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1712256841
transform 1 0 2288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1712256841
transform 1 0 2280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5236
timestamp 1712256841
transform 1 0 2240 0 -1 170
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1712256841
transform 1 0 2232 0 -1 170
box -8 -3 16 105
use FILL  FILL_5238
timestamp 1712256841
transform 1 0 2224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5239
timestamp 1712256841
transform 1 0 2216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1712256841
transform 1 0 2176 0 -1 170
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1712256841
transform 1 0 2168 0 -1 170
box -8 -3 16 105
use FILL  FILL_5242
timestamp 1712256841
transform 1 0 2160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5243
timestamp 1712256841
transform 1 0 2128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5244
timestamp 1712256841
transform 1 0 2120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1712256841
transform 1 0 2112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1712256841
transform 1 0 2080 0 -1 170
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1712256841
transform 1 0 2056 0 -1 170
box -8 -3 16 105
use FILL  FILL_5248
timestamp 1712256841
transform 1 0 2048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5249
timestamp 1712256841
transform 1 0 2040 0 -1 170
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1712256841
transform 1 0 2032 0 -1 170
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1712256841
transform 1 0 1992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5252
timestamp 1712256841
transform 1 0 1984 0 -1 170
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1712256841
transform 1 0 1976 0 -1 170
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1712256841
transform 1 0 1936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5255
timestamp 1712256841
transform 1 0 1928 0 -1 170
box -8 -3 16 105
use FILL  FILL_5256
timestamp 1712256841
transform 1 0 1920 0 -1 170
box -8 -3 16 105
use FILL  FILL_5257
timestamp 1712256841
transform 1 0 1912 0 -1 170
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1712256841
transform 1 0 1872 0 -1 170
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1712256841
transform 1 0 1864 0 -1 170
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1712256841
transform 1 0 1856 0 -1 170
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1712256841
transform 1 0 1824 0 -1 170
box -8 -3 16 105
use FILL  FILL_5262
timestamp 1712256841
transform 1 0 1816 0 -1 170
box -8 -3 16 105
use FILL  FILL_5263
timestamp 1712256841
transform 1 0 1808 0 -1 170
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1712256841
transform 1 0 1800 0 -1 170
box -8 -3 16 105
use FILL  FILL_5265
timestamp 1712256841
transform 1 0 1752 0 -1 170
box -8 -3 16 105
use FILL  FILL_5266
timestamp 1712256841
transform 1 0 1744 0 -1 170
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1712256841
transform 1 0 1736 0 -1 170
box -8 -3 16 105
use FILL  FILL_5268
timestamp 1712256841
transform 1 0 1696 0 -1 170
box -8 -3 16 105
use FILL  FILL_5269
timestamp 1712256841
transform 1 0 1688 0 -1 170
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1712256841
transform 1 0 1680 0 -1 170
box -8 -3 16 105
use FILL  FILL_5271
timestamp 1712256841
transform 1 0 1640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1712256841
transform 1 0 1632 0 -1 170
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1712256841
transform 1 0 1624 0 -1 170
box -8 -3 16 105
use FILL  FILL_5274
timestamp 1712256841
transform 1 0 1616 0 -1 170
box -8 -3 16 105
use FILL  FILL_5275
timestamp 1712256841
transform 1 0 1592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5276
timestamp 1712256841
transform 1 0 1560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1712256841
transform 1 0 1552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5278
timestamp 1712256841
transform 1 0 1544 0 -1 170
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1712256841
transform 1 0 1536 0 -1 170
box -8 -3 16 105
use FILL  FILL_5280
timestamp 1712256841
transform 1 0 1504 0 -1 170
box -8 -3 16 105
use FILL  FILL_5281
timestamp 1712256841
transform 1 0 1472 0 -1 170
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1712256841
transform 1 0 1464 0 -1 170
box -8 -3 16 105
use FILL  FILL_5283
timestamp 1712256841
transform 1 0 1456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5284
timestamp 1712256841
transform 1 0 1448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5285
timestamp 1712256841
transform 1 0 1440 0 -1 170
box -8 -3 16 105
use FILL  FILL_5286
timestamp 1712256841
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1712256841
transform 1 0 1384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1712256841
transform 1 0 1376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5289
timestamp 1712256841
transform 1 0 1368 0 -1 170
box -8 -3 16 105
use FILL  FILL_5290
timestamp 1712256841
transform 1 0 1328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1712256841
transform 1 0 1320 0 -1 170
box -8 -3 16 105
use FILL  FILL_5292
timestamp 1712256841
transform 1 0 1312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5293
timestamp 1712256841
transform 1 0 1288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5294
timestamp 1712256841
transform 1 0 1280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1712256841
transform 1 0 1272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1712256841
transform 1 0 1232 0 -1 170
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1712256841
transform 1 0 1224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1712256841
transform 1 0 1216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5299
timestamp 1712256841
transform 1 0 1208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5300
timestamp 1712256841
transform 1 0 1160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1712256841
transform 1 0 1152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5302
timestamp 1712256841
transform 1 0 1144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5303
timestamp 1712256841
transform 1 0 1136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5304
timestamp 1712256841
transform 1 0 1112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5305
timestamp 1712256841
transform 1 0 1072 0 -1 170
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1712256841
transform 1 0 1064 0 -1 170
box -8 -3 16 105
use FILL  FILL_5307
timestamp 1712256841
transform 1 0 1056 0 -1 170
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1712256841
transform 1 0 1048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5309
timestamp 1712256841
transform 1 0 1040 0 -1 170
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1712256841
transform 1 0 992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1712256841
transform 1 0 984 0 -1 170
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1712256841
transform 1 0 976 0 -1 170
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1712256841
transform 1 0 968 0 -1 170
box -8 -3 16 105
use FILL  FILL_5314
timestamp 1712256841
transform 1 0 960 0 -1 170
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1712256841
transform 1 0 912 0 -1 170
box -8 -3 16 105
use FILL  FILL_5316
timestamp 1712256841
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5317
timestamp 1712256841
transform 1 0 896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1712256841
transform 1 0 864 0 -1 170
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1712256841
transform 1 0 856 0 -1 170
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1712256841
transform 1 0 848 0 -1 170
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1712256841
transform 1 0 800 0 -1 170
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1712256841
transform 1 0 792 0 -1 170
box -8 -3 16 105
use FILL  FILL_5323
timestamp 1712256841
transform 1 0 784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5324
timestamp 1712256841
transform 1 0 776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1712256841
transform 1 0 768 0 -1 170
box -8 -3 16 105
use FILL  FILL_5326
timestamp 1712256841
transform 1 0 760 0 -1 170
box -8 -3 16 105
use FILL  FILL_5327
timestamp 1712256841
transform 1 0 712 0 -1 170
box -8 -3 16 105
use FILL  FILL_5328
timestamp 1712256841
transform 1 0 704 0 -1 170
box -8 -3 16 105
use FILL  FILL_5329
timestamp 1712256841
transform 1 0 696 0 -1 170
box -8 -3 16 105
use FILL  FILL_5330
timestamp 1712256841
transform 1 0 688 0 -1 170
box -8 -3 16 105
use FILL  FILL_5331
timestamp 1712256841
transform 1 0 648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5332
timestamp 1712256841
transform 1 0 640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5333
timestamp 1712256841
transform 1 0 632 0 -1 170
box -8 -3 16 105
use FILL  FILL_5334
timestamp 1712256841
transform 1 0 624 0 -1 170
box -8 -3 16 105
use FILL  FILL_5335
timestamp 1712256841
transform 1 0 600 0 -1 170
box -8 -3 16 105
use FILL  FILL_5336
timestamp 1712256841
transform 1 0 592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5337
timestamp 1712256841
transform 1 0 560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5338
timestamp 1712256841
transform 1 0 552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5339
timestamp 1712256841
transform 1 0 544 0 -1 170
box -8 -3 16 105
use FILL  FILL_5340
timestamp 1712256841
transform 1 0 536 0 -1 170
box -8 -3 16 105
use FILL  FILL_5341
timestamp 1712256841
transform 1 0 488 0 -1 170
box -8 -3 16 105
use FILL  FILL_5342
timestamp 1712256841
transform 1 0 480 0 -1 170
box -8 -3 16 105
use FILL  FILL_5343
timestamp 1712256841
transform 1 0 472 0 -1 170
box -8 -3 16 105
use FILL  FILL_5344
timestamp 1712256841
transform 1 0 464 0 -1 170
box -8 -3 16 105
use FILL  FILL_5345
timestamp 1712256841
transform 1 0 456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5346
timestamp 1712256841
transform 1 0 448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5347
timestamp 1712256841
transform 1 0 424 0 -1 170
box -8 -3 16 105
use FILL  FILL_5348
timestamp 1712256841
transform 1 0 392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5349
timestamp 1712256841
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5350
timestamp 1712256841
transform 1 0 376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5351
timestamp 1712256841
transform 1 0 368 0 -1 170
box -8 -3 16 105
use FILL  FILL_5352
timestamp 1712256841
transform 1 0 360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5353
timestamp 1712256841
transform 1 0 312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5354
timestamp 1712256841
transform 1 0 304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5355
timestamp 1712256841
transform 1 0 296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5356
timestamp 1712256841
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5357
timestamp 1712256841
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5358
timestamp 1712256841
transform 1 0 272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5359
timestamp 1712256841
transform 1 0 224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5360
timestamp 1712256841
transform 1 0 216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5361
timestamp 1712256841
transform 1 0 208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5362
timestamp 1712256841
transform 1 0 200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5363
timestamp 1712256841
transform 1 0 168 0 -1 170
box -8 -3 16 105
use FILL  FILL_5364
timestamp 1712256841
transform 1 0 160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5365
timestamp 1712256841
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5366
timestamp 1712256841
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5367
timestamp 1712256841
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5368
timestamp 1712256841
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5369
timestamp 1712256841
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5370
timestamp 1712256841
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5371
timestamp 1712256841
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5372
timestamp 1712256841
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_5373
timestamp 1712256841
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_5374
timestamp 1712256841
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_5375
timestamp 1712256841
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1712256841
transform 1 0 2896 0 1 770
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1712256841
transform 1 0 3112 0 1 770
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1712256841
transform 1 0 3232 0 -1 770
box -5 -3 84 105
use INVX2  INVX2_0
timestamp 1712256841
transform 1 0 3312 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1712256841
transform 1 0 3232 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1712256841
transform 1 0 3288 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1712256841
transform 1 0 2904 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1712256841
transform 1 0 1464 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1712256841
transform 1 0 2784 0 1 170
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1712256841
transform 1 0 2960 0 1 170
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1712256841
transform 1 0 3000 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1712256841
transform 1 0 3248 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1712256841
transform 1 0 3408 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1712256841
transform 1 0 1488 0 1 970
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1712256841
transform 1 0 2984 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1712256841
transform 1 0 3000 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1712256841
transform 1 0 1032 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1712256841
transform 1 0 1096 0 1 770
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1712256841
transform 1 0 2016 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1712256841
transform 1 0 2720 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1712256841
transform 1 0 1464 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1712256841
transform 1 0 792 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1712256841
transform 1 0 1784 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1712256841
transform 1 0 2776 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1712256841
transform 1 0 1464 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1712256841
transform 1 0 648 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1712256841
transform 1 0 1792 0 1 570
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1712256841
transform 1 0 2448 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1712256841
transform 1 0 2704 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1712256841
transform 1 0 1176 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1712256841
transform 1 0 1088 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1712256841
transform 1 0 1432 0 1 770
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1712256841
transform 1 0 1608 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1712256841
transform 1 0 2720 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1712256841
transform 1 0 1344 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1712256841
transform 1 0 2968 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1712256841
transform 1 0 760 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1712256841
transform 1 0 1520 0 1 570
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1712256841
transform 1 0 2352 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1712256841
transform 1 0 1232 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1712256841
transform 1 0 1560 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1712256841
transform 1 0 928 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1712256841
transform 1 0 1528 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1712256841
transform 1 0 2632 0 1 970
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1712256841
transform 1 0 3064 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1712256841
transform 1 0 1320 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1712256841
transform 1 0 1040 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1712256841
transform 1 0 992 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1712256841
transform 1 0 1864 0 1 970
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1712256841
transform 1 0 2768 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1712256841
transform 1 0 912 0 1 970
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1712256841
transform 1 0 1648 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1712256841
transform 1 0 2736 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1712256841
transform 1 0 2600 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1712256841
transform 1 0 1576 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1712256841
transform 1 0 1680 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1712256841
transform 1 0 2800 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1712256841
transform 1 0 2856 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1712256841
transform 1 0 2688 0 1 170
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1712256841
transform 1 0 2352 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1712256841
transform 1 0 2784 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1712256841
transform 1 0 2488 0 1 170
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1712256841
transform 1 0 872 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1712256841
transform 1 0 424 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1712256841
transform 1 0 1888 0 1 170
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1712256841
transform 1 0 2024 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1712256841
transform 1 0 2600 0 1 370
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1712256841
transform 1 0 656 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1712256841
transform 1 0 1424 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1712256841
transform 1 0 2952 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1712256841
transform 1 0 2616 0 1 370
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1712256841
transform 1 0 568 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1712256841
transform 1 0 2800 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1712256841
transform 1 0 2736 0 1 370
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1712256841
transform 1 0 1152 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1712256841
transform 1 0 368 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1712256841
transform 1 0 704 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1712256841
transform 1 0 2648 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1712256841
transform 1 0 2544 0 1 170
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1712256841
transform 1 0 920 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1712256841
transform 1 0 1568 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1712256841
transform 1 0 1240 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1712256841
transform 1 0 552 0 1 570
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1712256841
transform 1 0 544 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1712256841
transform 1 0 2024 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1712256841
transform 1 0 1552 0 1 170
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1712256841
transform 1 0 2016 0 1 170
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1712256841
transform 1 0 3080 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1712256841
transform 1 0 2528 0 1 170
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1712256841
transform 1 0 824 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1712256841
transform 1 0 320 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1712256841
transform 1 0 768 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1712256841
transform 1 0 504 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1712256841
transform 1 0 720 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1712256841
transform 1 0 824 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1712256841
transform 1 0 2640 0 1 770
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1712256841
transform 1 0 2984 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1712256841
transform 1 0 2536 0 1 370
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1712256841
transform 1 0 672 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1712256841
transform 1 0 248 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1712256841
transform 1 0 480 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1712256841
transform 1 0 488 0 1 570
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1712256841
transform 1 0 1248 0 1 370
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1712256841
transform 1 0 1296 0 1 370
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1712256841
transform 1 0 2912 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1712256841
transform 1 0 2696 0 1 970
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1712256841
transform 1 0 1848 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1712256841
transform 1 0 2640 0 1 370
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1712256841
transform 1 0 1504 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1712256841
transform 1 0 832 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1712256841
transform 1 0 808 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1712256841
transform 1 0 832 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1712256841
transform 1 0 536 0 1 570
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1712256841
transform 1 0 2536 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1712256841
transform 1 0 2416 0 1 370
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1712256841
transform 1 0 2536 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1712256841
transform 1 0 1536 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1712256841
transform 1 0 1048 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1712256841
transform 1 0 872 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1712256841
transform 1 0 480 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1712256841
transform 1 0 656 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1712256841
transform 1 0 416 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1712256841
transform 1 0 328 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1712256841
transform 1 0 448 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1712256841
transform 1 0 256 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1712256841
transform 1 0 264 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1712256841
transform 1 0 208 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1712256841
transform 1 0 176 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1712256841
transform 1 0 1056 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1712256841
transform 1 0 1192 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1712256841
transform 1 0 1256 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1712256841
transform 1 0 1312 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1712256841
transform 1 0 1464 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1712256841
transform 1 0 1488 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1712256841
transform 1 0 1704 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1712256841
transform 1 0 1864 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1712256841
transform 1 0 1760 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1712256841
transform 1 0 1976 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1712256841
transform 1 0 2072 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1712256841
transform 1 0 2240 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1712256841
transform 1 0 2008 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1712256841
transform 1 0 2416 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1712256841
transform 1 0 2648 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1712256841
transform 1 0 2696 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1712256841
transform 1 0 2544 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1712256841
transform 1 0 2872 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1712256841
transform 1 0 3104 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1712256841
transform 1 0 2688 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1712256841
transform 1 0 3144 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1712256841
transform 1 0 3024 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1712256841
transform 1 0 2976 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1712256841
transform 1 0 3192 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1712256841
transform 1 0 3240 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1712256841
transform 1 0 3160 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1712256841
transform 1 0 3272 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1712256841
transform 1 0 3312 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1712256841
transform 1 0 3288 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1712256841
transform 1 0 2912 0 1 570
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1712256841
transform 1 0 3048 0 1 570
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1712256841
transform 1 0 3112 0 1 570
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1712256841
transform 1 0 3200 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1712256841
transform 1 0 3320 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1712256841
transform 1 0 3184 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1712256841
transform 1 0 3360 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1712256841
transform 1 0 3160 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1712256841
transform 1 0 3280 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1712256841
transform 1 0 2056 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1712256841
transform 1 0 2328 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1712256841
transform 1 0 2016 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1712256841
transform 1 0 1992 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1712256841
transform 1 0 2056 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1712256841
transform 1 0 1944 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1712256841
transform 1 0 2136 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1712256841
transform 1 0 1896 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1712256841
transform 1 0 2272 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1712256841
transform 1 0 2184 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1712256841
transform 1 0 2312 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1712256841
transform 1 0 2256 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1712256841
transform 1 0 2408 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1712256841
transform 1 0 2408 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1712256841
transform 1 0 2440 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1712256841
transform 1 0 2552 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1712256841
transform 1 0 2456 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1712256841
transform 1 0 2632 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1712256841
transform 1 0 2360 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1712256841
transform 1 0 2112 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1712256841
transform 1 0 1552 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1712256841
transform 1 0 2624 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1712256841
transform 1 0 2464 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1712256841
transform 1 0 2440 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1712256841
transform 1 0 1232 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1712256841
transform 1 0 1632 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1712256841
transform 1 0 1008 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1712256841
transform 1 0 928 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1712256841
transform 1 0 1456 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1712256841
transform 1 0 872 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1712256841
transform 1 0 1664 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1712256841
transform 1 0 952 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1712256841
transform 1 0 2848 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1712256841
transform 1 0 1032 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1712256841
transform 1 0 1368 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1712256841
transform 1 0 1688 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1712256841
transform 1 0 672 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1712256841
transform 1 0 1336 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1712256841
transform 1 0 1264 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1712256841
transform 1 0 776 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1712256841
transform 1 0 680 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1712256841
transform 1 0 648 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1712256841
transform 1 0 1088 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1712256841
transform 1 0 672 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1712256841
transform 1 0 752 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1712256841
transform 1 0 536 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1712256841
transform 1 0 552 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1712256841
transform 1 0 480 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1712256841
transform 1 0 88 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1712256841
transform 1 0 528 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1712256841
transform 1 0 224 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1712256841
transform 1 0 560 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1712256841
transform 1 0 808 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1712256841
transform 1 0 304 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1712256841
transform 1 0 320 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1712256841
transform 1 0 760 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1712256841
transform 1 0 776 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1712256841
transform 1 0 624 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1712256841
transform 1 0 448 0 1 970
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1712256841
transform 1 0 96 0 1 970
box -9 -3 26 105
use INVX2  INVX2_223
timestamp 1712256841
transform 1 0 192 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1712256841
transform 1 0 376 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_225
timestamp 1712256841
transform 1 0 80 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_226
timestamp 1712256841
transform 1 0 672 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_227
timestamp 1712256841
transform 1 0 648 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_228
timestamp 1712256841
transform 1 0 128 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_229
timestamp 1712256841
transform 1 0 208 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_230
timestamp 1712256841
transform 1 0 632 0 1 970
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1712256841
transform 1 0 928 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_232
timestamp 1712256841
transform 1 0 1688 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1712256841
transform 1 0 928 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_234
timestamp 1712256841
transform 1 0 728 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_235
timestamp 1712256841
transform 1 0 648 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_236
timestamp 1712256841
transform 1 0 536 0 1 970
box -9 -3 26 105
use INVX2  INVX2_237
timestamp 1712256841
transform 1 0 440 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1712256841
transform 1 0 912 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_239
timestamp 1712256841
transform 1 0 2440 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1712256841
transform 1 0 584 0 1 170
box -9 -3 26 105
use INVX2  INVX2_241
timestamp 1712256841
transform 1 0 800 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_242
timestamp 1712256841
transform 1 0 968 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_243
timestamp 1712256841
transform 1 0 432 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_244
timestamp 1712256841
transform 1 0 608 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_245
timestamp 1712256841
transform 1 0 728 0 1 570
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1712256841
transform 1 0 1264 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_247
timestamp 1712256841
transform 1 0 1120 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_248
timestamp 1712256841
transform 1 0 1296 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_249
timestamp 1712256841
transform 1 0 1120 0 1 570
box -9 -3 26 105
use INVX2  INVX2_250
timestamp 1712256841
transform 1 0 1256 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_251
timestamp 1712256841
transform 1 0 1400 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_252
timestamp 1712256841
transform 1 0 1384 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_253
timestamp 1712256841
transform 1 0 1144 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_254
timestamp 1712256841
transform 1 0 1216 0 1 370
box -9 -3 26 105
use INVX2  INVX2_255
timestamp 1712256841
transform 1 0 1304 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_256
timestamp 1712256841
transform 1 0 1376 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_257
timestamp 1712256841
transform 1 0 1528 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_258
timestamp 1712256841
transform 1 0 1400 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_259
timestamp 1712256841
transform 1 0 1440 0 1 570
box -9 -3 26 105
use INVX2  INVX2_260
timestamp 1712256841
transform 1 0 1560 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_261
timestamp 1712256841
transform 1 0 1504 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_262
timestamp 1712256841
transform 1 0 1664 0 1 170
box -9 -3 26 105
use INVX2  INVX2_263
timestamp 1712256841
transform 1 0 1696 0 1 370
box -9 -3 26 105
use INVX2  INVX2_264
timestamp 1712256841
transform 1 0 1896 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_265
timestamp 1712256841
transform 1 0 1880 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_266
timestamp 1712256841
transform 1 0 1720 0 1 570
box -9 -3 26 105
use INVX2  INVX2_267
timestamp 1712256841
transform 1 0 1728 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_268
timestamp 1712256841
transform 1 0 2064 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_269
timestamp 1712256841
transform 1 0 2144 0 1 370
box -9 -3 26 105
use INVX2  INVX2_270
timestamp 1712256841
transform 1 0 2008 0 1 370
box -9 -3 26 105
use INVX2  INVX2_271
timestamp 1712256841
transform 1 0 1920 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_272
timestamp 1712256841
transform 1 0 1784 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_273
timestamp 1712256841
transform 1 0 2096 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_274
timestamp 1712256841
transform 1 0 1848 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_275
timestamp 1712256841
transform 1 0 1560 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_276
timestamp 1712256841
transform 1 0 1664 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_277
timestamp 1712256841
transform 1 0 2640 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_278
timestamp 1712256841
transform 1 0 2064 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_279
timestamp 1712256841
transform 1 0 1864 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_280
timestamp 1712256841
transform 1 0 2216 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_281
timestamp 1712256841
transform 1 0 1848 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_282
timestamp 1712256841
transform 1 0 1032 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_283
timestamp 1712256841
transform 1 0 2360 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_284
timestamp 1712256841
transform 1 0 2184 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_285
timestamp 1712256841
transform 1 0 2376 0 1 770
box -9 -3 26 105
use INVX2  INVX2_286
timestamp 1712256841
transform 1 0 1960 0 1 970
box -9 -3 26 105
use INVX2  INVX2_287
timestamp 1712256841
transform 1 0 2248 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_288
timestamp 1712256841
transform 1 0 2344 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_289
timestamp 1712256841
transform 1 0 2264 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_290
timestamp 1712256841
transform 1 0 2280 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_291
timestamp 1712256841
transform 1 0 2512 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_292
timestamp 1712256841
transform 1 0 2792 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_293
timestamp 1712256841
transform 1 0 2424 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_294
timestamp 1712256841
transform 1 0 3392 0 1 770
box -9 -3 26 105
use INVX2  INVX2_295
timestamp 1712256841
transform 1 0 3272 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_296
timestamp 1712256841
transform 1 0 3288 0 1 770
box -9 -3 26 105
use INVX2  INVX2_297
timestamp 1712256841
transform 1 0 3344 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_298
timestamp 1712256841
transform 1 0 3368 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_299
timestamp 1712256841
transform 1 0 3368 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_300
timestamp 1712256841
transform 1 0 3392 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_301
timestamp 1712256841
transform 1 0 3360 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_302
timestamp 1712256841
transform 1 0 3368 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_303
timestamp 1712256841
transform 1 0 2936 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_304
timestamp 1712256841
transform 1 0 3208 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_305
timestamp 1712256841
transform 1 0 2792 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_306
timestamp 1712256841
transform 1 0 2376 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_307
timestamp 1712256841
transform 1 0 3176 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_308
timestamp 1712256841
transform 1 0 1296 0 1 970
box -9 -3 26 105
use INVX2  INVX2_309
timestamp 1712256841
transform 1 0 3208 0 1 170
box -9 -3 26 105
use INVX2  INVX2_310
timestamp 1712256841
transform 1 0 2584 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_311
timestamp 1712256841
transform 1 0 1320 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_312
timestamp 1712256841
transform 1 0 2960 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_313
timestamp 1712256841
transform 1 0 2384 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_314
timestamp 1712256841
transform 1 0 2648 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_315
timestamp 1712256841
transform 1 0 2504 0 1 770
box -9 -3 26 105
use INVX2  INVX2_316
timestamp 1712256841
transform 1 0 2480 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_317
timestamp 1712256841
transform 1 0 2824 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_318
timestamp 1712256841
transform 1 0 1720 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_319
timestamp 1712256841
transform 1 0 2552 0 1 970
box -9 -3 26 105
use INVX2  INVX2_320
timestamp 1712256841
transform 1 0 2584 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_321
timestamp 1712256841
transform 1 0 3248 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_322
timestamp 1712256841
transform 1 0 376 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_323
timestamp 1712256841
transform 1 0 352 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_324
timestamp 1712256841
transform 1 0 480 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_325
timestamp 1712256841
transform 1 0 2272 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_326
timestamp 1712256841
transform 1 0 1600 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_327
timestamp 1712256841
transform 1 0 2696 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_328
timestamp 1712256841
transform 1 0 760 0 1 170
box -9 -3 26 105
use INVX2  INVX2_329
timestamp 1712256841
transform 1 0 3000 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_330
timestamp 1712256841
transform 1 0 3048 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_331
timestamp 1712256841
transform 1 0 2848 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_332
timestamp 1712256841
transform 1 0 2616 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_333
timestamp 1712256841
transform 1 0 2776 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_334
timestamp 1712256841
transform 1 0 2440 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_335
timestamp 1712256841
transform 1 0 2456 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_336
timestamp 1712256841
transform 1 0 2456 0 1 770
box -9 -3 26 105
use INVX2  INVX2_337
timestamp 1712256841
transform 1 0 2584 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_338
timestamp 1712256841
transform 1 0 3280 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_339
timestamp 1712256841
transform 1 0 3224 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_340
timestamp 1712256841
transform 1 0 3264 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_341
timestamp 1712256841
transform 1 0 2984 0 1 970
box -9 -3 26 105
use INVX2  INVX2_342
timestamp 1712256841
transform 1 0 1248 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_343
timestamp 1712256841
transform 1 0 2488 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_344
timestamp 1712256841
transform 1 0 2832 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_345
timestamp 1712256841
transform 1 0 2320 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_346
timestamp 1712256841
transform 1 0 2560 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_347
timestamp 1712256841
transform 1 0 2944 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_348
timestamp 1712256841
transform 1 0 1648 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_349
timestamp 1712256841
transform 1 0 2544 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_350
timestamp 1712256841
transform 1 0 3408 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_351
timestamp 1712256841
transform 1 0 3232 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_352
timestamp 1712256841
transform 1 0 3400 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_353
timestamp 1712256841
transform 1 0 3352 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_354
timestamp 1712256841
transform 1 0 3392 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_355
timestamp 1712256841
transform 1 0 3328 0 1 2170
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1712256841
transform 1 0 3268 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1712256841
transform 1 0 3108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1712256841
transform 1 0 3148 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1712256841
transform 1 0 2908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1712256841
transform 1 0 2924 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1712256841
transform 1 0 2844 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1712256841
transform 1 0 3132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1712256841
transform 1 0 2948 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1712256841
transform 1 0 2948 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1712256841
transform 1 0 2844 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1712256841
transform 1 0 2844 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1712256841
transform 1 0 2812 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1712256841
transform 1 0 3140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1712256841
transform 1 0 3004 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1712256841
transform 1 0 2924 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1712256841
transform 1 0 2836 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1712256841
transform 1 0 2820 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1712256841
transform 1 0 2780 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1712256841
transform 1 0 2764 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1712256841
transform 1 0 3092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1712256841
transform 1 0 2988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1712256841
transform 1 0 2812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1712256841
transform 1 0 2804 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1712256841
transform 1 0 2780 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1712256841
transform 1 0 2740 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1712256841
transform 1 0 2740 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1712256841
transform 1 0 2772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1712256841
transform 1 0 2716 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1712256841
transform 1 0 1492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1712256841
transform 1 0 1428 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1712256841
transform 1 0 2812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1712256841
transform 1 0 2732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1712256841
transform 1 0 1532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1712256841
transform 1 0 1444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1712256841
transform 1 0 1404 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1712256841
transform 1 0 3212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1712256841
transform 1 0 2860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1712256841
transform 1 0 2716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1712256841
transform 1 0 2572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1712256841
transform 1 0 2572 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1712256841
transform 1 0 2516 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1712256841
transform 1 0 2508 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1712256841
transform 1 0 2372 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1712256841
transform 1 0 1988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1712256841
transform 1 0 1980 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1712256841
transform 1 0 1340 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1712256841
transform 1 0 1316 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1712256841
transform 1 0 1260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1712256841
transform 1 0 1076 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1712256841
transform 1 0 1012 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1712256841
transform 1 0 748 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1712256841
transform 1 0 716 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1712256841
transform 1 0 692 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1712256841
transform 1 0 676 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1712256841
transform 1 0 636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1712256841
transform 1 0 596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1712256841
transform 1 0 3228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1712256841
transform 1 0 2844 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1712256841
transform 1 0 2732 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1712256841
transform 1 0 2692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1712256841
transform 1 0 2668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1712256841
transform 1 0 3308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1712256841
transform 1 0 3244 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1712256841
transform 1 0 3228 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1712256841
transform 1 0 3180 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1712256841
transform 1 0 3100 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1712256841
transform 1 0 2972 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1712256841
transform 1 0 2940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1712256841
transform 1 0 2892 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1712256841
transform 1 0 2844 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1712256841
transform 1 0 3068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1712256841
transform 1 0 2988 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1712256841
transform 1 0 2964 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1712256841
transform 1 0 2852 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1712256841
transform 1 0 2940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1712256841
transform 1 0 2788 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1712256841
transform 1 0 2756 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1712256841
transform 1 0 3428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1712256841
transform 1 0 3308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1712256841
transform 1 0 3284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1712256841
transform 1 0 3284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1712256841
transform 1 0 3252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1712256841
transform 1 0 3236 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1712256841
transform 1 0 3428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1712256841
transform 1 0 3308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1712256841
transform 1 0 3292 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1712256841
transform 1 0 2796 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1712256841
transform 1 0 2692 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1712256841
transform 1 0 3004 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1712256841
transform 1 0 2932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1712256841
transform 1 0 3228 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1712256841
transform 1 0 3108 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1712256841
transform 1 0 2900 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1712256841
transform 1 0 2876 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1712256841
transform 1 0 2684 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1712256841
transform 1 0 2548 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1712256841
transform 1 0 2796 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1712256841
transform 1 0 2652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1712256841
transform 1 0 2556 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1712256841
transform 1 0 2420 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1712256841
transform 1 0 2140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1712256841
transform 1 0 2012 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1712256841
transform 1 0 2364 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1712256841
transform 1 0 2244 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1712256841
transform 1 0 2196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1712256841
transform 1 0 2076 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1712256841
transform 1 0 2028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1712256841
transform 1 0 1980 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1712256841
transform 1 0 1884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1712256841
transform 1 0 1868 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1712256841
transform 1 0 1612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1712256841
transform 1 0 1492 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1712256841
transform 1 0 1372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1712256841
transform 1 0 1316 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1712256841
transform 1 0 1396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1712256841
transform 1 0 1260 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1712256841
transform 1 0 1196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1712256841
transform 1 0 1196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1712256841
transform 1 0 1140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1712256841
transform 1 0 1060 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1712256841
transform 1 0 332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1712256841
transform 1 0 260 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1712256841
transform 1 0 388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1712256841
transform 1 0 332 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1712256841
transform 1 0 500 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1712256841
transform 1 0 420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1712256841
transform 1 0 636 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1712256841
transform 1 0 636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1712256841
transform 1 0 876 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1712256841
transform 1 0 852 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1712256841
transform 1 0 3420 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1712256841
transform 1 0 3252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1712256841
transform 1 0 3340 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1712256841
transform 1 0 3284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1712256841
transform 1 0 3420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1712256841
transform 1 0 3316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1712256841
transform 1 0 3420 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1712256841
transform 1 0 3388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1712256841
transform 1 0 3180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1712256841
transform 1 0 3140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1712256841
transform 1 0 3388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1712256841
transform 1 0 3372 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1712256841
transform 1 0 3332 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1712256841
transform 1 0 3300 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1712256841
transform 1 0 2996 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1712256841
transform 1 0 2796 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1712256841
transform 1 0 3428 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1712256841
transform 1 0 3404 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1712256841
transform 1 0 3388 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1712256841
transform 1 0 3388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1712256841
transform 1 0 3092 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1712256841
transform 1 0 2980 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1712256841
transform 1 0 2756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1712256841
transform 1 0 2692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1712256841
transform 1 0 2948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1712256841
transform 1 0 2820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1712256841
transform 1 0 3044 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1712256841
transform 1 0 2860 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1712256841
transform 1 0 2852 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1712256841
transform 1 0 2780 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1712256841
transform 1 0 2660 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1712256841
transform 1 0 2604 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1712256841
transform 1 0 2564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1712256841
transform 1 0 2492 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1712256841
transform 1 0 2468 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1712256841
transform 1 0 2404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1712256841
transform 1 0 2180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1712256841
transform 1 0 2180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1712256841
transform 1 0 2004 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1712256841
transform 1 0 1988 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1712256841
transform 1 0 2372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1712256841
transform 1 0 2348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1712256841
transform 1 0 2276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1712256841
transform 1 0 2276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1712256841
transform 1 0 2084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1712256841
transform 1 0 2084 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1712256841
transform 1 0 1892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1712256841
transform 1 0 1884 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1712256841
transform 1 0 1788 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1712256841
transform 1 0 1788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1712256841
transform 1 0 1692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1712256841
transform 1 0 1692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1712256841
transform 1 0 1604 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1712256841
transform 1 0 1580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1712256841
transform 1 0 1244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1712256841
transform 1 0 1196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1712256841
transform 1 0 860 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1712256841
transform 1 0 860 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1712256841
transform 1 0 220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1712256841
transform 1 0 156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1712256841
transform 1 0 180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1712256841
transform 1 0 84 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1712256841
transform 1 0 204 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1712256841
transform 1 0 204 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1712256841
transform 1 0 300 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1712256841
transform 1 0 284 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1712256841
transform 1 0 380 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1712256841
transform 1 0 364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1712256841
transform 1 0 428 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1712256841
transform 1 0 428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1712256841
transform 1 0 524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1712256841
transform 1 0 516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1712256841
transform 1 0 636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1712256841
transform 1 0 612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1712256841
transform 1 0 748 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1712256841
transform 1 0 708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1712256841
transform 1 0 972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1712256841
transform 1 0 796 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1712256841
transform 1 0 1284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1712256841
transform 1 0 1204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1712256841
transform 1 0 2772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1712256841
transform 1 0 2764 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1712256841
transform 1 0 2972 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1712256841
transform 1 0 2876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1712256841
transform 1 0 2980 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1712256841
transform 1 0 2932 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1712256841
transform 1 0 2852 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1712256841
transform 1 0 2852 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1712256841
transform 1 0 2636 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1712256841
transform 1 0 2636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1712256841
transform 1 0 2732 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1712256841
transform 1 0 2564 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1712256841
transform 1 0 2500 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1712256841
transform 1 0 2476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1712256841
transform 1 0 2348 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1712256841
transform 1 0 2268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1712256841
transform 1 0 2044 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1712256841
transform 1 0 2044 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1712256841
transform 1 0 2380 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1712256841
transform 1 0 2316 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1712256841
transform 1 0 2308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1712256841
transform 1 0 2196 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1712256841
transform 1 0 2148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1712256841
transform 1 0 2148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1712256841
transform 1 0 1948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1712256841
transform 1 0 1948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1712256841
transform 1 0 1844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1712256841
transform 1 0 1844 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1712256841
transform 1 0 1740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1712256841
transform 1 0 1724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1712256841
transform 1 0 1644 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1712256841
transform 1 0 1644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1712256841
transform 1 0 1596 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1712256841
transform 1 0 1532 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1712256841
transform 1 0 1436 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1712256841
transform 1 0 1428 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1712256841
transform 1 0 1308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1712256841
transform 1 0 1300 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1712256841
transform 1 0 1084 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1712256841
transform 1 0 1084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1712256841
transform 1 0 980 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1712256841
transform 1 0 924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1712256841
transform 1 0 220 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1712256841
transform 1 0 220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1712256841
transform 1 0 164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1712256841
transform 1 0 148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1712256841
transform 1 0 276 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1712256841
transform 1 0 276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1712256841
transform 1 0 388 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1712256841
transform 1 0 356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1712256841
transform 1 0 404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1712256841
transform 1 0 404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1712256841
transform 1 0 500 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1712256841
transform 1 0 492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1712256841
transform 1 0 548 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1712256841
transform 1 0 532 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1712256841
transform 1 0 652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1712256841
transform 1 0 644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1712256841
transform 1 0 756 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1712256841
transform 1 0 748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1712256841
transform 1 0 868 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1712256841
transform 1 0 860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1712256841
transform 1 0 1236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1712256841
transform 1 0 1212 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1712256841
transform 1 0 3324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1712256841
transform 1 0 3228 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1712256841
transform 1 0 3220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1712256841
transform 1 0 3204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1712256841
transform 1 0 3196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1712256841
transform 1 0 3164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1712256841
transform 1 0 3084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1712256841
transform 1 0 3268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1712256841
transform 1 0 3220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1712256841
transform 1 0 3204 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1712256841
transform 1 0 3204 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1712256841
transform 1 0 3204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1712256841
transform 1 0 3188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1712256841
transform 1 0 3172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1712256841
transform 1 0 3100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1712256841
transform 1 0 3092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1712256841
transform 1 0 3092 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1712256841
transform 1 0 3092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1712256841
transform 1 0 3052 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1712256841
transform 1 0 3052 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1712256841
transform 1 0 3020 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1712256841
transform 1 0 2972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1712256841
transform 1 0 2908 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1712256841
transform 1 0 2844 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1712256841
transform 1 0 2740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1712256841
transform 1 0 2908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1712256841
transform 1 0 2908 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1712256841
transform 1 0 2892 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1712256841
transform 1 0 2892 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1712256841
transform 1 0 2780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1712256841
transform 1 0 2780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1712256841
transform 1 0 3404 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1712256841
transform 1 0 3364 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1712256841
transform 1 0 3364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1712256841
transform 1 0 3292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1712256841
transform 1 0 3180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1712256841
transform 1 0 3276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1712256841
transform 1 0 3276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1712256841
transform 1 0 3180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1712256841
transform 1 0 3372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1712256841
transform 1 0 3356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1712256841
transform 1 0 3356 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1712256841
transform 1 0 3284 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1712256841
transform 1 0 3404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1712256841
transform 1 0 3364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1712256841
transform 1 0 3300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1712256841
transform 1 0 3292 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1712256841
transform 1 0 3428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1712256841
transform 1 0 3340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1712256841
transform 1 0 3260 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1712256841
transform 1 0 3244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1712256841
transform 1 0 3428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1712256841
transform 1 0 3364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1712256841
transform 1 0 3300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1712256841
transform 1 0 3316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1712256841
transform 1 0 3268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1712256841
transform 1 0 3244 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1712256841
transform 1 0 3204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1712256841
transform 1 0 3164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1712256841
transform 1 0 3060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1712256841
transform 1 0 3012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1712256841
transform 1 0 2980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1712256841
transform 1 0 2932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1712256841
transform 1 0 2892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1712256841
transform 1 0 2876 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1712256841
transform 1 0 2828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1712256841
transform 1 0 3348 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1712256841
transform 1 0 3292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1712256841
transform 1 0 3284 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1712256841
transform 1 0 3276 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1712256841
transform 1 0 3236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1712256841
transform 1 0 3220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1712256841
transform 1 0 3220 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1712256841
transform 1 0 3196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1712256841
transform 1 0 3060 0 1 2645
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1712256841
transform 1 0 3044 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1712256841
transform 1 0 3420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1712256841
transform 1 0 3276 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1712256841
transform 1 0 3260 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1712256841
transform 1 0 3228 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1712256841
transform 1 0 3156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1712256841
transform 1 0 3268 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1712256841
transform 1 0 3236 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1712256841
transform 1 0 3236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1712256841
transform 1 0 3180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1712256841
transform 1 0 3172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1712256841
transform 1 0 3172 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1712256841
transform 1 0 3132 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1712256841
transform 1 0 3164 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1712256841
transform 1 0 3068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1712256841
transform 1 0 2860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1712256841
transform 1 0 3228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1712256841
transform 1 0 3228 0 1 755
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1712256841
transform 1 0 3188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1712256841
transform 1 0 3116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1712256841
transform 1 0 3100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1712256841
transform 1 0 3356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1712256841
transform 1 0 3228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1712256841
transform 1 0 2708 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1712256841
transform 1 0 2612 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1712256841
transform 1 0 2356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1712256841
transform 1 0 1700 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1712256841
transform 1 0 1452 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1712256841
transform 1 0 1236 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1712256841
transform 1 0 3324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1712256841
transform 1 0 3316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1712256841
transform 1 0 3244 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1712256841
transform 1 0 3244 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1712256841
transform 1 0 3236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1712256841
transform 1 0 3172 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1712256841
transform 1 0 3044 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1712256841
transform 1 0 3044 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1712256841
transform 1 0 2908 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1712256841
transform 1 0 2908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1712256841
transform 1 0 3316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1712256841
transform 1 0 3300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1712256841
transform 1 0 3292 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1712256841
transform 1 0 3204 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1712256841
transform 1 0 3108 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1712256841
transform 1 0 3004 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1712256841
transform 1 0 3004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1712256841
transform 1 0 2980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1712256841
transform 1 0 2948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1712256841
transform 1 0 2764 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1712256841
transform 1 0 2668 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1712256841
transform 1 0 2660 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1712256841
transform 1 0 2652 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1712256841
transform 1 0 2628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1712256841
transform 1 0 2620 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1712256841
transform 1 0 2572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1712256841
transform 1 0 2540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1712256841
transform 1 0 2444 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1712256841
transform 1 0 2196 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1712256841
transform 1 0 1852 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1712256841
transform 1 0 1804 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1712256841
transform 1 0 1788 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1712256841
transform 1 0 1772 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1712256841
transform 1 0 1748 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1712256841
transform 1 0 1740 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1712256841
transform 1 0 1740 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1712256841
transform 1 0 1388 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1712256841
transform 1 0 1372 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1712256841
transform 1 0 1068 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1712256841
transform 1 0 1020 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1712256841
transform 1 0 844 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1712256841
transform 1 0 796 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1712256841
transform 1 0 796 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1712256841
transform 1 0 2596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1712256841
transform 1 0 2596 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1712256841
transform 1 0 2580 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1712256841
transform 1 0 2572 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1712256841
transform 1 0 2516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1712256841
transform 1 0 2396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1712256841
transform 1 0 2132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1712256841
transform 1 0 1556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1712256841
transform 1 0 1556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1712256841
transform 1 0 1532 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1712256841
transform 1 0 1492 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1712256841
transform 1 0 1452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1712256841
transform 1 0 1428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1712256841
transform 1 0 1428 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1712256841
transform 1 0 1420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1712256841
transform 1 0 1332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1712256841
transform 1 0 1284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1712256841
transform 1 0 1052 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1712256841
transform 1 0 980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1712256841
transform 1 0 980 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1712256841
transform 1 0 964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1712256841
transform 1 0 948 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1712256841
transform 1 0 1484 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1712256841
transform 1 0 1452 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1712256841
transform 1 0 1172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1712256841
transform 1 0 2876 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1712256841
transform 1 0 2780 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1712256841
transform 1 0 2756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1712256841
transform 1 0 3028 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1712256841
transform 1 0 2924 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1712256841
transform 1 0 2908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1712256841
transform 1 0 3092 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1712256841
transform 1 0 3060 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1712256841
transform 1 0 3316 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1712256841
transform 1 0 3316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1712256841
transform 1 0 3244 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1712256841
transform 1 0 3180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1712256841
transform 1 0 3428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1712256841
transform 1 0 3428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1712256841
transform 1 0 3372 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1712256841
transform 1 0 3332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1712256841
transform 1 0 2972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1712256841
transform 1 0 2948 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1712256841
transform 1 0 2924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1712256841
transform 1 0 2836 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1712256841
transform 1 0 2836 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1712256841
transform 1 0 2820 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1712256841
transform 1 0 2812 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1712256841
transform 1 0 2804 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1712256841
transform 1 0 2764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1712256841
transform 1 0 2756 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1712256841
transform 1 0 2756 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1712256841
transform 1 0 2748 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1712256841
transform 1 0 2748 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1712256841
transform 1 0 1476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1712256841
transform 1 0 1452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1712256841
transform 1 0 2524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1712256841
transform 1 0 2492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1712256841
transform 1 0 2492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1712256841
transform 1 0 2444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1712256841
transform 1 0 2332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1712256841
transform 1 0 2308 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1712256841
transform 1 0 2300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1712256841
transform 1 0 2260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1712256841
transform 1 0 2060 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1712256841
transform 1 0 1956 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1712256841
transform 1 0 1948 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1712256841
transform 1 0 1932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1712256841
transform 1 0 1836 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1712256841
transform 1 0 1836 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1712256841
transform 1 0 1700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1712256841
transform 1 0 1700 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1712256841
transform 1 0 1668 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1712256841
transform 1 0 1628 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1712256841
transform 1 0 1612 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1712256841
transform 1 0 2988 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1712256841
transform 1 0 2964 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1712256841
transform 1 0 2892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1712256841
transform 1 0 2884 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1712256841
transform 1 0 2860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1712256841
transform 1 0 3012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1712256841
transform 1 0 2916 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1712256841
transform 1 0 2860 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1712256841
transform 1 0 2836 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1712256841
transform 1 0 2796 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1712256841
transform 1 0 2772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1712256841
transform 1 0 1012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1712256841
transform 1 0 908 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1712256841
transform 1 0 1252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1712256841
transform 1 0 1076 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1712256841
transform 1 0 1028 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1712256841
transform 1 0 1028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1712256841
transform 1 0 916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1712256841
transform 1 0 2044 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1712256841
transform 1 0 2028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1712256841
transform 1 0 1924 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1712256841
transform 1 0 1740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1712256841
transform 1 0 1668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1712256841
transform 1 0 2700 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1712256841
transform 1 0 2676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1712256841
transform 1 0 1468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1712256841
transform 1 0 1428 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1712256841
transform 1 0 820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1712256841
transform 1 0 820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1712256841
transform 1 0 692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1712256841
transform 1 0 644 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1712256841
transform 1 0 1780 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1712256841
transform 1 0 1764 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1712256841
transform 1 0 1668 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1712256841
transform 1 0 1620 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1712256841
transform 1 0 3068 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1712256841
transform 1 0 2972 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1712256841
transform 1 0 2788 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1712256841
transform 1 0 2788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1712256841
transform 1 0 2572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1712256841
transform 1 0 2412 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1712256841
transform 1 0 2396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1712256841
transform 1 0 2364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1712256841
transform 1 0 1700 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1712256841
transform 1 0 1500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1712256841
transform 1 0 1500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1712256841
transform 1 0 1476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1712256841
transform 1 0 1460 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1712256841
transform 1 0 1452 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1712256841
transform 1 0 652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1712256841
transform 1 0 620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1712256841
transform 1 0 620 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1712256841
transform 1 0 1948 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1712256841
transform 1 0 1796 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1712256841
transform 1 0 1772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1712256841
transform 1 0 2652 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1712256841
transform 1 0 2620 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1712256841
transform 1 0 2436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1712256841
transform 1 0 2412 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1712256841
transform 1 0 2796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1712256841
transform 1 0 2748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1712256841
transform 1 0 1292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1712256841
transform 1 0 1188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1712256841
transform 1 0 1108 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1712256841
transform 1 0 1084 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1712256841
transform 1 0 956 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1712256841
transform 1 0 1404 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1712256841
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1712256841
transform 1 0 1092 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1712256841
transform 1 0 2620 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1712256841
transform 1 0 1628 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1712256841
transform 1 0 1628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1712256841
transform 1 0 2916 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1712256841
transform 1 0 2676 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1712256841
transform 1 0 1916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1712256841
transform 1 0 1484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1712256841
transform 1 0 1340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1712256841
transform 1 0 1268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1712256841
transform 1 0 1188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1712256841
transform 1 0 1124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1712256841
transform 1 0 2940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1712256841
transform 1 0 2908 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1712256841
transform 1 0 2876 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1712256841
transform 1 0 2764 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1712256841
transform 1 0 2756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1712256841
transform 1 0 756 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1712256841
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1712256841
transform 1 0 1604 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1712256841
transform 1 0 1532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1712256841
transform 1 0 1500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1712256841
transform 1 0 2332 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1712256841
transform 1 0 2332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1712256841
transform 1 0 2300 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1712256841
transform 1 0 1564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1712256841
transform 1 0 1540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1712256841
transform 1 0 916 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1712256841
transform 1 0 916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1712256841
transform 1 0 756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1712256841
transform 1 0 724 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1712256841
transform 1 0 1532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1712256841
transform 1 0 1492 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1712256841
transform 1 0 1308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1712256841
transform 1 0 1284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1712256841
transform 1 0 1284 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1712256841
transform 1 0 2772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1712256841
transform 1 0 2636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1712256841
transform 1 0 1684 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1712256841
transform 1 0 3084 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1712256841
transform 1 0 3084 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1712256841
transform 1 0 3068 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1712256841
transform 1 0 3068 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1712256841
transform 1 0 2916 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1712256841
transform 1 0 2292 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1712256841
transform 1 0 2132 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1712256841
transform 1 0 2108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1712256841
transform 1 0 1404 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1712256841
transform 1 0 1332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1712256841
transform 1 0 1300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1712256841
transform 1 0 1300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1712256841
transform 1 0 1276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1712256841
transform 1 0 1268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1712256841
transform 1 0 1116 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1712256841
transform 1 0 1092 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1712256841
transform 1 0 1052 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1712256841
transform 1 0 1004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1712256841
transform 1 0 1068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1712256841
transform 1 0 972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1712256841
transform 1 0 780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1712256841
transform 1 0 676 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1712256841
transform 1 0 676 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1712256841
transform 1 0 1972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1712256841
transform 1 0 1868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1712256841
transform 1 0 1868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1712256841
transform 1 0 1860 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1712256841
transform 1 0 1828 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1712256841
transform 1 0 2892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1712256841
transform 1 0 2836 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1712256841
transform 1 0 2780 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1712256841
transform 1 0 2780 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1712256841
transform 1 0 2652 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1712256841
transform 1 0 2548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1712256841
transform 1 0 2540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1712256841
transform 1 0 1060 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1712256841
transform 1 0 908 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1712256841
transform 1 0 684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1712256841
transform 1 0 1884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1712256841
transform 1 0 1684 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1712256841
transform 1 0 1636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1712256841
transform 1 0 1420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1712256841
transform 1 0 2740 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1712256841
transform 1 0 2716 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1712256841
transform 1 0 2660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1712256841
transform 1 0 2692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1712256841
transform 1 0 2636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1712256841
transform 1 0 1588 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1712256841
transform 1 0 1556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1712256841
transform 1 0 1556 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1712256841
transform 1 0 1500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1712256841
transform 1 0 1484 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1712256841
transform 1 0 3380 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1712256841
transform 1 0 3324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1712256841
transform 1 0 3244 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1712256841
transform 1 0 3228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1712256841
transform 1 0 3148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1712256841
transform 1 0 3076 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1712256841
transform 1 0 2900 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1712256841
transform 1 0 2900 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1712256841
transform 1 0 2748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1712256841
transform 1 0 2748 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1712256841
transform 1 0 2868 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1712256841
transform 1 0 2804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1712256841
transform 1 0 2796 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1712256841
transform 1 0 2780 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1712256841
transform 1 0 3020 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1712256841
transform 1 0 2820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1712256841
transform 1 0 2748 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1712256841
transform 1 0 2724 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1712256841
transform 1 0 2700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1712256841
transform 1 0 2692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1712256841
transform 1 0 2668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1712256841
transform 1 0 2628 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1712256841
transform 1 0 2604 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1712256841
transform 1 0 2604 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1712256841
transform 1 0 2364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1712256841
transform 1 0 2348 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1712256841
transform 1 0 3084 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1712256841
transform 1 0 2796 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1712256841
transform 1 0 2716 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1712256841
transform 1 0 2660 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1712256841
transform 1 0 2604 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1712256841
transform 1 0 2572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1712256841
transform 1 0 2524 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1712256841
transform 1 0 2524 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1712256841
transform 1 0 2500 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1712256841
transform 1 0 2500 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1712256841
transform 1 0 2468 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1712256841
transform 1 0 2468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1712256841
transform 1 0 1260 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1712256841
transform 1 0 1244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1712256841
transform 1 0 1148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1712256841
transform 1 0 1132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1712256841
transform 1 0 980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1712256841
transform 1 0 948 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1712256841
transform 1 0 892 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1712256841
transform 1 0 884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1712256841
transform 1 0 524 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1712256841
transform 1 0 508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1712256841
transform 1 0 1340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1712256841
transform 1 0 812 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1712256841
transform 1 0 580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1712256841
transform 1 0 444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1712256841
transform 1 0 308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1712256841
transform 1 0 300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1712256841
transform 1 0 148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1712256841
transform 1 0 84 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1712256841
transform 1 0 1900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1712256841
transform 1 0 1788 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1712256841
transform 1 0 1636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1712256841
transform 1 0 1636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1712256841
transform 1 0 1564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1712256841
transform 1 0 1388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1712256841
transform 1 0 2108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1712256841
transform 1 0 2092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1712256841
transform 1 0 2060 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1712256841
transform 1 0 2052 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1712256841
transform 1 0 2036 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1712256841
transform 1 0 2036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1712256841
transform 1 0 2012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1712256841
transform 1 0 1932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1712256841
transform 1 0 2556 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1712256841
transform 1 0 2556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1712256841
transform 1 0 2308 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1712256841
transform 1 0 1036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1712256841
transform 1 0 1036 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1712256841
transform 1 0 1380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1712256841
transform 1 0 1356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1712256841
transform 1 0 700 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1712256841
transform 1 0 692 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1712256841
transform 1 0 612 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1712256841
transform 1 0 1436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1712256841
transform 1 0 1372 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1712256841
transform 1 0 1036 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1712256841
transform 1 0 876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1712256841
transform 1 0 756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1712256841
transform 1 0 692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1712256841
transform 1 0 3116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1712256841
transform 1 0 3052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1712256841
transform 1 0 2924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1712256841
transform 1 0 2756 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1712256841
transform 1 0 2284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1712256841
transform 1 0 1996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1712256841
transform 1 0 1932 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1712256841
transform 1 0 2628 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1712256841
transform 1 0 2620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1712256841
transform 1 0 2316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1712256841
transform 1 0 1324 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1712256841
transform 1 0 1220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1712256841
transform 1 0 1196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1712256841
transform 1 0 1060 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1712256841
transform 1 0 1012 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1712256841
transform 1 0 972 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1712256841
transform 1 0 940 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1712256841
transform 1 0 868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1712256841
transform 1 0 604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1712256841
transform 1 0 492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1712256841
transform 1 0 3100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1712256841
transform 1 0 2788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1712256841
transform 1 0 2412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1712256841
transform 1 0 2356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1712256841
transform 1 0 2276 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1712256841
transform 1 0 2244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1712256841
transform 1 0 2740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1712256841
transform 1 0 2700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1712256841
transform 1 0 2532 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1712256841
transform 1 0 1156 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1712256841
transform 1 0 1116 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1712256841
transform 1 0 1268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1712256841
transform 1 0 1260 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1712256841
transform 1 0 1156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1712256841
transform 1 0 1148 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1712256841
transform 1 0 1132 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1712256841
transform 1 0 1604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1712256841
transform 1 0 932 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1712256841
transform 1 0 692 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1712256841
transform 1 0 660 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1712256841
transform 1 0 348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1712256841
transform 1 0 276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1712256841
transform 1 0 740 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1712256841
transform 1 0 724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1712256841
transform 1 0 652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1712256841
transform 1 0 580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1712256841
transform 1 0 148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1712256841
transform 1 0 148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1712256841
transform 1 0 2644 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1712256841
transform 1 0 2620 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1712256841
transform 1 0 2596 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1712256841
transform 1 0 2564 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1712256841
transform 1 0 2564 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1712256841
transform 1 0 2556 0 1 295
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1712256841
transform 1 0 2596 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1712256841
transform 1 0 2588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1712256841
transform 1 0 2580 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1712256841
transform 1 0 1140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1712256841
transform 1 0 1012 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1712256841
transform 1 0 1076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1712256841
transform 1 0 1028 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1712256841
transform 1 0 972 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1712256841
transform 1 0 916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1712256841
transform 1 0 916 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1712256841
transform 1 0 1652 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1712256841
transform 1 0 1604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1712256841
transform 1 0 1236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1712256841
transform 1 0 1220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1712256841
transform 1 0 132 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1712256841
transform 1 0 132 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1712256841
transform 1 0 612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1712256841
transform 1 0 452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1712256841
transform 1 0 420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1712256841
transform 1 0 364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1712256841
transform 1 0 364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1712256841
transform 1 0 516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1712256841
transform 1 0 516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1712256841
transform 1 0 484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1712256841
transform 1 0 404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1712256841
transform 1 0 380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1712256841
transform 1 0 2036 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1712256841
transform 1 0 2028 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1712256841
transform 1 0 1964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1712256841
transform 1 0 1940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1712256841
transform 1 0 1804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1712256841
transform 1 0 1588 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1712256841
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1712256841
transform 1 0 1548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1712256841
transform 1 0 1324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1712256841
transform 1 0 1284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1712256841
transform 1 0 1252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1712256841
transform 1 0 2004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1712256841
transform 1 0 2004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1712256841
transform 1 0 3068 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1712256841
transform 1 0 2980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1712256841
transform 1 0 2396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1712256841
transform 1 0 2172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1712256841
transform 1 0 2076 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1712256841
transform 1 0 1996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1712256841
transform 1 0 2620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1712256841
transform 1 0 2508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1712256841
transform 1 0 1412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1712256841
transform 1 0 1244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1712256841
transform 1 0 1244 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1712256841
transform 1 0 1564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1712256841
transform 1 0 1532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1712256841
transform 1 0 1164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1712256841
transform 1 0 844 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1712256841
transform 1 0 804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1712256841
transform 1 0 668 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1712256841
transform 1 0 708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1712256841
transform 1 0 676 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1712256841
transform 1 0 628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1712256841
transform 1 0 548 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1712256841
transform 1 0 452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1712256841
transform 1 0 340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1712256841
transform 1 0 220 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1712256841
transform 1 0 188 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1712256841
transform 1 0 988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1712256841
transform 1 0 820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1712256841
transform 1 0 748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1712256841
transform 1 0 748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1712256841
transform 1 0 732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1712256841
transform 1 0 492 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1712256841
transform 1 0 492 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1712256841
transform 1 0 428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1712256841
transform 1 0 412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1712256841
transform 1 0 380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1712256841
transform 1 0 732 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1712256841
transform 1 0 708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1712256841
transform 1 0 660 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1712256841
transform 1 0 460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1712256841
transform 1 0 356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1712256841
transform 1 0 348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1712256841
transform 1 0 836 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1712256841
transform 1 0 756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1712256841
transform 1 0 428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1712256841
transform 1 0 276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1712256841
transform 1 0 276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1712256841
transform 1 0 2620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1712256841
transform 1 0 2596 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1712256841
transform 1 0 2388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1712256841
transform 1 0 2268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1712256841
transform 1 0 2956 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1712256841
transform 1 0 2620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1712256841
transform 1 0 2572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1712256841
transform 1 0 2500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1712256841
transform 1 0 2388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1712256841
transform 1 0 2556 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1712256841
transform 1 0 2540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1712256841
transform 1 0 1596 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1712256841
transform 1 0 1100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1712256841
transform 1 0 1084 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1712256841
transform 1 0 1364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1712256841
transform 1 0 1332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1712256841
transform 1 0 684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1712256841
transform 1 0 628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1712256841
transform 1 0 508 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1712256841
transform 1 0 596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1712256841
transform 1 0 524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1712256841
transform 1 0 428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1712256841
transform 1 0 284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1712256841
transform 1 0 284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1712256841
transform 1 0 124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1712256841
transform 1 0 92 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1712256841
transform 1 0 484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1712256841
transform 1 0 460 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1712256841
transform 1 0 460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1712256841
transform 1 0 436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1712256841
transform 1 0 380 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1712256841
transform 1 0 1316 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1712256841
transform 1 0 524 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1712256841
transform 1 0 476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1712256841
transform 1 0 436 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1712256841
transform 1 0 404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1712256841
transform 1 0 1244 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1712256841
transform 1 0 996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1712256841
transform 1 0 988 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1712256841
transform 1 0 1340 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1712256841
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1712256841
transform 1 0 1268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1712256841
transform 1 0 1020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1712256841
transform 1 0 964 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1712256841
transform 1 0 2988 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1712256841
transform 1 0 2956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1712256841
transform 1 0 2772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1712256841
transform 1 0 2228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1712256841
transform 1 0 2212 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1712256841
transform 1 0 2188 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1712256841
transform 1 0 2044 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1712256841
transform 1 0 2012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1712256841
transform 1 0 2012 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1712256841
transform 1 0 1996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1712256841
transform 1 0 1884 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1712256841
transform 1 0 2652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1712256841
transform 1 0 2580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1712256841
transform 1 0 2508 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1712256841
transform 1 0 2444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1712256841
transform 1 0 2444 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1712256841
transform 1 0 1852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1712256841
transform 1 0 1844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1712256841
transform 1 0 1764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1712256841
transform 1 0 1724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1712256841
transform 1 0 1604 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1712256841
transform 1 0 2644 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1712256841
transform 1 0 2636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1712256841
transform 1 0 2516 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1712256841
transform 1 0 2500 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1712256841
transform 1 0 2484 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1712256841
transform 1 0 1332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1712256841
transform 1 0 1756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1712256841
transform 1 0 1484 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1712256841
transform 1 0 1308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1712256841
transform 1 0 1492 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1712256841
transform 1 0 1452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1712256841
transform 1 0 1044 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1712256841
transform 1 0 804 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1712256841
transform 1 0 788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1712256841
transform 1 0 820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1712256841
transform 1 0 628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1712256841
transform 1 0 580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1712256841
transform 1 0 548 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1712256841
transform 1 0 228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1712256841
transform 1 0 228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1712256841
transform 1 0 196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1712256841
transform 1 0 1972 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1712256841
transform 1 0 860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1712256841
transform 1 0 508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1712256841
transform 1 0 404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1712256841
transform 1 0 404 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1712256841
transform 1 0 548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1712256841
transform 1 0 548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1712256841
transform 1 0 508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1712256841
transform 1 0 460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1712256841
transform 1 0 364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1712256841
transform 1 0 356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1712256841
transform 1 0 2572 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1712256841
transform 1 0 2572 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1712256841
transform 1 0 2484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1712256841
transform 1 0 2364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1712256841
transform 1 0 2300 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1712256841
transform 1 0 2268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1712256841
transform 1 0 2260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1712256841
transform 1 0 2500 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1712256841
transform 1 0 2428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1712256841
transform 1 0 2420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1712256841
transform 1 0 1956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1712256841
transform 1 0 1948 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1712256841
transform 1 0 2652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1712256841
transform 1 0 2540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1712256841
transform 1 0 2484 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1712256841
transform 1 0 2476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1712256841
transform 1 0 2428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1712256841
transform 1 0 2404 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1712256841
transform 1 0 2868 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1712256841
transform 1 0 2188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1712256841
transform 1 0 1572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1712256841
transform 1 0 1484 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1712256841
transform 1 0 1468 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1712256841
transform 1 0 1084 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1712256841
transform 1 0 1060 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1712256841
transform 1 0 1028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1712256841
transform 1 0 884 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1712256841
transform 1 0 852 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1712256841
transform 1 0 852 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1712256841
transform 1 0 508 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1712256841
transform 1 0 508 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1712256841
transform 1 0 652 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1712256841
transform 1 0 644 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1712256841
transform 1 0 620 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1712256841
transform 1 0 468 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1712256841
transform 1 0 444 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1712256841
transform 1 0 404 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1712256841
transform 1 0 356 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1712256841
transform 1 0 476 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1712256841
transform 1 0 444 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1712256841
transform 1 0 308 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1712256841
transform 1 0 268 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1712256841
transform 1 0 292 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1712256841
transform 1 0 284 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1712256841
transform 1 0 196 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1712256841
transform 1 0 228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1712256841
transform 1 0 140 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1712256841
transform 1 0 188 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1712256841
transform 1 0 164 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1712256841
transform 1 0 1148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1712256841
transform 1 0 1068 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1712256841
transform 1 0 1068 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1712256841
transform 1 0 1204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1712256841
transform 1 0 1196 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1712256841
transform 1 0 1172 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1712256841
transform 1 0 1276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1712256841
transform 1 0 1260 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1712256841
transform 1 0 1236 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1712256841
transform 1 0 1404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1712256841
transform 1 0 1404 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1712256841
transform 1 0 1380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1712256841
transform 1 0 1356 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1712256841
transform 1 0 1476 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1712256841
transform 1 0 1452 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1712256841
transform 1 0 1444 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1712256841
transform 1 0 1540 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1712256841
transform 1 0 1524 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1712256841
transform 1 0 1516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1712256841
transform 1 0 1724 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1712256841
transform 1 0 1644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1712256841
transform 1 0 1900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1712256841
transform 1 0 1884 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1712256841
transform 1 0 1804 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1712256841
transform 1 0 1772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1712256841
transform 1 0 1772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1712256841
transform 1 0 2036 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1712256841
transform 1 0 2028 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1712256841
transform 1 0 2148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1712256841
transform 1 0 2068 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1712256841
transform 1 0 2052 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1712256841
transform 1 0 2236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1712256841
transform 1 0 2220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1712256841
transform 1 0 2220 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1712256841
transform 1 0 2036 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1712256841
transform 1 0 1972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1712256841
transform 1 0 1956 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1712256841
transform 1 0 2412 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1712256841
transform 1 0 2396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1712256841
transform 1 0 2380 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1712256841
transform 1 0 2380 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1712256841
transform 1 0 2740 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1712256841
transform 1 0 2660 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1712256841
transform 1 0 2612 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1712256841
transform 1 0 2708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1712256841
transform 1 0 2700 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1712256841
transform 1 0 2652 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1712256841
transform 1 0 2580 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1712256841
transform 1 0 2580 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1712256841
transform 1 0 2540 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1712256841
transform 1 0 2524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1712256841
transform 1 0 2876 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1712256841
transform 1 0 2836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1712256841
transform 1 0 2812 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1712256841
transform 1 0 3132 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1712256841
transform 1 0 3132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1712256841
transform 1 0 2980 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1712256841
transform 1 0 2732 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1712256841
transform 1 0 2700 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1712256841
transform 1 0 2700 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1712256841
transform 1 0 3156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1712256841
transform 1 0 3156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1712256841
transform 1 0 3116 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1712256841
transform 1 0 3116 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1712256841
transform 1 0 2996 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1712256841
transform 1 0 2860 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1712256841
transform 1 0 2972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1712256841
transform 1 0 2956 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1712256841
transform 1 0 2924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1712256841
transform 1 0 2908 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1712256841
transform 1 0 2892 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1712256841
transform 1 0 3252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1712256841
transform 1 0 3252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1712256841
transform 1 0 3188 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1712256841
transform 1 0 3188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1712256841
transform 1 0 3164 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1712256841
transform 1 0 3164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1712256841
transform 1 0 3396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1712256841
transform 1 0 3364 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1712256841
transform 1 0 3252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1712256841
transform 1 0 3196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1712256841
transform 1 0 3132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1712256841
transform 1 0 3084 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1712256841
transform 1 0 3084 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1712256841
transform 1 0 3020 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1712256841
transform 1 0 3260 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1712256841
transform 1 0 3228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1712256841
transform 1 0 3228 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1712256841
transform 1 0 3372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1712256841
transform 1 0 3292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1712256841
transform 1 0 3284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1712256841
transform 1 0 3260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1712256841
transform 1 0 3284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1712256841
transform 1 0 3188 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1712256841
transform 1 0 3372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1712256841
transform 1 0 3300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1712256841
transform 1 0 3292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1712256841
transform 1 0 3276 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1712256841
transform 1 0 3236 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1712256841
transform 1 0 2876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1712256841
transform 1 0 2844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1712256841
transform 1 0 3044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1712256841
transform 1 0 3028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1712256841
transform 1 0 3004 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1712256841
transform 1 0 2996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1712256841
transform 1 0 3132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1712256841
transform 1 0 3116 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1712256841
transform 1 0 3108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1712256841
transform 1 0 3108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1712256841
transform 1 0 3404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1712256841
transform 1 0 3404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1712256841
transform 1 0 3372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1712256841
transform 1 0 3356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1712256841
transform 1 0 3340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1712256841
transform 1 0 3212 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1712256841
transform 1 0 3204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1712256841
transform 1 0 3372 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1712256841
transform 1 0 3348 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1712256841
transform 1 0 3332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1712256841
transform 1 0 3244 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1712256841
transform 1 0 3260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1712256841
transform 1 0 3236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1712256841
transform 1 0 3212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1712256841
transform 1 0 3204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1712256841
transform 1 0 3196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1712256841
transform 1 0 3180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1712256841
transform 1 0 3140 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1712256841
transform 1 0 3052 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1712256841
transform 1 0 3364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1712256841
transform 1 0 3324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1712256841
transform 1 0 3148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1712256841
transform 1 0 3140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1712256841
transform 1 0 3076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1712256841
transform 1 0 2636 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1712256841
transform 1 0 1740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1712256841
transform 1 0 3356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1712256841
transform 1 0 3292 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1712256841
transform 1 0 3284 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1712256841
transform 1 0 3180 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1712256841
transform 1 0 3148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1712256841
transform 1 0 3060 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1712256841
transform 1 0 3028 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1712256841
transform 1 0 2100 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1712256841
transform 1 0 2084 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1712256841
transform 1 0 2020 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1712256841
transform 1 0 1932 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1712256841
transform 1 0 1932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1712256841
transform 1 0 1932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1712256841
transform 1 0 2100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1712256841
transform 1 0 1964 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1712256841
transform 1 0 1940 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1712256841
transform 1 0 1900 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1712256841
transform 1 0 1852 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1712256841
transform 1 0 1956 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1712256841
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1712256841
transform 1 0 2300 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1712256841
transform 1 0 2284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1712256841
transform 1 0 2308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1712256841
transform 1 0 2244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1712256841
transform 1 0 2204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1712256841
transform 1 0 2284 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1712256841
transform 1 0 2260 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1712256841
transform 1 0 2228 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1712256841
transform 1 0 2172 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1712256841
transform 1 0 2148 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1712256841
transform 1 0 2428 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1712256841
transform 1 0 2428 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1712256841
transform 1 0 2476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1712256841
transform 1 0 2460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1712256841
transform 1 0 2548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1712256841
transform 1 0 2420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1712256841
transform 1 0 2412 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1712256841
transform 1 0 2444 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1712256841
transform 1 0 2444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1712256841
transform 1 0 2412 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1712256841
transform 1 0 2380 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1712256841
transform 1 0 2292 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1712256841
transform 1 0 2652 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1712256841
transform 1 0 2628 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1712256841
transform 1 0 2124 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1712256841
transform 1 0 1996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1712256841
transform 1 0 1556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1712256841
transform 1 0 1532 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1712256841
transform 1 0 2596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1712256841
transform 1 0 2580 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1712256841
transform 1 0 2580 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1712256841
transform 1 0 1380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1712256841
transform 1 0 1268 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1712256841
transform 1 0 1268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1712256841
transform 1 0 1228 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1712256841
transform 1 0 1228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1712256841
transform 1 0 868 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1712256841
transform 1 0 1636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1712256841
transform 1 0 1604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1712256841
transform 1 0 1164 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1712256841
transform 1 0 1156 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1712256841
transform 1 0 1132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1712256841
transform 1 0 1020 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1712256841
transform 1 0 940 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1712256841
transform 1 0 940 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1712256841
transform 1 0 1452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1712256841
transform 1 0 1420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1712256841
transform 1 0 1156 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1712256841
transform 1 0 1116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1712256841
transform 1 0 1084 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1712256841
transform 1 0 1084 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1712256841
transform 1 0 1060 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1712256841
transform 1 0 1060 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1712256841
transform 1 0 1372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1712256841
transform 1 0 1364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1712256841
transform 1 0 1748 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1712256841
transform 1 0 1716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1712256841
transform 1 0 1276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1712256841
transform 1 0 1188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1712256841
transform 1 0 692 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1712256841
transform 1 0 628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1712256841
transform 1 0 484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1712256841
transform 1 0 1172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1712256841
transform 1 0 1116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1712256841
transform 1 0 836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1712256841
transform 1 0 772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1712256841
transform 1 0 748 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1712256841
transform 1 0 564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1712256841
transform 1 0 796 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1712256841
transform 1 0 500 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1712256841
transform 1 0 100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1712256841
transform 1 0 100 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1712256841
transform 1 0 284 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1712256841
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1712256841
transform 1 0 260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1712256841
transform 1 0 260 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1712256841
transform 1 0 316 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1712256841
transform 1 0 300 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1712256841
transform 1 0 316 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1712256841
transform 1 0 316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1712256841
transform 1 0 252 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1712256841
transform 1 0 204 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1712256841
transform 1 0 188 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1712256841
transform 1 0 756 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1712256841
transform 1 0 740 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1712256841
transform 1 0 652 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1712256841
transform 1 0 636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1712256841
transform 1 0 444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1712256841
transform 1 0 428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1712256841
transform 1 0 300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1712256841
transform 1 0 116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1712256841
transform 1 0 108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1712256841
transform 1 0 340 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1712256841
transform 1 0 260 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1712256841
transform 1 0 204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1712256841
transform 1 0 180 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1712256841
transform 1 0 420 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1712256841
transform 1 0 388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1712256841
transform 1 0 132 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1712256841
transform 1 0 132 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1712256841
transform 1 0 692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1712256841
transform 1 0 652 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1712256841
transform 1 0 132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1712256841
transform 1 0 68 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1712256841
transform 1 0 268 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1712256841
transform 1 0 220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1712256841
transform 1 0 220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1712256841
transform 1 0 220 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1712256841
transform 1 0 1772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1712256841
transform 1 0 1684 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1712256841
transform 1 0 1644 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1712256841
transform 1 0 916 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1712256841
transform 1 0 884 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1712256841
transform 1 0 748 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1712256841
transform 1 0 692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1712256841
transform 1 0 676 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1712256841
transform 1 0 668 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1712256841
transform 1 0 724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1712256841
transform 1 0 692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1712256841
transform 1 0 580 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1712256841
transform 1 0 580 0 1 1045
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1712256841
transform 1 0 508 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1712256841
transform 1 0 476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1712256841
transform 1 0 868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1712256841
transform 1 0 788 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1712256841
transform 1 0 740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1712256841
transform 1 0 1044 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1712256841
transform 1 0 492 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1712256841
transform 1 0 780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1712256841
transform 1 0 772 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1712256841
transform 1 0 764 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1712256841
transform 1 0 1212 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1712256841
transform 1 0 1164 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1712256841
transform 1 0 1388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1712256841
transform 1 0 1124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1712256841
transform 1 0 1060 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1712256841
transform 1 0 1500 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1712256841
transform 1 0 1420 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1712256841
transform 1 0 1708 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1712256841
transform 1 0 1580 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1712256841
transform 1 0 1340 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1712256841
transform 1 0 1116 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1712256841
transform 1 0 1548 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1712256841
transform 1 0 1212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1712256841
transform 1 0 1140 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1712256841
transform 1 0 1108 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1712256841
transform 1 0 1108 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1712256841
transform 1 0 1084 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1712256841
transform 1 0 988 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1712256841
transform 1 0 1636 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1712256841
transform 1 0 1228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1712256841
transform 1 0 1540 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1712256841
transform 1 0 1500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1712256841
transform 1 0 1444 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1712256841
transform 1 0 1404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1712256841
transform 1 0 1404 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1712256841
transform 1 0 1252 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1712256841
transform 1 0 1684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1712256841
transform 1 0 1604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1712256841
transform 1 0 1700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1712256841
transform 1 0 1684 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1712256841
transform 1 0 1732 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1712256841
transform 1 0 1708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1712256841
transform 1 0 1708 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1712256841
transform 1 0 1684 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1712256841
transform 1 0 1684 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1712256841
transform 1 0 1668 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1712256841
transform 1 0 1988 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1712256841
transform 1 0 1908 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1712256841
transform 1 0 1916 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1712256841
transform 1 0 1900 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1712256841
transform 1 0 2108 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1712256841
transform 1 0 2092 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1712256841
transform 1 0 2172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1712256841
transform 1 0 2156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1712256841
transform 1 0 2220 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1712256841
transform 1 0 2204 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1712256841
transform 1 0 2164 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1712256841
transform 1 0 1988 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1712256841
transform 1 0 1988 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1712256841
transform 1 0 1908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1712256841
transform 1 0 1892 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1712256841
transform 1 0 2148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1712256841
transform 1 0 2084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1712256841
transform 1 0 1604 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1712256841
transform 1 0 1580 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1712256841
transform 1 0 1548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1712256841
transform 1 0 1524 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1712256841
transform 1 0 1788 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1712256841
transform 1 0 1732 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1712256841
transform 1 0 1676 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1712256841
transform 1 0 1676 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1712256841
transform 1 0 2660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1712256841
transform 1 0 2660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1712256841
transform 1 0 1924 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1712256841
transform 1 0 1876 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1712256841
transform 1 0 1820 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1712256841
transform 1 0 1716 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1712256841
transform 1 0 1716 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1712256841
transform 1 0 2092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1712256841
transform 1 0 1860 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1712256841
transform 1 0 1756 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1712256841
transform 1 0 1756 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1712256841
transform 1 0 1012 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1712256841
transform 1 0 996 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1712256841
transform 1 0 2436 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1712256841
transform 1 0 2372 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1712256841
transform 1 0 2324 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1712256841
transform 1 0 2180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1712256841
transform 1 0 2172 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1712256841
transform 1 0 2036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1712256841
transform 1 0 1964 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1712256841
transform 1 0 1964 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1712256841
transform 1 0 2900 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1712256841
transform 1 0 2580 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1712256841
transform 1 0 2356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1712256841
transform 1 0 2260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1712256841
transform 1 0 2188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1712256841
transform 1 0 2084 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1712256841
transform 1 0 2812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1712256841
transform 1 0 2716 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1712256841
transform 1 0 2324 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1712256841
transform 1 0 2492 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1712256841
transform 1 0 2484 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1712256841
transform 1 0 2452 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1712256841
transform 1 0 2788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1712256841
transform 1 0 2788 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1712256841
transform 1 0 3404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1712256841
transform 1 0 3348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1712256841
transform 1 0 3292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1712256841
transform 1 0 3404 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1712256841
transform 1 0 3364 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1712256841
transform 1 0 3300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1712256841
transform 1 0 3300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1712256841
transform 1 0 3348 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1712256841
transform 1 0 3332 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1712256841
transform 1 0 3316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1712256841
transform 1 0 3276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1712256841
transform 1 0 3388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1712256841
transform 1 0 3388 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1712256841
transform 1 0 3412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1712256841
transform 1 0 3372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1712256841
transform 1 0 3364 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1712256841
transform 1 0 3404 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1712256841
transform 1 0 3380 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1712256841
transform 1 0 3348 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1712256841
transform 1 0 3308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1712256841
transform 1 0 2972 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1712256841
transform 1 0 2972 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1712256841
transform 1 0 2956 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1712256841
transform 1 0 2892 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1712256841
transform 1 0 2620 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1712256841
transform 1 0 2572 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1712256841
transform 1 0 3292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1712256841
transform 1 0 3260 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1712256841
transform 1 0 3220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1712256841
transform 1 0 3220 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1712256841
transform 1 0 3196 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1712256841
transform 1 0 3188 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1712256841
transform 1 0 3148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1712256841
transform 1 0 3140 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1712256841
transform 1 0 3036 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1712256841
transform 1 0 2780 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1712256841
transform 1 0 2740 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1712256841
transform 1 0 2356 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1712256841
transform 1 0 1492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1712256841
transform 1 0 1468 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1712256841
transform 1 0 884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1712256841
transform 1 0 3220 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1712256841
transform 1 0 3196 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1712256841
transform 1 0 3260 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1712256841
transform 1 0 3228 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1712256841
transform 1 0 3284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1712256841
transform 1 0 3236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1712256841
transform 1 0 3340 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1712256841
transform 1 0 3340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1712256841
transform 1 0 3332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1712256841
transform 1 0 2476 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1712256841
transform 1 0 2284 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1712256841
transform 1 0 2116 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1712256841
transform 1 0 2060 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1712256841
transform 1 0 1948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1712256841
transform 1 0 1804 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1712256841
transform 1 0 1676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1712256841
transform 1 0 1588 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1712256841
transform 1 0 1532 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1712256841
transform 1 0 1372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1712256841
transform 1 0 1316 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1712256841
transform 1 0 1292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1712256841
transform 1 0 1116 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1712256841
transform 1 0 3260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1712256841
transform 1 0 3236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1712256841
transform 1 0 3060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1712256841
transform 1 0 3036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1712256841
transform 1 0 1060 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1712256841
transform 1 0 940 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1712256841
transform 1 0 740 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1712256841
transform 1 0 532 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1712256841
transform 1 0 420 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1712256841
transform 1 0 372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1712256841
transform 1 0 356 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1712256841
transform 1 0 308 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1712256841
transform 1 0 252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1712256841
transform 1 0 172 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1712256841
transform 1 0 92 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1712256841
transform 1 0 92 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1712256841
transform 1 0 3348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1712256841
transform 1 0 3348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1712256841
transform 1 0 3340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1712256841
transform 1 0 3340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1712256841
transform 1 0 3268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1712256841
transform 1 0 3228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1712256841
transform 1 0 3132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1712256841
transform 1 0 3132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1712256841
transform 1 0 3100 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1712256841
transform 1 0 3052 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1712256841
transform 1 0 3004 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1712256841
transform 1 0 2988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1712256841
transform 1 0 2860 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1712256841
transform 1 0 2732 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1712256841
transform 1 0 2716 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1712256841
transform 1 0 2692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1712256841
transform 1 0 3348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1712256841
transform 1 0 3340 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1712256841
transform 1 0 3268 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1712256841
transform 1 0 3252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1712256841
transform 1 0 3156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1712256841
transform 1 0 2900 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1712256841
transform 1 0 2892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1712256841
transform 1 0 2772 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1712256841
transform 1 0 2692 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1712256841
transform 1 0 2652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1712256841
transform 1 0 2540 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1712256841
transform 1 0 2420 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1712256841
transform 1 0 2396 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1712256841
transform 1 0 2268 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1712256841
transform 1 0 2220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1712256841
transform 1 0 2204 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1712256841
transform 1 0 2116 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1712256841
transform 1 0 2068 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1712256841
transform 1 0 1964 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1712256841
transform 1 0 1860 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1712256841
transform 1 0 1756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1712256841
transform 1 0 1660 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1712256841
transform 1 0 1548 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1712256841
transform 1 0 1444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1712256841
transform 1 0 1332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1712256841
transform 1 0 1228 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1712256841
transform 1 0 1004 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1712256841
transform 1 0 900 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1712256841
transform 1 0 3052 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1712256841
transform 1 0 2948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1712256841
transform 1 0 2356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1712256841
transform 1 0 1116 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1712256841
transform 1 0 788 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1712256841
transform 1 0 676 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1712256841
transform 1 0 572 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1712256841
transform 1 0 436 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1712256841
transform 1 0 420 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1712256841
transform 1 0 308 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1712256841
transform 1 0 300 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1712256841
transform 1 0 196 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1712256841
transform 1 0 140 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1712256841
transform 1 0 84 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1712256841
transform 1 0 2964 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1712256841
transform 1 0 2868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1712256841
transform 1 0 2772 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1712256841
transform 1 0 2676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1712256841
transform 1 0 2580 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1712256841
transform 1 0 2484 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1712256841
transform 1 0 2388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1712256841
transform 1 0 2292 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1712256841
transform 1 0 2196 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1712256841
transform 1 0 2100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1712256841
transform 1 0 2004 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1712256841
transform 1 0 1996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1712256841
transform 1 0 1908 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1712256841
transform 1 0 1812 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1712256841
transform 1 0 1876 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1712256841
transform 1 0 1708 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1712256841
transform 1 0 1596 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1712256841
transform 1 0 1484 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1712256841
transform 1 0 1468 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1712256841
transform 1 0 1316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1712256841
transform 1 0 1100 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1712256841
transform 1 0 940 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1712256841
transform 1 0 780 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1712256841
transform 1 0 300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1712256841
transform 1 0 220 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1712256841
transform 1 0 140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1712256841
transform 1 0 100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1712256841
transform 1 0 92 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1712256841
transform 1 0 3348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1712256841
transform 1 0 3340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1712256841
transform 1 0 3236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1712256841
transform 1 0 3180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1712256841
transform 1 0 3124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1712256841
transform 1 0 2932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1712256841
transform 1 0 2812 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1712256841
transform 1 0 1972 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1712256841
transform 1 0 1204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1712256841
transform 1 0 892 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1712256841
transform 1 0 668 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1712256841
transform 1 0 556 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1712256841
transform 1 0 444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1712256841
transform 1 0 332 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1712256841
transform 1 0 2364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1712256841
transform 1 0 2340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1712256841
transform 1 0 2188 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1712256841
transform 1 0 2180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1712256841
transform 1 0 2172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1712256841
transform 1 0 1980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1712256841
transform 1 0 1924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1712256841
transform 1 0 1860 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1712256841
transform 1 0 2628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1712256841
transform 1 0 2556 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1712256841
transform 1 0 2532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1712256841
transform 1 0 2508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1712256841
transform 1 0 2476 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1712256841
transform 1 0 2452 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1712256841
transform 1 0 2644 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1712256841
transform 1 0 2388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1712256841
transform 1 0 2284 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1712256841
transform 1 0 2468 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1712256841
transform 1 0 2052 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1712256841
transform 1 0 1892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1712256841
transform 1 0 1748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1712256841
transform 1 0 1668 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1712256841
transform 1 0 1612 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1712256841
transform 1 0 1556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1712256841
transform 1 0 1412 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1712256841
transform 1 0 2780 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1712256841
transform 1 0 2524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1712256841
transform 1 0 1252 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1712256841
transform 1 0 1028 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1712256841
transform 1 0 868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1712256841
transform 1 0 236 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1712256841
transform 1 0 124 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1712256841
transform 1 0 92 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1712256841
transform 1 0 2812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1712256841
transform 1 0 2620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1712256841
transform 1 0 708 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1712256841
transform 1 0 564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1712256841
transform 1 0 460 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1712256841
transform 1 0 412 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1712256841
transform 1 0 324 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1712256841
transform 1 0 300 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1712256841
transform 1 0 2732 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1712256841
transform 1 0 2500 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1712256841
transform 1 0 1204 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1712256841
transform 1 0 804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1712256841
transform 1 0 2580 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1712256841
transform 1 0 2564 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1712256841
transform 1 0 2548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1712256841
transform 1 0 2524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1712256841
transform 1 0 2500 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1712256841
transform 1 0 2436 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1712256841
transform 1 0 2412 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1712256841
transform 1 0 2428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1712256841
transform 1 0 2324 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1712256841
transform 1 0 2188 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1712256841
transform 1 0 2020 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1712256841
transform 1 0 2884 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1712256841
transform 1 0 2804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1712256841
transform 1 0 2596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1712256841
transform 1 0 1228 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1712256841
transform 1 0 820 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1712256841
transform 1 0 732 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1712256841
transform 1 0 636 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1712256841
transform 1 0 572 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1712256841
transform 1 0 452 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1712256841
transform 1 0 388 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1712256841
transform 1 0 316 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1712256841
transform 1 0 252 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1712256841
transform 1 0 180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1712256841
transform 1 0 140 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1712256841
transform 1 0 3004 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1712256841
transform 1 0 2980 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1712256841
transform 1 0 3060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1712256841
transform 1 0 2996 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1712256841
transform 1 0 2940 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1712256841
transform 1 0 3012 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1712256841
transform 1 0 3012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1712256841
transform 1 0 2724 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1712256841
transform 1 0 2628 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1712256841
transform 1 0 2604 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1712256841
transform 1 0 1972 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1712256841
transform 1 0 1900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1712256841
transform 1 0 1740 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1712256841
transform 1 0 1540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1712256841
transform 1 0 1476 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1712256841
transform 1 0 1460 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1712256841
transform 1 0 1252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1712256841
transform 1 0 1188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1712256841
transform 1 0 1092 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1712256841
transform 1 0 324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1712256841
transform 1 0 212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1712256841
transform 1 0 180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1712256841
transform 1 0 164 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1712256841
transform 1 0 3076 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1712256841
transform 1 0 3012 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1712256841
transform 1 0 2956 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1712256841
transform 1 0 2492 0 1 3085
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1712256841
transform 1 0 2492 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1712256841
transform 1 0 2644 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1712256841
transform 1 0 2476 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1712256841
transform 1 0 2324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1712256841
transform 1 0 2252 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1712256841
transform 1 0 2108 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1712256841
transform 1 0 2044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1712256841
transform 1 0 1932 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1712256841
transform 1 0 1828 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1712256841
transform 1 0 1684 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1712256841
transform 1 0 1628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1712256841
transform 1 0 1476 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1712256841
transform 1 0 1364 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1712256841
transform 1 0 1340 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1712256841
transform 1 0 1268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1712256841
transform 1 0 1236 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1712256841
transform 1 0 1036 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1712256841
transform 1 0 1004 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1712256841
transform 1 0 916 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1712256841
transform 1 0 772 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1712256841
transform 1 0 756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1712256841
transform 1 0 660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1712256841
transform 1 0 644 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1712256841
transform 1 0 620 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1712256841
transform 1 0 580 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1712256841
transform 1 0 548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1712256841
transform 1 0 540 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1712256841
transform 1 0 2868 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1712256841
transform 1 0 2852 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1712256841
transform 1 0 2836 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1712256841
transform 1 0 3060 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1712256841
transform 1 0 2892 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1712256841
transform 1 0 2844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1712256841
transform 1 0 2828 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1712256841
transform 1 0 2724 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1712256841
transform 1 0 2516 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1712256841
transform 1 0 2372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1712256841
transform 1 0 2212 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1712256841
transform 1 0 2156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1712256841
transform 1 0 2044 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1712256841
transform 1 0 1980 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1712256841
transform 1 0 1892 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1712256841
transform 1 0 1740 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1712256841
transform 1 0 1620 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1712256841
transform 1 0 1540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1712256841
transform 1 0 1436 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1712256841
transform 1 0 1388 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1712256841
transform 1 0 1268 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1712256841
transform 1 0 1212 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1712256841
transform 1 0 1172 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1712256841
transform 1 0 2300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1712256841
transform 1 0 2276 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1712256841
transform 1 0 2220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1712256841
transform 1 0 2172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1712256841
transform 1 0 2148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1712256841
transform 1 0 2132 0 1 1445
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1712256841
transform 1 0 2132 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1712256841
transform 1 0 2124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1712256841
transform 1 0 2092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1712256841
transform 1 0 2084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1712256841
transform 1 0 1788 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1712256841
transform 1 0 1756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1712256841
transform 1 0 1756 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1712256841
transform 1 0 1692 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1712256841
transform 1 0 1684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1712256841
transform 1 0 1492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1712256841
transform 1 0 1100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1712256841
transform 1 0 764 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1712256841
transform 1 0 612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1712256841
transform 1 0 500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1712256841
transform 1 0 212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1712256841
transform 1 0 132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1712256841
transform 1 0 92 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1712256841
transform 1 0 92 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1712256841
transform 1 0 92 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1712256841
transform 1 0 92 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1712256841
transform 1 0 92 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1712256841
transform 1 0 92 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1712256841
transform 1 0 84 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1712256841
transform 1 0 2196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1712256841
transform 1 0 1716 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1712256841
transform 1 0 1652 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1712256841
transform 1 0 1388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1712256841
transform 1 0 548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1712256841
transform 1 0 380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1712256841
transform 1 0 356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1712256841
transform 1 0 308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1712256841
transform 1 0 268 0 1 585
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1712256841
transform 1 0 268 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1712256841
transform 1 0 244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1712256841
transform 1 0 244 0 1 585
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1712256841
transform 1 0 236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1712256841
transform 1 0 228 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1712256841
transform 1 0 228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1712256841
transform 1 0 204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1712256841
transform 1 0 180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1712256841
transform 1 0 2428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1712256841
transform 1 0 2420 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1712256841
transform 1 0 2348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1712256841
transform 1 0 2348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1712256841
transform 1 0 2284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1712256841
transform 1 0 2204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1712256841
transform 1 0 1924 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1712256841
transform 1 0 1860 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1712256841
transform 1 0 1796 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1712256841
transform 1 0 1748 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1712256841
transform 1 0 1508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1712256841
transform 1 0 1204 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1712256841
transform 1 0 956 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1712256841
transform 1 0 2148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1712256841
transform 1 0 2068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1712256841
transform 1 0 2012 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1712256841
transform 1 0 2012 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1712256841
transform 1 0 1924 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1712256841
transform 1 0 1308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1712256841
transform 1 0 612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1712256841
transform 1 0 532 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1712256841
transform 1 0 268 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1712256841
transform 1 0 172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1712256841
transform 1 0 140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1712256841
transform 1 0 124 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1712256841
transform 1 0 124 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1712256841
transform 1 0 124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1712256841
transform 1 0 124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1712256841
transform 1 0 123 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1712256841
transform 1 0 2324 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1712256841
transform 1 0 2252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1712256841
transform 1 0 2236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1712256841
transform 1 0 2188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1712256841
transform 1 0 2180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1712256841
transform 1 0 2180 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1712256841
transform 1 0 2180 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1712256841
transform 1 0 2108 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1712256841
transform 1 0 2084 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1712256841
transform 1 0 1844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1712256841
transform 1 0 1828 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1712256841
transform 1 0 1756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1712256841
transform 1 0 1652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1712256841
transform 1 0 1524 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1712256841
transform 1 0 1164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1712256841
transform 1 0 860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1712256841
transform 1 0 2692 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1712256841
transform 1 0 2660 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1712256841
transform 1 0 3068 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1712256841
transform 1 0 3004 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1712256841
transform 1 0 2972 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1712256841
transform 1 0 2884 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1712256841
transform 1 0 2588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1712256841
transform 1 0 2460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1712256841
transform 1 0 1780 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1712256841
transform 1 0 1372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1712256841
transform 1 0 1156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1712256841
transform 1 0 1140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1712256841
transform 1 0 2460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1712256841
transform 1 0 2436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1712256841
transform 1 0 2436 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1712256841
transform 1 0 2388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1712256841
transform 1 0 2380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1712256841
transform 1 0 2316 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1712256841
transform 1 0 2276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1712256841
transform 1 0 2084 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1712256841
transform 1 0 2020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1712256841
transform 1 0 1844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1712256841
transform 1 0 1700 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1712256841
transform 1 0 1484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1712256841
transform 1 0 1468 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1712256841
transform 1 0 1132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1712256841
transform 1 0 1044 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1712256841
transform 1 0 972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1712256841
transform 1 0 956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1712256841
transform 1 0 804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1712256841
transform 1 0 684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1712256841
transform 1 0 636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1712256841
transform 1 0 612 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1712256841
transform 1 0 612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1712256841
transform 1 0 596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1712256841
transform 1 0 596 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1712256841
transform 1 0 588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1712256841
transform 1 0 548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1712256841
transform 1 0 532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1712256841
transform 1 0 3140 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1712256841
transform 1 0 2796 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1712256841
transform 1 0 2780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1712256841
transform 1 0 3156 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1712256841
transform 1 0 3148 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1712256841
transform 1 0 3108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1712256841
transform 1 0 3012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1712256841
transform 1 0 2876 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1712256841
transform 1 0 2588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1712256841
transform 1 0 3188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1712256841
transform 1 0 3116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1712256841
transform 1 0 2876 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1712256841
transform 1 0 2844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1712256841
transform 1 0 2596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1712256841
transform 1 0 2380 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1712256841
transform 1 0 2364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1712256841
transform 1 0 2364 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1712256841
transform 1 0 2364 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1712256841
transform 1 0 2348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1712256841
transform 1 0 2340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1712256841
transform 1 0 2276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1712256841
transform 1 0 2252 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1712256841
transform 1 0 2244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1712256841
transform 1 0 2036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1712256841
transform 1 0 1812 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1712256841
transform 1 0 1668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1712256841
transform 1 0 1452 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1712256841
transform 1 0 1100 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1712256841
transform 1 0 924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1712256841
transform 1 0 772 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1712256841
transform 1 0 620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1712256841
transform 1 0 556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1712256841
transform 1 0 2780 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1712256841
transform 1 0 2708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1712256841
transform 1 0 2508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1712256841
transform 1 0 1964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1712256841
transform 1 0 1540 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1712256841
transform 1 0 1532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1712256841
transform 1 0 1244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1712256841
transform 1 0 1164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1712256841
transform 1 0 988 0 1 1885
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1712256841
transform 1 0 980 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1712256841
transform 1 0 916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1712256841
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1712256841
transform 1 0 548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1712256841
transform 1 0 548 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1712256841
transform 1 0 548 0 1 1455
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1712256841
transform 1 0 532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1712256841
transform 1 0 500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1712256841
transform 1 0 492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1712256841
transform 1 0 2684 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1712256841
transform 1 0 2612 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1712256841
transform 1 0 2444 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1712256841
transform 1 0 3132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1712256841
transform 1 0 3036 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1712256841
transform 1 0 2996 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1712256841
transform 1 0 2980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1712256841
transform 1 0 2444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1712256841
transform 1 0 2396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1712256841
transform 1 0 2372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1712256841
transform 1 0 2284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1712256841
transform 1 0 2268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1712256841
transform 1 0 2228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1712256841
transform 1 0 2164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1712256841
transform 1 0 1868 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1712256841
transform 1 0 1812 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1712256841
transform 1 0 1740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1712256841
transform 1 0 1444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1712256841
transform 1 0 1172 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1712256841
transform 1 0 900 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1712256841
transform 1 0 340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1712256841
transform 1 0 276 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1712256841
transform 1 0 236 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1712256841
transform 1 0 2492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1712256841
transform 1 0 2468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1712256841
transform 1 0 2172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1712256841
transform 1 0 1508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1712256841
transform 1 0 1492 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1712256841
transform 1 0 1212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1712256841
transform 1 0 1132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1712256841
transform 1 0 956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1712256841
transform 1 0 540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1712256841
transform 1 0 236 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1712256841
transform 1 0 212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1712256841
transform 1 0 204 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1712256841
transform 1 0 204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1712256841
transform 1 0 196 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1712256841
transform 1 0 148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1712256841
transform 1 0 148 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1712256841
transform 1 0 140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1712256841
transform 1 0 2844 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1712256841
transform 1 0 2820 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1712256841
transform 1 0 2620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1712256841
transform 1 0 1668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1712256841
transform 1 0 1580 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1712256841
transform 1 0 1340 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1712256841
transform 1 0 1324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1712256841
transform 1 0 2628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1712256841
transform 1 0 2628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1712256841
transform 1 0 2548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1712256841
transform 1 0 2548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1712256841
transform 1 0 2516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1712256841
transform 1 0 2492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1712256841
transform 1 0 2348 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1712256841
transform 1 0 2236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1712256841
transform 1 0 2156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1712256841
transform 1 0 1972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1712256841
transform 1 0 1932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1712256841
transform 1 0 1884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1712256841
transform 1 0 1772 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1712256841
transform 1 0 1476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1712256841
transform 1 0 1332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1712256841
transform 1 0 1132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1712256841
transform 1 0 996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1712256841
transform 1 0 924 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1712256841
transform 1 0 756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1712256841
transform 1 0 508 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1712256841
transform 1 0 508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1712256841
transform 1 0 492 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1712256841
transform 1 0 484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1712256841
transform 1 0 468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1712256841
transform 1 0 468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1712256841
transform 1 0 452 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1712256841
transform 1 0 452 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1712256841
transform 1 0 436 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1712256841
transform 1 0 428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1712256841
transform 1 0 428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1712256841
transform 1 0 380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1712256841
transform 1 0 3156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1712256841
transform 1 0 3068 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1712256841
transform 1 0 3012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1712256841
transform 1 0 2988 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1712256841
transform 1 0 3308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1712256841
transform 1 0 3292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1712256841
transform 1 0 3196 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1712256841
transform 1 0 2860 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1712256841
transform 1 0 3068 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1712256841
transform 1 0 2988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1712256841
transform 1 0 2924 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1712256841
transform 1 0 2900 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1712256841
transform 1 0 2780 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1712256841
transform 1 0 2564 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1712256841
transform 1 0 2388 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1712256841
transform 1 0 2356 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1712256841
transform 1 0 2324 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1712256841
transform 1 0 2316 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1712256841
transform 1 0 2300 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1712256841
transform 1 0 2228 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1712256841
transform 1 0 2076 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1712256841
transform 1 0 1956 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1712256841
transform 1 0 1852 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1712256841
transform 1 0 1796 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1712256841
transform 1 0 1772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1712256841
transform 1 0 1756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1712256841
transform 1 0 1612 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1712256841
transform 1 0 1564 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1712256841
transform 1 0 1524 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1712256841
transform 1 0 1268 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1712256841
transform 1 0 1196 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1712256841
transform 1 0 1108 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1712256841
transform 1 0 1020 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1712256841
transform 1 0 892 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1712256841
transform 1 0 644 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1712256841
transform 1 0 556 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1712256841
transform 1 0 388 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1712256841
transform 1 0 300 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1712256841
transform 1 0 260 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1712256841
transform 1 0 252 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1712256841
transform 1 0 252 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1712256841
transform 1 0 252 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1712256841
transform 1 0 236 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1712256841
transform 1 0 156 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1712256841
transform 1 0 156 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1712256841
transform 1 0 116 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1712256841
transform 1 0 2676 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1712256841
transform 1 0 2676 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1712256841
transform 1 0 2668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1712256841
transform 1 0 2628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1712256841
transform 1 0 2476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1712256841
transform 1 0 2460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1712256841
transform 1 0 2060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1712256841
transform 1 0 1876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1712256841
transform 1 0 1572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1712256841
transform 1 0 1284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1712256841
transform 1 0 1188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1712256841
transform 1 0 1188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1712256841
transform 1 0 1180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1712256841
transform 1 0 1164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1712256841
transform 1 0 2572 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1712256841
transform 1 0 2564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1712256841
transform 1 0 2460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1712256841
transform 1 0 2276 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1712256841
transform 1 0 2116 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1712256841
transform 1 0 2044 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1712256841
transform 1 0 2036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1712256841
transform 1 0 2004 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1712256841
transform 1 0 1804 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1712256841
transform 1 0 1636 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1712256841
transform 1 0 1596 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1712256841
transform 1 0 1516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1712256841
transform 1 0 1260 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1712256841
transform 1 0 1148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1712256841
transform 1 0 1140 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1712256841
transform 1 0 1132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1712256841
transform 1 0 1124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1712256841
transform 1 0 1124 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1712256841
transform 1 0 3308 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1712256841
transform 1 0 3252 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1712256841
transform 1 0 3180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1712256841
transform 1 0 1756 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1712256841
transform 1 0 1100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1712256841
transform 1 0 1044 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1712256841
transform 1 0 980 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1712256841
transform 1 0 740 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1712256841
transform 1 0 676 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1712256841
transform 1 0 572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1712256841
transform 1 0 428 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1712256841
transform 1 0 380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1712256841
transform 1 0 300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1712256841
transform 1 0 260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1712256841
transform 1 0 204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1712256841
transform 1 0 132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1712256841
transform 1 0 92 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1712256841
transform 1 0 2852 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1712256841
transform 1 0 2652 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1712256841
transform 1 0 2420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1712256841
transform 1 0 2300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1712256841
transform 1 0 2244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1712256841
transform 1 0 2084 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1712256841
transform 1 0 2020 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1712256841
transform 1 0 1988 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1712256841
transform 1 0 1844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1712256841
transform 1 0 1788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1712256841
transform 1 0 1676 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1712256841
transform 1 0 1468 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1712256841
transform 1 0 1396 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1712256841
transform 1 0 1364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1712256841
transform 1 0 3324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1712256841
transform 1 0 3276 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1712256841
transform 1 0 3268 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1712256841
transform 1 0 3156 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1712256841
transform 1 0 3092 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1712256841
transform 1 0 3028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1712256841
transform 1 0 2988 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1712256841
transform 1 0 2964 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1712256841
transform 1 0 2836 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1712256841
transform 1 0 2804 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1712256841
transform 1 0 2700 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1712256841
transform 1 0 2604 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1712256841
transform 1 0 2460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1712256841
transform 1 0 1316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1712256841
transform 1 0 1788 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1712256841
transform 1 0 1532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1712256841
transform 1 0 1308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1712256841
transform 1 0 1228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1712256841
transform 1 0 1196 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1712256841
transform 1 0 1004 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1712256841
transform 1 0 740 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1712256841
transform 1 0 700 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1712256841
transform 1 0 628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1712256841
transform 1 0 588 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1712256841
transform 1 0 588 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1712256841
transform 1 0 548 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1712256841
transform 1 0 508 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1712256841
transform 1 0 500 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1712256841
transform 1 0 2580 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1712256841
transform 1 0 2548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1712256841
transform 1 0 2404 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1712256841
transform 1 0 2292 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1712256841
transform 1 0 2212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1712256841
transform 1 0 2068 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1712256841
transform 1 0 2012 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1712256841
transform 1 0 1868 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1712256841
transform 1 0 1636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1712256841
transform 1 0 1572 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1712256841
transform 1 0 1492 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1712256841
transform 1 0 1420 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1712256841
transform 1 0 1332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1712256841
transform 1 0 972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1712256841
transform 1 0 3348 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1712256841
transform 1 0 3292 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1712256841
transform 1 0 3284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1712256841
transform 1 0 3260 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1712256841
transform 1 0 3244 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1712256841
transform 1 0 3228 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1712256841
transform 1 0 3188 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1712256841
transform 1 0 3180 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1712256841
transform 1 0 3140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1712256841
transform 1 0 3036 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1712256841
transform 1 0 3036 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1712256841
transform 1 0 2884 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1712256841
transform 1 0 2684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1712256841
transform 1 0 1628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1712256841
transform 1 0 1444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1712256841
transform 1 0 1404 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1712256841
transform 1 0 1364 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1712256841
transform 1 0 2876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1712256841
transform 1 0 2876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1712256841
transform 1 0 2804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1712256841
transform 1 0 2620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1712256841
transform 1 0 2532 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1712256841
transform 1 0 2412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1712256841
transform 1 0 2148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1712256841
transform 1 0 1612 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1712256841
transform 1 0 1572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1712256841
transform 1 0 1476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1712256841
transform 1 0 1452 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1712256841
transform 1 0 1380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1712256841
transform 1 0 1300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1712256841
transform 1 0 1204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1712256841
transform 1 0 1092 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1712256841
transform 1 0 996 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1712256841
transform 1 0 996 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1712256841
transform 1 0 980 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1712256841
transform 1 0 2620 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1712256841
transform 1 0 2580 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1712256841
transform 1 0 2548 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1712256841
transform 1 0 2540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1712256841
transform 1 0 2380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1712256841
transform 1 0 2380 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1712256841
transform 1 0 2380 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1712256841
transform 1 0 2380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1712256841
transform 1 0 2164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1712256841
transform 1 0 1804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1712256841
transform 1 0 1796 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1712256841
transform 1 0 1772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1712256841
transform 1 0 1660 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1712256841
transform 1 0 1660 0 1 695
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1712256841
transform 1 0 1364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1712256841
transform 1 0 1276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1712256841
transform 1 0 1108 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1712256841
transform 1 0 1076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1712256841
transform 1 0 1012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1712256841
transform 1 0 996 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1712256841
transform 1 0 884 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1712256841
transform 1 0 820 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1712256841
transform 1 0 812 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1712256841
transform 1 0 812 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1712256841
transform 1 0 3092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1712256841
transform 1 0 3060 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1712256841
transform 1 0 3036 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1712256841
transform 1 0 3020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1712256841
transform 1 0 2444 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1712256841
transform 1 0 2188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1712256841
transform 1 0 2164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1712256841
transform 1 0 2052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1712256841
transform 1 0 1980 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1712256841
transform 1 0 1956 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1712256841
transform 1 0 1956 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1712256841
transform 1 0 1924 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1712256841
transform 1 0 3060 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1712256841
transform 1 0 2948 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1712256841
transform 1 0 2940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1712256841
transform 1 0 2708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1712256841
transform 1 0 2116 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1712256841
transform 1 0 2092 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1712256841
transform 1 0 1972 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1712256841
transform 1 0 1876 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1712256841
transform 1 0 1764 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1712256841
transform 1 0 1740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1712256841
transform 1 0 1724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1712256841
transform 1 0 2428 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1712256841
transform 1 0 2412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1712256841
transform 1 0 2372 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1712256841
transform 1 0 2308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1712256841
transform 1 0 2276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1712256841
transform 1 0 2276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1712256841
transform 1 0 2212 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1712256841
transform 1 0 2204 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1712256841
transform 1 0 2156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1712256841
transform 1 0 2084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1712256841
transform 1 0 2228 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1712256841
transform 1 0 2172 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1712256841
transform 1 0 2132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1712256841
transform 1 0 2108 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1712256841
transform 1 0 1916 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1712256841
transform 1 0 1884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1712256841
transform 1 0 1772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1712256841
transform 1 0 1764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1712256841
transform 1 0 1748 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1712256841
transform 1 0 1628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1712256841
transform 1 0 1628 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1712256841
transform 1 0 2348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1712256841
transform 1 0 2276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1712256841
transform 1 0 2244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1712256841
transform 1 0 1668 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1712256841
transform 1 0 1532 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1712256841
transform 1 0 1356 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1712256841
transform 1 0 1212 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1712256841
transform 1 0 1060 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1712256841
transform 1 0 772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1712256841
transform 1 0 764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1712256841
transform 1 0 668 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1712256841
transform 1 0 1364 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1712256841
transform 1 0 1316 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1712256841
transform 1 0 1316 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1712256841
transform 1 0 1276 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1712256841
transform 1 0 1276 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1712256841
transform 1 0 1236 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1712256841
transform 1 0 1236 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1712256841
transform 1 0 980 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1712256841
transform 1 0 948 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1712256841
transform 1 0 940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1712256841
transform 1 0 916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1712256841
transform 1 0 884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1712256841
transform 1 0 860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1712256841
transform 1 0 788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1712256841
transform 1 0 780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1712256841
transform 1 0 764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1712256841
transform 1 0 636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1712256841
transform 1 0 620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1712256841
transform 1 0 580 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1712256841
transform 1 0 580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1712256841
transform 1 0 564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1712256841
transform 1 0 396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1712256841
transform 1 0 236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1712256841
transform 1 0 196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1712256841
transform 1 0 1700 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1712256841
transform 1 0 1660 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1712256841
transform 1 0 1396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1712256841
transform 1 0 1204 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1712256841
transform 1 0 764 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1712256841
transform 1 0 372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1712256841
transform 1 0 372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1712256841
transform 1 0 340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1712256841
transform 1 0 308 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1712256841
transform 1 0 252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1712256841
transform 1 0 220 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1712256841
transform 1 0 924 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1712256841
transform 1 0 852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1712256841
transform 1 0 772 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1712256841
transform 1 0 588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1712256841
transform 1 0 460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1712256841
transform 1 0 444 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1712256841
transform 1 0 364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1712256841
transform 1 0 324 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1712256841
transform 1 0 300 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1712256841
transform 1 0 108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1712256841
transform 1 0 1260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1712256841
transform 1 0 1220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1712256841
transform 1 0 700 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1712256841
transform 1 0 612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1712256841
transform 1 0 508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1712256841
transform 1 0 300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1712256841
transform 1 0 300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1712256841
transform 1 0 292 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1712256841
transform 1 0 236 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1712256841
transform 1 0 236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1712256841
transform 1 0 1372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1712256841
transform 1 0 1332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1712256841
transform 1 0 1332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1712256841
transform 1 0 1316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1712256841
transform 1 0 1300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1712256841
transform 1 0 1300 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1712256841
transform 1 0 1292 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1712256841
transform 1 0 1284 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1712256841
transform 1 0 1204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1712256841
transform 1 0 1140 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1712256841
transform 1 0 1092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1712256841
transform 1 0 1092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1712256841
transform 1 0 924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1712256841
transform 1 0 852 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1712256841
transform 1 0 788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1712256841
transform 1 0 780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1712256841
transform 1 0 684 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1712256841
transform 1 0 684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1712256841
transform 1 0 652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1712256841
transform 1 0 3388 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1712256841
transform 1 0 3380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1712256841
transform 1 0 3356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1712256841
transform 1 0 3348 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1712256841
transform 1 0 3260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1712256841
transform 1 0 3220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1712256841
transform 1 0 3212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1712256841
transform 1 0 3188 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1712256841
transform 1 0 3092 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1712256841
transform 1 0 3396 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1712256841
transform 1 0 3172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1712256841
transform 1 0 3132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1712256841
transform 1 0 3116 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1712256841
transform 1 0 3308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1712256841
transform 1 0 2948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1712256841
transform 1 0 2644 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1712256841
transform 1 0 1764 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1712256841
transform 1 0 3252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1712256841
transform 1 0 3100 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1712256841
transform 1 0 2564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1712256841
transform 1 0 2484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1712256841
transform 1 0 2692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1712256841
transform 1 0 2652 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1712256841
transform 1 0 2636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1712256841
transform 1 0 2588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1712256841
transform 1 0 1668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1712256841
transform 1 0 1668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1712256841
transform 1 0 1652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1712256841
transform 1 0 1636 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1712256841
transform 1 0 1412 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1712256841
transform 1 0 1108 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1712256841
transform 1 0 1444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1712256841
transform 1 0 1412 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1712256841
transform 1 0 1316 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1712256841
transform 1 0 1220 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1712256841
transform 1 0 1204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1712256841
transform 1 0 2940 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1712256841
transform 1 0 2924 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1712256841
transform 1 0 2924 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1712256841
transform 1 0 2860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1712256841
transform 1 0 2660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1712256841
transform 1 0 2388 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1712256841
transform 1 0 1532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1712256841
transform 1 0 1532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1712256841
transform 1 0 1516 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1712256841
transform 1 0 1484 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1712256841
transform 1 0 1388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1712256841
transform 1 0 3228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1712256841
transform 1 0 3172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1712256841
transform 1 0 3140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1712256841
transform 1 0 3108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1712256841
transform 1 0 3060 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1712256841
transform 1 0 3220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1712256841
transform 1 0 2796 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1712256841
transform 1 0 1636 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1712256841
transform 1 0 3332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1712256841
transform 1 0 3252 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1712256841
transform 1 0 3164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1712256841
transform 1 0 3148 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1712256841
transform 1 0 3196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1712256841
transform 1 0 2324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1712256841
transform 1 0 2868 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1712256841
transform 1 0 2836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1712256841
transform 1 0 3388 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1712256841
transform 1 0 3388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1712256841
transform 1 0 3340 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1712256841
transform 1 0 3332 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1712256841
transform 1 0 1468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1712256841
transform 1 0 1292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1712256841
transform 1 0 1292 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1712256841
transform 1 0 1212 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1712256841
transform 1 0 1164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1712256841
transform 1 0 1436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1712256841
transform 1 0 1380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1712256841
transform 1 0 852 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1712256841
transform 1 0 756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1712256841
transform 1 0 756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1712256841
transform 1 0 1348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1712256841
transform 1 0 1252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1712256841
transform 1 0 1220 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1712256841
transform 1 0 1036 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1712256841
transform 1 0 1020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1712256841
transform 1 0 1020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1712256841
transform 1 0 1004 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1712256841
transform 1 0 964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1712256841
transform 1 0 868 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1712256841
transform 1 0 2332 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1712256841
transform 1 0 2332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1712256841
transform 1 0 2244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1712256841
transform 1 0 2244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1712256841
transform 1 0 2084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1712256841
transform 1 0 1916 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1712256841
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1712256841
transform 1 0 1612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1712256841
transform 1 0 1604 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1712256841
transform 1 0 1532 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1712256841
transform 1 0 1436 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1712256841
transform 1 0 1420 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1712256841
transform 1 0 964 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1712256841
transform 1 0 724 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1712256841
transform 1 0 1052 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1712256841
transform 1 0 636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1712256841
transform 1 0 564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1712256841
transform 1 0 500 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1712256841
transform 1 0 468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1712256841
transform 1 0 276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1712256841
transform 1 0 236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1712256841
transform 1 0 3036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1712256841
transform 1 0 3036 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1712256841
transform 1 0 2996 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1712256841
transform 1 0 2684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1712256841
transform 1 0 2636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1712256841
transform 1 0 2116 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1712256841
transform 1 0 1956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1712256841
transform 1 0 1028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1712256841
transform 1 0 828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1712256841
transform 1 0 596 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1712256841
transform 1 0 564 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1712256841
transform 1 0 356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1712256841
transform 1 0 260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1712256841
transform 1 0 212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1712256841
transform 1 0 2700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1712256841
transform 1 0 2596 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1712256841
transform 1 0 2492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1712256841
transform 1 0 2484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1712256841
transform 1 0 2444 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1712256841
transform 1 0 2444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1712256841
transform 1 0 2276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1712256841
transform 1 0 2172 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1712256841
transform 1 0 2092 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1712256841
transform 1 0 2036 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1712256841
transform 1 0 1860 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1712256841
transform 1 0 1852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1712256841
transform 1 0 1724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1712256841
transform 1 0 1628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1712256841
transform 1 0 1332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1712256841
transform 1 0 1300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1712256841
transform 1 0 1100 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1712256841
transform 1 0 964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1712256841
transform 1 0 716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1712256841
transform 1 0 452 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1712256841
transform 1 0 444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1712256841
transform 1 0 436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1712256841
transform 1 0 420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1712256841
transform 1 0 420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1712256841
transform 1 0 420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1712256841
transform 1 0 396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1712256841
transform 1 0 396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1712256841
transform 1 0 348 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1712256841
transform 1 0 2716 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1712256841
transform 1 0 2692 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1712256841
transform 1 0 2668 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1712256841
transform 1 0 2588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1712256841
transform 1 0 2204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1712256841
transform 1 0 2196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1712256841
transform 1 0 2188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1712256841
transform 1 0 2188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1712256841
transform 1 0 3372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1712256841
transform 1 0 3276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1712256841
transform 1 0 3276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1712256841
transform 1 0 3268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1712256841
transform 1 0 3156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1712256841
transform 1 0 3148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1712256841
transform 1 0 3052 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1712256841
transform 1 0 2972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1712256841
transform 1 0 2868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1712256841
transform 1 0 2844 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1712256841
transform 1 0 3356 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1712256841
transform 1 0 3316 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1712256841
transform 1 0 3188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1712256841
transform 1 0 3180 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1712256841
transform 1 0 3004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1712256841
transform 1 0 2988 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1712256841
transform 1 0 2940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1712256841
transform 1 0 2892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1712256841
transform 1 0 3436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1712256841
transform 1 0 3388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1712256841
transform 1 0 3276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1712256841
transform 1 0 3268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1712256841
transform 1 0 3148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1712256841
transform 1 0 3140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1712256841
transform 1 0 3044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1712256841
transform 1 0 3036 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1712256841
transform 1 0 2964 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1712256841
transform 1 0 2908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1712256841
transform 1 0 3396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1712256841
transform 1 0 3388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1712256841
transform 1 0 3412 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1712256841
transform 1 0 3372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1712256841
transform 1 0 3420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1712256841
transform 1 0 3372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1712256841
transform 1 0 3356 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1712256841
transform 1 0 2964 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1712256841
transform 1 0 2876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1712256841
transform 1 0 2780 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1712256841
transform 1 0 2724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1712256841
transform 1 0 3348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1712256841
transform 1 0 3276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1712256841
transform 1 0 2772 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1712256841
transform 1 0 2676 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1712256841
transform 1 0 2676 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1712256841
transform 1 0 2676 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1712256841
transform 1 0 2652 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1712256841
transform 1 0 3196 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1712256841
transform 1 0 2788 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1712256841
transform 1 0 2724 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1712256841
transform 1 0 2628 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1712256841
transform 1 0 2612 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1712256841
transform 1 0 2604 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1712256841
transform 1 0 3204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1712256841
transform 1 0 3108 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1712256841
transform 1 0 2732 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1712256841
transform 1 0 2708 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1712256841
transform 1 0 2692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1712256841
transform 1 0 2692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1712256841
transform 1 0 2684 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1712256841
transform 1 0 2580 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1712256841
transform 1 0 2580 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1712256841
transform 1 0 2940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1712256841
transform 1 0 2828 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1712256841
transform 1 0 2796 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1712256841
transform 1 0 2724 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1712256841
transform 1 0 2692 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1712256841
transform 1 0 2796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1712256841
transform 1 0 2780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1712256841
transform 1 0 2772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1712256841
transform 1 0 2756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1712256841
transform 1 0 2740 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1712256841
transform 1 0 2700 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1712256841
transform 1 0 3364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1712256841
transform 1 0 3364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1712256841
transform 1 0 3260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1712256841
transform 1 0 3060 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1712256841
transform 1 0 3196 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1712256841
transform 1 0 3172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1712256841
transform 1 0 3004 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1712256841
transform 1 0 2980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1712256841
transform 1 0 2852 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1712256841
transform 1 0 2852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1712256841
transform 1 0 3372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1712256841
transform 1 0 3300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1712256841
transform 1 0 3284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1712256841
transform 1 0 3228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1712256841
transform 1 0 2724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1712256841
transform 1 0 2716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1712256841
transform 1 0 2892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1712256841
transform 1 0 2892 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1712256841
transform 1 0 2996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1712256841
transform 1 0 2996 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1712256841
transform 1 0 2844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1712256841
transform 1 0 2820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1712256841
transform 1 0 2628 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1712256841
transform 1 0 2628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1712256841
transform 1 0 2508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1712256841
transform 1 0 2508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1712256841
transform 1 0 2444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1712256841
transform 1 0 2436 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1712256841
transform 1 0 2124 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1712256841
transform 1 0 2108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1712256841
transform 1 0 2012 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1712256841
transform 1 0 1956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1712256841
transform 1 0 2324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1712256841
transform 1 0 2324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1712256841
transform 1 0 2268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1712256841
transform 1 0 2244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1712256841
transform 1 0 2140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1712256841
transform 1 0 2052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1712256841
transform 1 0 1892 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1712256841
transform 1 0 1860 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1712256841
transform 1 0 1828 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1712256841
transform 1 0 1756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1712256841
transform 1 0 1700 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1712256841
transform 1 0 1644 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1712256841
transform 1 0 1508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1712256841
transform 1 0 1508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1712256841
transform 1 0 1492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1712256841
transform 1 0 1468 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1712256841
transform 1 0 1388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1712256841
transform 1 0 1364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1712256841
transform 1 0 1148 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1712256841
transform 1 0 1140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1712256841
transform 1 0 1028 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1712256841
transform 1 0 980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1712256841
transform 1 0 804 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1712256841
transform 1 0 652 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1712256841
transform 1 0 188 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1712256841
transform 1 0 188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1712256841
transform 1 0 124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1712256841
transform 1 0 124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1712256841
transform 1 0 252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1712256841
transform 1 0 132 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1712256841
transform 1 0 284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1712256841
transform 1 0 268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1712256841
transform 1 0 364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1712256841
transform 1 0 348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1712256841
transform 1 0 420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1712256841
transform 1 0 380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1712256841
transform 1 0 492 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1712256841
transform 1 0 492 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1712256841
transform 1 0 724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1712256841
transform 1 0 604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1712256841
transform 1 0 796 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1712256841
transform 1 0 708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1712256841
transform 1 0 1092 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1712256841
transform 1 0 940 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1712256841
transform 1 0 1340 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1712256841
transform 1 0 1252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1712256841
transform 1 0 2988 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1712256841
transform 1 0 2972 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1712256841
transform 1 0 2092 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1712256841
transform 1 0 1636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1712256841
transform 1 0 2540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1712256841
transform 1 0 2524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1712256841
transform 1 0 3412 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1712256841
transform 1 0 3372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1712256841
transform 1 0 3196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1712256841
transform 1 0 3100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1712256841
transform 1 0 2964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1712256841
transform 1 0 2940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1712256841
transform 1 0 3228 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1712256841
transform 1 0 3228 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1712256841
transform 1 0 3180 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1712256841
transform 1 0 2756 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1712256841
transform 1 0 2676 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1712256841
transform 1 0 2564 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1712256841
transform 1 0 3412 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1712256841
transform 1 0 3372 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1712256841
transform 1 0 3308 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1712256841
transform 1 0 3340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1712256841
transform 1 0 3300 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1712256841
transform 1 0 3284 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1712256841
transform 1 0 2900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1712256841
transform 1 0 1612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1712256841
transform 1 0 1692 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1712256841
transform 1 0 1580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1712256841
transform 1 0 1572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1712256841
transform 1 0 1500 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1712256841
transform 1 0 1452 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1712256841
transform 1 0 1452 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1712256841
transform 1 0 1532 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1712256841
transform 1 0 1444 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1712256841
transform 1 0 1492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1712256841
transform 1 0 1468 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1712256841
transform 1 0 1572 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1712256841
transform 1 0 1484 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1712256841
transform 1 0 1532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1712256841
transform 1 0 1532 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1712256841
transform 1 0 1508 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1712256841
transform 1 0 1476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1712256841
transform 1 0 2116 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1712256841
transform 1 0 1508 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1712256841
transform 1 0 1492 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1712256841
transform 1 0 860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1712256841
transform 1 0 836 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1712256841
transform 1 0 268 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1712256841
transform 1 0 868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1712256841
transform 1 0 860 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1712256841
transform 1 0 860 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1712256841
transform 1 0 860 0 1 1885
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1712256841
transform 1 0 1044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1712256841
transform 1 0 844 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1712256841
transform 1 0 844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1712256841
transform 1 0 668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1712256841
transform 1 0 852 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1712256841
transform 1 0 852 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1712256841
transform 1 0 1724 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1712256841
transform 1 0 828 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1712256841
transform 1 0 660 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1712256841
transform 1 0 1020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1712256841
transform 1 0 868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1712256841
transform 1 0 1540 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1712256841
transform 1 0 1508 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1712256841
transform 1 0 1476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1712256841
transform 1 0 1300 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1712256841
transform 1 0 1004 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1712256841
transform 1 0 1324 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1712256841
transform 1 0 1196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1712256841
transform 1 0 1044 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1712256841
transform 1 0 1036 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1712256841
transform 1 0 660 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1712256841
transform 1 0 524 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1712256841
transform 1 0 356 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1712256841
transform 1 0 740 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1712256841
transform 1 0 684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1712256841
transform 1 0 588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1712256841
transform 1 0 1172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1712256841
transform 1 0 1012 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1712256841
transform 1 0 972 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1712256841
transform 1 0 900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1712256841
transform 1 0 1284 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1712256841
transform 1 0 1108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1712256841
transform 1 0 1108 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1712256841
transform 1 0 1084 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1712256841
transform 1 0 220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1712256841
transform 1 0 180 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1712256841
transform 1 0 236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1712256841
transform 1 0 196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1712256841
transform 1 0 300 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1712256841
transform 1 0 188 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1712256841
transform 1 0 268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1712256841
transform 1 0 268 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1712256841
transform 1 0 180 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1712256841
transform 1 0 300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1712256841
transform 1 0 292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1712256841
transform 1 0 324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1712256841
transform 1 0 236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1712256841
transform 1 0 204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1712256841
transform 1 0 524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1712256841
transform 1 0 308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1712256841
transform 1 0 308 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1712256841
transform 1 0 284 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1712256841
transform 1 0 284 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1712256841
transform 1 0 244 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1712256841
transform 1 0 220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1712256841
transform 1 0 180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1712256841
transform 1 0 268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1712256841
transform 1 0 212 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1712256841
transform 1 0 204 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1712256841
transform 1 0 540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1712256841
transform 1 0 180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1712256841
transform 1 0 156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1712256841
transform 1 0 252 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1712256841
transform 1 0 252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1712256841
transform 1 0 220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1712256841
transform 1 0 2108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1712256841
transform 1 0 2108 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1712256841
transform 1 0 2212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1712256841
transform 1 0 2180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1712256841
transform 1 0 2252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1712256841
transform 1 0 2228 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1712256841
transform 1 0 2220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1712256841
transform 1 0 1820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1712256841
transform 1 0 1780 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1712256841
transform 1 0 2276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1712256841
transform 1 0 2268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1712256841
transform 1 0 2260 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1712256841
transform 1 0 2268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1712256841
transform 1 0 2164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1712256841
transform 1 0 2164 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1712256841
transform 1 0 2092 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1712256841
transform 1 0 2084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1712256841
transform 1 0 2332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1712256841
transform 1 0 2116 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1712256841
transform 1 0 2404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1712256841
transform 1 0 2324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1712256841
transform 1 0 2324 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1712256841
transform 1 0 2324 0 1 685
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1712256841
transform 1 0 2300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1712256841
transform 1 0 2404 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1712256841
transform 1 0 2404 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1712256841
transform 1 0 2340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1712256841
transform 1 0 2212 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1712256841
transform 1 0 2164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1712256841
transform 1 0 2084 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1712256841
transform 1 0 2100 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1712256841
transform 1 0 1908 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1712256841
transform 1 0 1860 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1712256841
transform 1 0 1500 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1712256841
transform 1 0 1484 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1712256841
transform 1 0 1500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1712256841
transform 1 0 1116 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1712256841
transform 1 0 1108 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1712256841
transform 1 0 1020 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1712256841
transform 1 0 1140 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1712256841
transform 1 0 1052 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1712256841
transform 1 0 1012 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1712256841
transform 1 0 1028 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1712256841
transform 1 0 892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1712256841
transform 1 0 892 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1712256841
transform 1 0 444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1712256841
transform 1 0 428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1712256841
transform 1 0 332 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1712256841
transform 1 0 1612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1712256841
transform 1 0 1516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1712256841
transform 1 0 2228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1712256841
transform 1 0 1564 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1712256841
transform 1 0 2492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1712256841
transform 1 0 2388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1712256841
transform 1 0 2212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1712256841
transform 1 0 2284 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1712256841
transform 1 0 2236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1712256841
transform 1 0 2180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1712256841
transform 1 0 1740 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1712256841
transform 1 0 1708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1712256841
transform 1 0 1604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1712256841
transform 1 0 1620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1712256841
transform 1 0 1420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1712256841
transform 1 0 1380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1712256841
transform 1 0 1812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1712256841
transform 1 0 1516 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1712256841
transform 1 0 1660 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1712256841
transform 1 0 1548 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1712256841
transform 1 0 1516 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1712256841
transform 1 0 644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1712256841
transform 1 0 588 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1712256841
transform 1 0 540 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1712256841
transform 1 0 612 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1712256841
transform 1 0 500 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1712256841
transform 1 0 412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1712256841
transform 1 0 404 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1712256841
transform 1 0 460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1712256841
transform 1 0 412 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1712256841
transform 1 0 668 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1712256841
transform 1 0 444 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1712256841
transform 1 0 796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1712256841
transform 1 0 684 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1712256841
transform 1 0 924 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1712256841
transform 1 0 916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1712256841
transform 1 0 780 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1712256841
transform 1 0 820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1712256841
transform 1 0 820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1712256841
transform 1 0 780 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1712256841
transform 1 0 2964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1712256841
transform 1 0 2844 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1712256841
transform 1 0 2580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1712256841
transform 1 0 2564 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1712256841
transform 1 0 2556 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1712256841
transform 1 0 2476 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1712256841
transform 1 0 1652 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1712256841
transform 1 0 1516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1712256841
transform 1 0 1516 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1712256841
transform 1 0 2596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1712256841
transform 1 0 2540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1712256841
transform 1 0 1684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1712256841
transform 1 0 484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1712256841
transform 1 0 444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1712256841
transform 1 0 404 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1712256841
transform 1 0 444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1712256841
transform 1 0 420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1712256841
transform 1 0 388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1712256841
transform 1 0 388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1712256841
transform 1 0 380 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1712256841
transform 1 0 492 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1712256841
transform 1 0 452 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1712256841
transform 1 0 444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1712256841
transform 1 0 468 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1712256841
transform 1 0 444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1712256841
transform 1 0 980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1712256841
transform 1 0 516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1712256841
transform 1 0 508 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1712256841
transform 1 0 508 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1712256841
transform 1 0 484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1712256841
transform 1 0 468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1712256841
transform 1 0 436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1712256841
transform 1 0 452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1712256841
transform 1 0 444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1712256841
transform 1 0 476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1712256841
transform 1 0 460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1712256841
transform 1 0 436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1712256841
transform 1 0 468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1712256841
transform 1 0 468 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1712256841
transform 1 0 1124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1712256841
transform 1 0 1012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1712256841
transform 1 0 972 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1712256841
transform 1 0 988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1712256841
transform 1 0 988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1712256841
transform 1 0 956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1712256841
transform 1 0 500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1712256841
transform 1 0 412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1712256841
transform 1 0 452 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1712256841
transform 1 0 420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1712256841
transform 1 0 420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1712256841
transform 1 0 1780 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1712256841
transform 1 0 1636 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1712256841
transform 1 0 1748 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1712256841
transform 1 0 1668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1712256841
transform 1 0 1748 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1712256841
transform 1 0 1716 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1712256841
transform 1 0 1716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1712256841
transform 1 0 1748 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1712256841
transform 1 0 1588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1712256841
transform 1 0 1572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1712256841
transform 1 0 1468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1712256841
transform 1 0 1244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1712256841
transform 1 0 932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1712256841
transform 1 0 596 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1712256841
transform 1 0 1548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1712256841
transform 1 0 1348 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1712256841
transform 1 0 1332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1712256841
transform 1 0 1604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1712256841
transform 1 0 1572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1712256841
transform 1 0 1388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1712256841
transform 1 0 996 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1712256841
transform 1 0 644 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1712256841
transform 1 0 164 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1712256841
transform 1 0 156 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1712256841
transform 1 0 1596 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1712256841
transform 1 0 1596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1712256841
transform 1 0 1588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1712256841
transform 1 0 1764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1712256841
transform 1 0 1740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1712256841
transform 1 0 2140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1712256841
transform 1 0 1820 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1712256841
transform 1 0 2500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1712256841
transform 1 0 2324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1712256841
transform 1 0 2132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1712256841
transform 1 0 2124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1712256841
transform 1 0 2380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1712256841
transform 1 0 2340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1712256841
transform 1 0 2132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1712256841
transform 1 0 2588 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1712256841
transform 1 0 2244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1712256841
transform 1 0 2172 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1712256841
transform 1 0 2164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1712256841
transform 1 0 2164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1712256841
transform 1 0 2228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1712256841
transform 1 0 2196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1712256841
transform 1 0 2196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1712256841
transform 1 0 2548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1712256841
transform 1 0 2140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1712256841
transform 1 0 1836 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1712256841
transform 1 0 1828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1712256841
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1712256841
transform 1 0 1940 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1712256841
transform 1 0 1924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1712256841
transform 1 0 1732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1712256841
transform 1 0 1652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1712256841
transform 1 0 1316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1712256841
transform 1 0 1316 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1712256841
transform 1 0 2548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1712256841
transform 1 0 1828 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1712256841
transform 1 0 1860 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1712256841
transform 1 0 1852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1712256841
transform 1 0 1804 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1712256841
transform 1 0 1372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1712256841
transform 1 0 1372 0 1 355
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1712256841
transform 1 0 2156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1712256841
transform 1 0 2156 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1712256841
transform 1 0 1884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1712256841
transform 1 0 1844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1712256841
transform 1 0 1796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1712256841
transform 1 0 1692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1712256841
transform 1 0 1556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1712256841
transform 1 0 1980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1712256841
transform 1 0 1900 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1712256841
transform 1 0 2148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1712256841
transform 1 0 2100 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1712256841
transform 1 0 1972 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1712256841
transform 1 0 1988 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1712256841
transform 1 0 1876 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1712256841
transform 1 0 1772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1712256841
transform 1 0 2636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1712256841
transform 1 0 2524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1712256841
transform 1 0 2540 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1712256841
transform 1 0 2540 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1712256841
transform 1 0 2620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1712256841
transform 1 0 2516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1712256841
transform 1 0 2508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1712256841
transform 1 0 2548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1712256841
transform 1 0 2500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1712256841
transform 1 0 2356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1712256841
transform 1 0 2660 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1712256841
transform 1 0 2508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1712256841
transform 1 0 2420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1712256841
transform 1 0 1596 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1712256841
transform 1 0 1508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1712256841
transform 1 0 1484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1712256841
transform 1 0 948 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1712256841
transform 1 0 884 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1712256841
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1712256841
transform 1 0 924 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1712256841
transform 1 0 884 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1712256841
transform 1 0 900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1712256841
transform 1 0 900 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1712256841
transform 1 0 868 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1712256841
transform 1 0 588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1712256841
transform 1 0 1556 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1712256841
transform 1 0 916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1712256841
transform 1 0 1556 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1712256841
transform 1 0 1028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1712256841
transform 1 0 1108 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1712256841
transform 1 0 980 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1712256841
transform 1 0 932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1712256841
transform 1 0 1212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1712256841
transform 1 0 1052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1712256841
transform 1 0 1020 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1712256841
transform 1 0 2556 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1712256841
transform 1 0 2524 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1712256841
transform 1 0 1556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1712256841
transform 1 0 532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1712256841
transform 1 0 484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1712256841
transform 1 0 580 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1712256841
transform 1 0 516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1712256841
transform 1 0 668 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1712256841
transform 1 0 564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1712256841
transform 1 0 500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1712256841
transform 1 0 532 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1712256841
transform 1 0 532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1712256841
transform 1 0 628 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1712256841
transform 1 0 556 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1712256841
transform 1 0 500 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1712256841
transform 1 0 468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1712256841
transform 1 0 652 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1712256841
transform 1 0 540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1712256841
transform 1 0 540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1712256841
transform 1 0 1004 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1712256841
transform 1 0 868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1712256841
transform 1 0 884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1712256841
transform 1 0 724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1712256841
transform 1 0 780 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1712256841
transform 1 0 780 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1712256841
transform 1 0 740 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1712256841
transform 1 0 716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1712256841
transform 1 0 732 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1712256841
transform 1 0 732 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1712256841
transform 1 0 628 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1712256841
transform 1 0 988 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1712256841
transform 1 0 988 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1712256841
transform 1 0 956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1712256841
transform 1 0 932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1712256841
transform 1 0 1076 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1712256841
transform 1 0 1060 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1712256841
transform 1 0 1052 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1712256841
transform 1 0 1988 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1712256841
transform 1 0 1988 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1712256841
transform 1 0 1820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1712256841
transform 1 0 1404 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1712256841
transform 1 0 1316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1712256841
transform 1 0 1252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1712256841
transform 1 0 1244 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1712256841
transform 1 0 612 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1712256841
transform 1 0 508 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1712256841
transform 1 0 508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1712256841
transform 1 0 540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1712256841
transform 1 0 532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1712256841
transform 1 0 596 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1712256841
transform 1 0 508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1712256841
transform 1 0 508 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1712256841
transform 1 0 692 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1712256841
transform 1 0 612 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1712256841
transform 1 0 1572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1712256841
transform 1 0 1572 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1712256841
transform 1 0 2132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1712256841
transform 1 0 1580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1712256841
transform 1 0 1732 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1712256841
transform 1 0 1588 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1712256841
transform 1 0 2396 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1712256841
transform 1 0 1708 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1712256841
transform 1 0 1724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1712256841
transform 1 0 1724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1712256841
transform 1 0 1956 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1712256841
transform 1 0 1748 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1712256841
transform 1 0 2028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1712256841
transform 1 0 1924 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1712256841
transform 1 0 1924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1712256841
transform 1 0 1972 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1712256841
transform 1 0 1820 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1712256841
transform 1 0 2276 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1712256841
transform 1 0 2244 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1712256841
transform 1 0 2212 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1712256841
transform 1 0 2124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1712256841
transform 1 0 2124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1712256841
transform 1 0 2044 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1712256841
transform 1 0 2004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1712256841
transform 1 0 2004 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1712256841
transform 1 0 1980 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1712256841
transform 1 0 1948 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1712256841
transform 1 0 1564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1712256841
transform 1 0 1444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1712256841
transform 1 0 2436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1712256841
transform 1 0 2412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1712256841
transform 1 0 2460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1712256841
transform 1 0 2452 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1712256841
transform 1 0 2428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1712256841
transform 1 0 2404 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1712256841
transform 1 0 1996 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1712256841
transform 1 0 2476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1712256841
transform 1 0 2356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1712256841
transform 1 0 2140 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1712256841
transform 1 0 2404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1712256841
transform 1 0 2356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1712256841
transform 1 0 2132 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1712256841
transform 1 0 2452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1712256841
transform 1 0 2268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1712256841
transform 1 0 2076 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1712256841
transform 1 0 2356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1712256841
transform 1 0 2108 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1712256841
transform 1 0 2156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1712256841
transform 1 0 2116 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1712256841
transform 1 0 2180 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1712256841
transform 1 0 2140 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1712256841
transform 1 0 1996 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1712256841
transform 1 0 2252 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1712256841
transform 1 0 2220 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1712256841
transform 1 0 2204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1712256841
transform 1 0 2476 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1712256841
transform 1 0 2340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1712256841
transform 1 0 2332 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1712256841
transform 1 0 1532 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1712256841
transform 1 0 1260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1712256841
transform 1 0 1628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1712256841
transform 1 0 1548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1712256841
transform 1 0 1740 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1712256841
transform 1 0 1668 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1712256841
transform 1 0 1620 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1712256841
transform 1 0 1636 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1712256841
transform 1 0 1540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1712256841
transform 1 0 1332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1712256841
transform 1 0 1252 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1712256841
transform 1 0 1236 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1712256841
transform 1 0 1068 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1712256841
transform 1 0 1268 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1712256841
transform 1 0 1156 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1712256841
transform 1 0 1124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1712256841
transform 1 0 1476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1712256841
transform 1 0 1388 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1712256841
transform 1 0 1028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1712256841
transform 1 0 588 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1712256841
transform 1 0 564 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1712256841
transform 1 0 156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1712256841
transform 1 0 140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1712256841
transform 1 0 1964 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1712256841
transform 1 0 1388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1712256841
transform 1 0 1404 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1712256841
transform 1 0 772 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1712256841
transform 1 0 708 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1712256841
transform 1 0 668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1712256841
transform 1 0 716 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1712256841
transform 1 0 716 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1712256841
transform 1 0 788 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1712256841
transform 1 0 756 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1712256841
transform 1 0 908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1712256841
transform 1 0 812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1712256841
transform 1 0 1244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1712256841
transform 1 0 1244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1712256841
transform 1 0 924 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1712256841
transform 1 0 868 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1712256841
transform 1 0 868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1712256841
transform 1 0 332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1712256841
transform 1 0 260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1712256841
transform 1 0 908 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1712256841
transform 1 0 884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1712256841
transform 1 0 1092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1712256841
transform 1 0 1028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1712256841
transform 1 0 924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1712256841
transform 1 0 860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1712256841
transform 1 0 932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1712256841
transform 1 0 892 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1712256841
transform 1 0 892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1712256841
transform 1 0 948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1712256841
transform 1 0 756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1712256841
transform 1 0 772 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1712256841
transform 1 0 692 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1712256841
transform 1 0 1012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1712256841
transform 1 0 844 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1712256841
transform 1 0 740 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1712256841
transform 1 0 644 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1712256841
transform 1 0 604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1712256841
transform 1 0 740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1712256841
transform 1 0 732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1712256841
transform 1 0 708 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1712256841
transform 1 0 700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1712256841
transform 1 0 676 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1712256841
transform 1 0 604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1712256841
transform 1 0 1156 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1712256841
transform 1 0 1060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1712256841
transform 1 0 996 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1712256841
transform 1 0 916 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1712256841
transform 1 0 916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1712256841
transform 1 0 900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1712256841
transform 1 0 900 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1712256841
transform 1 0 1356 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1712256841
transform 1 0 1268 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1712256841
transform 1 0 1060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1712256841
transform 1 0 980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1712256841
transform 1 0 980 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1712256841
transform 1 0 764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1712256841
transform 1 0 700 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1712256841
transform 1 0 644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1712256841
transform 1 0 572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1712256841
transform 1 0 836 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1712256841
transform 1 0 772 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1712256841
transform 1 0 700 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1712256841
transform 1 0 564 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1712256841
transform 1 0 564 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1712256841
transform 1 0 540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1712256841
transform 1 0 524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1712256841
transform 1 0 964 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1712256841
transform 1 0 884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1712256841
transform 1 0 644 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1712256841
transform 1 0 628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1712256841
transform 1 0 620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1712256841
transform 1 0 2524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1712256841
transform 1 0 2492 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1712256841
transform 1 0 2412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1712256841
transform 1 0 2380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1712256841
transform 1 0 1468 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1712256841
transform 1 0 1164 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1712256841
transform 1 0 1044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1712256841
transform 1 0 1004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1712256841
transform 1 0 1004 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1712256841
transform 1 0 732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1712256841
transform 1 0 700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1712256841
transform 1 0 660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1712256841
transform 1 0 652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1712256841
transform 1 0 1092 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1712256841
transform 1 0 940 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1712256841
transform 1 0 700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1712256841
transform 1 0 636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1712256841
transform 1 0 588 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1712256841
transform 1 0 588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1712256841
transform 1 0 852 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1712256841
transform 1 0 852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1712256841
transform 1 0 812 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1712256841
transform 1 0 756 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1712256841
transform 1 0 580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1712256841
transform 1 0 564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1712256841
transform 1 0 852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1712256841
transform 1 0 700 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1712256841
transform 1 0 692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1712256841
transform 1 0 692 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1712256841
transform 1 0 612 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1712256841
transform 1 0 564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1712256841
transform 1 0 2084 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1712256841
transform 1 0 1940 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1712256841
transform 1 0 2460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1712256841
transform 1 0 1932 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1712256841
transform 1 0 1956 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1712256841
transform 1 0 1924 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1712256841
transform 1 0 1892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1712256841
transform 1 0 1892 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1712256841
transform 1 0 1956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1712256841
transform 1 0 1884 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1712256841
transform 1 0 1900 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1712256841
transform 1 0 1436 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1712256841
transform 1 0 2252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1712256841
transform 1 0 2244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1712256841
transform 1 0 2244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1712256841
transform 1 0 2244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1712256841
transform 1 0 2220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1712256841
transform 1 0 2196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1712256841
transform 1 0 1828 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1712256841
transform 1 0 1780 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1712256841
transform 1 0 1764 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1712256841
transform 1 0 1716 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1712256841
transform 1 0 1620 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1712256841
transform 1 0 1428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1712256841
transform 1 0 1420 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1712256841
transform 1 0 1436 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1712256841
transform 1 0 1404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1712256841
transform 1 0 1484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1712256841
transform 1 0 1468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1712256841
transform 1 0 1396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1712256841
transform 1 0 1380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1712256841
transform 1 0 1276 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1712256841
transform 1 0 1220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1712256841
transform 1 0 1500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1712256841
transform 1 0 1412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1712256841
transform 1 0 1212 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1712256841
transform 1 0 1188 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1712256841
transform 1 0 1124 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1712256841
transform 1 0 1092 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1712256841
transform 1 0 1948 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1712256841
transform 1 0 1948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1712256841
transform 1 0 2228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1712256841
transform 1 0 1988 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1712256841
transform 1 0 2516 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1712256841
transform 1 0 2372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1712256841
transform 1 0 2188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1712256841
transform 1 0 2060 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1712256841
transform 1 0 1612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1712256841
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1712256841
transform 1 0 2308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1712256841
transform 1 0 2300 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1712256841
transform 1 0 2268 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1712256841
transform 1 0 2268 0 1 755
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1712256841
transform 1 0 2244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1712256841
transform 1 0 2188 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1712256841
transform 1 0 1932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1712256841
transform 1 0 1908 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1712256841
transform 1 0 1828 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1712256841
transform 1 0 2076 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1712256841
transform 1 0 1940 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1712256841
transform 1 0 1932 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1712256841
transform 1 0 1932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1712256841
transform 1 0 1900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1712256841
transform 1 0 1852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1712256841
transform 1 0 1956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1712256841
transform 1 0 1844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1712256841
transform 1 0 1732 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1712256841
transform 1 0 1716 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1712256841
transform 1 0 1708 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1712256841
transform 1 0 1620 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1712256841
transform 1 0 1588 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1712256841
transform 1 0 2612 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1712256841
transform 1 0 2460 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1712256841
transform 1 0 2428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1712256841
transform 1 0 2404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1712256841
transform 1 0 2452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1712256841
transform 1 0 2444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1712256841
transform 1 0 2372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1712256841
transform 1 0 2356 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1712256841
transform 1 0 2316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1712256841
transform 1 0 2284 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1712256841
transform 1 0 2676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1712256841
transform 1 0 2628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1712256841
transform 1 0 2524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1712256841
transform 1 0 2508 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1712256841
transform 1 0 2436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1712256841
transform 1 0 2412 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1712256841
transform 1 0 2092 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1712256841
transform 1 0 2084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1712256841
transform 1 0 3068 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1712256841
transform 1 0 3012 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1712256841
transform 1 0 2932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1712256841
transform 1 0 2916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1712256841
transform 1 0 2548 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1712256841
transform 1 0 2540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1712256841
transform 1 0 2276 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1712256841
transform 1 0 2236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1712256841
transform 1 0 2236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1712256841
transform 1 0 2220 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1712256841
transform 1 0 2220 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1712256841
transform 1 0 2188 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1712256841
transform 1 0 2092 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1712256841
transform 1 0 2044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1712256841
transform 1 0 2020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1712256841
transform 1 0 2060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1712256841
transform 1 0 1972 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1712256841
transform 1 0 1972 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1712256841
transform 1 0 1932 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1712256841
transform 1 0 1860 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1712256841
transform 1 0 1780 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1712256841
transform 1 0 1724 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1712256841
transform 1 0 2204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1712256841
transform 1 0 2092 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1712256841
transform 1 0 2076 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1712256841
transform 1 0 2060 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1712256841
transform 1 0 2036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1712256841
transform 1 0 2028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1712256841
transform 1 0 2012 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1712256841
transform 1 0 1716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1712256841
transform 1 0 1660 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1712256841
transform 1 0 1700 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1712256841
transform 1 0 1676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1712256841
transform 1 0 1636 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1712256841
transform 1 0 1612 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1712256841
transform 1 0 3244 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1712256841
transform 1 0 1908 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1712256841
transform 1 0 1604 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1712256841
transform 1 0 1596 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1712256841
transform 1 0 1596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1712256841
transform 1 0 1380 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1712256841
transform 1 0 1620 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1712256841
transform 1 0 1620 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1712256841
transform 1 0 1596 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1712256841
transform 1 0 1580 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1712256841
transform 1 0 1836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1712256841
transform 1 0 1604 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1712256841
transform 1 0 1548 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1712256841
transform 1 0 372 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1712256841
transform 1 0 1580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1712256841
transform 1 0 1436 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1712256841
transform 1 0 1468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1712256841
transform 1 0 1420 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1712256841
transform 1 0 1468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1712256841
transform 1 0 1420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1712256841
transform 1 0 1412 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1712256841
transform 1 0 1380 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1712256841
transform 1 0 772 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1712256841
transform 1 0 724 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1712256841
transform 1 0 724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1712256841
transform 1 0 724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1712256841
transform 1 0 540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1712256841
transform 1 0 420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1712256841
transform 1 0 484 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1712256841
transform 1 0 412 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1712256841
transform 1 0 412 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1712256841
transform 1 0 428 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1712256841
transform 1 0 356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1712256841
transform 1 0 1444 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1712256841
transform 1 0 1340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1712256841
transform 1 0 1284 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1712256841
transform 1 0 1284 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1712256841
transform 1 0 2044 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1712256841
transform 1 0 1996 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1712256841
transform 1 0 1532 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1712256841
transform 1 0 372 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1712256841
transform 1 0 348 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1712256841
transform 1 0 356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1712256841
transform 1 0 348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1712256841
transform 1 0 436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1712256841
transform 1 0 340 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1712256841
transform 1 0 404 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1712256841
transform 1 0 404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1712256841
transform 1 0 396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1712256841
transform 1 0 316 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1712256841
transform 1 0 316 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1712256841
transform 1 0 388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1712256841
transform 1 0 380 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1712256841
transform 1 0 428 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1712256841
transform 1 0 348 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1712256841
transform 1 0 348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1712256841
transform 1 0 468 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1712256841
transform 1 0 404 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1712256841
transform 1 0 356 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1712256841
transform 1 0 436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1712256841
transform 1 0 436 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1712256841
transform 1 0 332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1712256841
transform 1 0 364 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1712256841
transform 1 0 364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1712256841
transform 1 0 524 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1712256841
transform 1 0 340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1712256841
transform 1 0 340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1712256841
transform 1 0 420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1712256841
transform 1 0 340 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1712256841
transform 1 0 1876 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1712256841
transform 1 0 1860 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1712256841
transform 1 0 2684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1712256841
transform 1 0 1884 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1712256841
transform 1 0 2892 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1712256841
transform 1 0 2660 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1712256841
transform 1 0 2652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1712256841
transform 1 0 2644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1712256841
transform 1 0 2684 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1712256841
transform 1 0 2612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1712256841
transform 1 0 2588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1712256841
transform 1 0 2588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1712256841
transform 1 0 2228 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1712256841
transform 1 0 2628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1712256841
transform 1 0 2420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1712256841
transform 1 0 2268 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1712256841
transform 1 0 2644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1712256841
transform 1 0 2476 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1712256841
transform 1 0 2452 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1712256841
transform 1 0 1852 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1712256841
transform 1 0 1836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1712256841
transform 1 0 2148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1712256841
transform 1 0 1916 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1712256841
transform 1 0 2428 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1712256841
transform 1 0 2308 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1712256841
transform 1 0 2132 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1712256841
transform 1 0 2236 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1712256841
transform 1 0 2204 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1712256841
transform 1 0 2188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1712256841
transform 1 0 1948 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1712256841
transform 1 0 1908 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1712256841
transform 1 0 1820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1712256841
transform 1 0 1852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1712256841
transform 1 0 1788 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1712256841
transform 1 0 1732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1712256841
transform 1 0 2028 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1712256841
transform 1 0 1572 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1712256841
transform 1 0 1588 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1712256841
transform 1 0 1292 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1712256841
transform 1 0 1268 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1712256841
transform 1 0 1260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1712256841
transform 1 0 1260 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1712256841
transform 1 0 1244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1712256841
transform 1 0 1276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1712256841
transform 1 0 1108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1712256841
transform 1 0 1124 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1712256841
transform 1 0 940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1712256841
transform 1 0 940 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1712256841
transform 1 0 2492 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1712256841
transform 1 0 2060 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1712256841
transform 1 0 2476 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1712256841
transform 1 0 2476 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1712256841
transform 1 0 2476 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1712256841
transform 1 0 2508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1712256841
transform 1 0 2212 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1712256841
transform 1 0 2132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1712256841
transform 1 0 1900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1712256841
transform 1 0 1860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1712256841
transform 1 0 1804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1712256841
transform 1 0 1700 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1712256841
transform 1 0 1364 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1712256841
transform 1 0 204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1712256841
transform 1 0 1364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1712256841
transform 1 0 684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1712256841
transform 1 0 1628 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1712256841
transform 1 0 1372 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1712256841
transform 1 0 1988 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1712256841
transform 1 0 1660 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1712256841
transform 1 0 1676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1712256841
transform 1 0 1676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1712256841
transform 1 0 2172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1712256841
transform 1 0 1644 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1712256841
transform 1 0 1668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1712256841
transform 1 0 1660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1712256841
transform 1 0 1660 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1712256841
transform 1 0 1620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1712256841
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1712256841
transform 1 0 1724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1712256841
transform 1 0 1604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1712256841
transform 1 0 1644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1712256841
transform 1 0 1516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1712256841
transform 1 0 1492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1712256841
transform 1 0 1204 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1712256841
transform 1 0 1148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1712256841
transform 1 0 1100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1712256841
transform 1 0 2140 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1712256841
transform 1 0 2116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1712256841
transform 1 0 2012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1712256841
transform 1 0 2220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1712256841
transform 1 0 2196 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1712256841
transform 1 0 2244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1712256841
transform 1 0 2204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1712256841
transform 1 0 2204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1712256841
transform 1 0 2228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1712256841
transform 1 0 2228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1712256841
transform 1 0 2148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1712256841
transform 1 0 2028 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1712256841
transform 1 0 1972 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1712256841
transform 1 0 2244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1712256841
transform 1 0 1972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1712256841
transform 1 0 1980 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1712256841
transform 1 0 1980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1712256841
transform 1 0 2108 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1712256841
transform 1 0 2060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1712256841
transform 1 0 2052 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1712256841
transform 1 0 2052 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1712256841
transform 1 0 1964 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1712256841
transform 1 0 2012 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1712256841
transform 1 0 2004 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1712256841
transform 1 0 2156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1712256841
transform 1 0 1988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1712256841
transform 1 0 1988 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1712256841
transform 1 0 2020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1712256841
transform 1 0 1820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1712256841
transform 1 0 1820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1712256841
transform 1 0 2484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1712256841
transform 1 0 2196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1712256841
transform 1 0 2068 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1712256841
transform 1 0 2332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1712256841
transform 1 0 2284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1712256841
transform 1 0 2172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1712256841
transform 1 0 2116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1712256841
transform 1 0 2020 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1712256841
transform 1 0 2036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1712256841
transform 1 0 1892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1712256841
transform 1 0 668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1712256841
transform 1 0 652 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1712256841
transform 1 0 668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1712256841
transform 1 0 316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1712256841
transform 1 0 260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1712256841
transform 1 0 116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1712256841
transform 1 0 100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1712256841
transform 1 0 284 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1712256841
transform 1 0 220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1712256841
transform 1 0 228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1712256841
transform 1 0 164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1712256841
transform 1 0 116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1712256841
transform 1 0 708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1712256841
transform 1 0 684 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1712256841
transform 1 0 836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1712256841
transform 1 0 812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1712256841
transform 1 0 700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1712256841
transform 1 0 724 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1712256841
transform 1 0 524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1712256841
transform 1 0 524 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1712256841
transform 1 0 540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1712256841
transform 1 0 196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1712256841
transform 1 0 172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1712256841
transform 1 0 164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1712256841
transform 1 0 260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1712256841
transform 1 0 116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1712256841
transform 1 0 1140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1712256841
transform 1 0 132 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1712256841
transform 1 0 84 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1712256841
transform 1 0 276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1712256841
transform 1 0 260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1712256841
transform 1 0 252 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1712256841
transform 1 0 604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1712256841
transform 1 0 476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1712256841
transform 1 0 268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1712256841
transform 1 0 148 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1712256841
transform 1 0 108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1712256841
transform 1 0 148 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1712256841
transform 1 0 100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1712256841
transform 1 0 132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1712256841
transform 1 0 132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1712256841
transform 1 0 116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1712256841
transform 1 0 116 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1712256841
transform 1 0 108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1712256841
transform 1 0 84 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1712256841
transform 1 0 1796 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1712256841
transform 1 0 1668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1712256841
transform 1 0 1652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1712256841
transform 1 0 1436 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1712256841
transform 1 0 3156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1712256841
transform 1 0 1724 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1712256841
transform 1 0 1708 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1712256841
transform 1 0 1700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1712256841
transform 1 0 1452 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1712256841
transform 1 0 1388 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1712256841
transform 1 0 1372 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1712256841
transform 1 0 820 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1712256841
transform 1 0 1420 0 1 1445
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1712256841
transform 1 0 1420 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1712256841
transform 1 0 1404 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1712256841
transform 1 0 364 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1712256841
transform 1 0 340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1712256841
transform 1 0 332 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1712256841
transform 1 0 380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1712256841
transform 1 0 348 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1712256841
transform 1 0 1052 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1712256841
transform 1 0 1052 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1712256841
transform 1 0 1036 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1712256841
transform 1 0 1036 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1712256841
transform 1 0 492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1712256841
transform 1 0 300 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1712256841
transform 1 0 300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1712256841
transform 1 0 411 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1712256841
transform 1 0 348 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1712256841
transform 1 0 348 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1712256841
transform 1 0 292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1712256841
transform 1 0 428 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1712256841
transform 1 0 308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1712256841
transform 1 0 308 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1712256841
transform 1 0 1660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1712256841
transform 1 0 1500 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1712256841
transform 1 0 1428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1712256841
transform 1 0 796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1712256841
transform 1 0 556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1712256841
transform 1 0 1964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1712256841
transform 1 0 1732 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1712256841
transform 1 0 1716 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1712256841
transform 1 0 564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1712256841
transform 1 0 548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1712256841
transform 1 0 276 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1712256841
transform 1 0 276 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1712256841
transform 1 0 220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1712256841
transform 1 0 364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1712256841
transform 1 0 332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1712256841
transform 1 0 356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1712256841
transform 1 0 300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1712256841
transform 1 0 380 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1712256841
transform 1 0 348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1712256841
transform 1 0 284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1712256841
transform 1 0 316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1712256841
transform 1 0 316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1712256841
transform 1 0 260 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1712256841
transform 1 0 260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1712256841
transform 1 0 2148 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1712256841
transform 1 0 2108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1712256841
transform 1 0 2100 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1712256841
transform 1 0 748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1712256841
transform 1 0 724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1712256841
transform 1 0 2076 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1712256841
transform 1 0 2076 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1712256841
transform 1 0 2036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1712256841
transform 1 0 860 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1712256841
transform 1 0 828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1712256841
transform 1 0 308 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1712256841
transform 1 0 276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1712256841
transform 1 0 380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1712256841
transform 1 0 252 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1712256841
transform 1 0 212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1712256841
transform 1 0 2116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1712256841
transform 1 0 2108 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1712256841
transform 1 0 2036 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1712256841
transform 1 0 572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1712256841
transform 1 0 540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1712256841
transform 1 0 532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1712256841
transform 1 0 852 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1712256841
transform 1 0 756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1712256841
transform 1 0 588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1712256841
transform 1 0 444 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1712256841
transform 1 0 428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1712256841
transform 1 0 388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1712256841
transform 1 0 388 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1712256841
transform 1 0 388 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1712256841
transform 1 0 436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1712256841
transform 1 0 260 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1712256841
transform 1 0 228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1712256841
transform 1 0 1020 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1712256841
transform 1 0 932 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3699
timestamp 1712256841
transform 1 0 828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1712256841
transform 1 0 572 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1712256841
transform 1 0 508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3702
timestamp 1712256841
transform 1 0 500 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1712256841
transform 1 0 484 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1712256841
transform 1 0 484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1712256841
transform 1 0 780 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1712256841
transform 1 0 676 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3707
timestamp 1712256841
transform 1 0 556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3708
timestamp 1712256841
transform 1 0 516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1712256841
transform 1 0 508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1712256841
transform 1 0 772 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1712256841
transform 1 0 748 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1712256841
transform 1 0 668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1712256841
transform 1 0 636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1712256841
transform 1 0 564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1712256841
transform 1 0 564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1712256841
transform 1 0 1476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1712256841
transform 1 0 1436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1712256841
transform 1 0 1988 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1712256841
transform 1 0 1620 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1712256841
transform 1 0 1460 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1712256841
transform 1 0 1484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1712256841
transform 1 0 1380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1712256841
transform 1 0 1340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1712256841
transform 1 0 884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1712256841
transform 1 0 836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1712256841
transform 1 0 644 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1712256841
transform 1 0 140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1712256841
transform 1 0 116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1712256841
transform 1 0 1476 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1712256841
transform 1 0 1452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1712256841
transform 1 0 1628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1712256841
transform 1 0 1532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1712256841
transform 1 0 1428 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1712256841
transform 1 0 1460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1712256841
transform 1 0 1444 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1712256841
transform 1 0 1364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1712256841
transform 1 0 1388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1712256841
transform 1 0 1372 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1712256841
transform 1 0 2332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1712256841
transform 1 0 1780 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1712256841
transform 1 0 1804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1712256841
transform 1 0 1780 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1712256841
transform 1 0 1836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1712256841
transform 1 0 1788 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1712256841
transform 1 0 1972 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1712256841
transform 1 0 1828 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1712256841
transform 1 0 1860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1712256841
transform 1 0 1396 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1712256841
transform 1 0 1364 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1712256841
transform 1 0 1332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1712256841
transform 1 0 1468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1712256841
transform 1 0 1412 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3753
timestamp 1712256841
transform 1 0 1308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1712256841
transform 1 0 1348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1712256841
transform 1 0 1220 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1712256841
transform 1 0 1220 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1712256841
transform 1 0 1828 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1712256841
transform 1 0 1796 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1712256841
transform 1 0 1732 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1712256841
transform 1 0 1540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1712256841
transform 1 0 1300 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1712256841
transform 1 0 1300 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1712256841
transform 1 0 1004 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1712256841
transform 1 0 1004 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1712256841
transform 1 0 2412 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3766
timestamp 1712256841
transform 1 0 1988 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1712256841
transform 1 0 2396 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1712256841
transform 1 0 2364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1712256841
transform 1 0 2364 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1712256841
transform 1 0 2436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1712256841
transform 1 0 2340 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1712256841
transform 1 0 2308 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1712256841
transform 1 0 2436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1712256841
transform 1 0 2396 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1712256841
transform 1 0 2364 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1712256841
transform 1 0 2356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1712256841
transform 1 0 2028 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1712256841
transform 1 0 2564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1712256841
transform 1 0 2540 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1712256841
transform 1 0 2524 0 1 1895
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1712256841
transform 1 0 2524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1712256841
transform 1 0 1852 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1712256841
transform 1 0 1788 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1712256841
transform 1 0 1756 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3785
timestamp 1712256841
transform 1 0 2276 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1712256841
transform 1 0 1772 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1712256841
transform 1 0 1820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1712256841
transform 1 0 1788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1712256841
transform 1 0 1908 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1712256841
transform 1 0 1844 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1712256841
transform 1 0 1804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1712256841
transform 1 0 2020 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1712256841
transform 1 0 1892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1712256841
transform 1 0 1844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1712256841
transform 1 0 2884 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1712256841
transform 1 0 2884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1712256841
transform 1 0 2852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1712256841
transform 1 0 2556 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1712256841
transform 1 0 2540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1712256841
transform 1 0 2524 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1712256841
transform 1 0 2500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1712256841
transform 1 0 2020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1712256841
transform 1 0 1972 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1712256841
transform 1 0 1972 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1712256841
transform 1 0 3084 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1712256841
transform 1 0 3036 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1712256841
transform 1 0 3020 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3808
timestamp 1712256841
transform 1 0 2572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1712256841
transform 1 0 2572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1712256841
transform 1 0 2772 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1712256841
transform 1 0 2044 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1712256841
transform 1 0 1852 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1712256841
transform 1 0 2300 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1712256841
transform 1 0 2244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1712256841
transform 1 0 2236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1712256841
transform 1 0 2484 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1712256841
transform 1 0 2428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1712256841
transform 1 0 2308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1712256841
transform 1 0 3068 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1712256841
transform 1 0 3068 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1712256841
transform 1 0 2796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1712256841
transform 1 0 2612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1712256841
transform 1 0 2604 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1712256841
transform 1 0 2508 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1712256841
transform 1 0 2412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3826
timestamp 1712256841
transform 1 0 2396 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1712256841
transform 1 0 2372 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1712256841
transform 1 0 2308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1712256841
transform 1 0 2404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1712256841
transform 1 0 2380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1712256841
transform 1 0 2364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1712256841
transform 1 0 2260 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1712256841
transform 1 0 2228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1712256841
transform 1 0 2412 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1712256841
transform 1 0 2284 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1712256841
transform 1 0 2180 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1712256841
transform 1 0 2836 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1712256841
transform 1 0 2764 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1712256841
transform 1 0 2700 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1712256841
transform 1 0 3140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1712256841
transform 1 0 3004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1712256841
transform 1 0 2988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1712256841
transform 1 0 1796 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1712256841
transform 1 0 1692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1712256841
transform 1 0 1700 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1712256841
transform 1 0 204 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1712256841
transform 1 0 140 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1712256841
transform 1 0 108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1712256841
transform 1 0 156 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1712256841
transform 1 0 108 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1712256841
transform 1 0 684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1712256841
transform 1 0 92 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1712256841
transform 1 0 116 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1712256841
transform 1 0 116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1712256841
transform 1 0 140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1712256841
transform 1 0 132 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1712256841
transform 1 0 84 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1712256841
transform 1 0 2196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1712256841
transform 1 0 2156 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1712256841
transform 1 0 1716 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1712256841
transform 1 0 1292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1712256841
transform 1 0 1292 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1712256841
transform 1 0 708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1712256841
transform 1 0 524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1712256841
transform 1 0 396 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1712256841
transform 1 0 380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1712256841
transform 1 0 324 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1712256841
transform 1 0 100 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1712256841
transform 1 0 164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1712256841
transform 1 0 140 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1712256841
transform 1 0 124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1712256841
transform 1 0 124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1712256841
transform 1 0 124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1712256841
transform 1 0 172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1712256841
transform 1 0 164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1712256841
transform 1 0 92 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1712256841
transform 1 0 740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1712256841
transform 1 0 724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1712256841
transform 1 0 1092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1712256841
transform 1 0 1012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1712256841
transform 1 0 732 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1712256841
transform 1 0 804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1712256841
transform 1 0 804 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1712256841
transform 1 0 540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1712256841
transform 1 0 508 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1712256841
transform 1 0 164 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1712256841
transform 1 0 84 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1712256841
transform 1 0 84 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1712256841
transform 1 0 84 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1712256841
transform 1 0 84 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1712256841
transform 1 0 156 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1712256841
transform 1 0 84 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1712256841
transform 1 0 172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1712256841
transform 1 0 116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1712256841
transform 1 0 100 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1712256841
transform 1 0 172 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1712256841
transform 1 0 172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1712256841
transform 1 0 84 0 1 1095
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1712256841
transform 1 0 196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1712256841
transform 1 0 92 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1712256841
transform 1 0 516 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1712256841
transform 1 0 180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1712256841
transform 1 0 180 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3904
timestamp 1712256841
transform 1 0 212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1712256841
transform 1 0 212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1712256841
transform 1 0 100 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1712256841
transform 1 0 1116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1712256841
transform 1 0 1116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1712256841
transform 1 0 1220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3910
timestamp 1712256841
transform 1 0 1124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1712256841
transform 1 0 1380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1712256841
transform 1 0 1340 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1712256841
transform 1 0 1196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1712256841
transform 1 0 1188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1712256841
transform 1 0 1244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3916
timestamp 1712256841
transform 1 0 1244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1712256841
transform 1 0 1356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1712256841
transform 1 0 1332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1712256841
transform 1 0 1260 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1712256841
transform 1 0 1212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1712256841
transform 1 0 1436 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1712256841
transform 1 0 1340 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_3923
timestamp 1712256841
transform 1 0 1188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1712256841
transform 1 0 1108 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3925
timestamp 1712256841
transform 1 0 1620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3926
timestamp 1712256841
transform 1 0 1508 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1712256841
transform 1 0 1308 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3928
timestamp 1712256841
transform 1 0 1124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1712256841
transform 1 0 1956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1712256841
transform 1 0 1772 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1712256841
transform 1 0 1772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1712256841
transform 1 0 1764 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1712256841
transform 1 0 1812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3934
timestamp 1712256841
transform 1 0 1756 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3935
timestamp 1712256841
transform 1 0 2108 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1712256841
transform 1 0 1860 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3937
timestamp 1712256841
transform 1 0 1900 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1712256841
transform 1 0 1876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3939
timestamp 1712256841
transform 1 0 1852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1712256841
transform 1 0 1532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1712256841
transform 1 0 1356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3942
timestamp 1712256841
transform 1 0 2476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3943
timestamp 1712256841
transform 1 0 2428 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1712256841
transform 1 0 2364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1712256841
transform 1 0 2332 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3946
timestamp 1712256841
transform 1 0 2044 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3947
timestamp 1712256841
transform 1 0 2028 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1712256841
transform 1 0 1948 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1712256841
transform 1 0 1932 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1712256841
transform 1 0 1892 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1712256841
transform 1 0 1892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3952
timestamp 1712256841
transform 1 0 1884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1712256841
transform 1 0 1924 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1712256841
transform 1 0 1916 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1712256841
transform 1 0 2100 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1712256841
transform 1 0 2020 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1712256841
transform 1 0 1948 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1712256841
transform 1 0 1916 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1712256841
transform 1 0 1932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1712256841
transform 1 0 1732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3961
timestamp 1712256841
transform 1 0 2932 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1712256841
transform 1 0 2612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1712256841
transform 1 0 2540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3964
timestamp 1712256841
transform 1 0 2508 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3965
timestamp 1712256841
transform 1 0 2468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1712256841
transform 1 0 2188 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3967
timestamp 1712256841
transform 1 0 2132 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1712256841
transform 1 0 2092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1712256841
transform 1 0 2060 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1712256841
transform 1 0 1996 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1712256841
transform 1 0 1980 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1712256841
transform 1 0 1980 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1712256841
transform 1 0 1980 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_3974
timestamp 1712256841
transform 1 0 2156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3975
timestamp 1712256841
transform 1 0 2132 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1712256841
transform 1 0 2148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1712256841
transform 1 0 2148 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1712256841
transform 1 0 2076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1712256841
transform 1 0 2076 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3980
timestamp 1712256841
transform 1 0 2196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1712256841
transform 1 0 2164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3982
timestamp 1712256841
transform 1 0 2164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1712256841
transform 1 0 2164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1712256841
transform 1 0 2084 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1712256841
transform 1 0 1700 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1712256841
transform 1 0 1596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3987
timestamp 1712256841
transform 1 0 2228 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1712256841
transform 1 0 1724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1712256841
transform 1 0 2148 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1712256841
transform 1 0 2148 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1712256841
transform 1 0 2300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1712256841
transform 1 0 2300 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1712256841
transform 1 0 1996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1712256841
transform 1 0 1676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3995
timestamp 1712256841
transform 1 0 1580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1712256841
transform 1 0 1628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1712256841
transform 1 0 1076 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1712256841
transform 1 0 652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1712256841
transform 1 0 2108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1712256841
transform 1 0 2108 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1712256841
transform 1 0 2044 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1712256841
transform 1 0 1940 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1712256841
transform 1 0 1900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1712256841
transform 1 0 1892 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1712256841
transform 1 0 1852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4006
timestamp 1712256841
transform 1 0 1804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1712256841
transform 1 0 1788 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1712256841
transform 1 0 1916 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1712256841
transform 1 0 1836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4010
timestamp 1712256841
transform 1 0 1820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1712256841
transform 1 0 1572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4012
timestamp 1712256841
transform 1 0 1356 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1712256841
transform 1 0 1612 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1712256841
transform 1 0 1540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1712256841
transform 1 0 1492 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1712256841
transform 1 0 1460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1712256841
transform 1 0 1516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1712256841
transform 1 0 1460 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1712256841
transform 1 0 1324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1712256841
transform 1 0 1324 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1712256841
transform 1 0 1308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4022
timestamp 1712256841
transform 1 0 1300 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1712256841
transform 1 0 1300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1712256841
transform 1 0 852 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1712256841
transform 1 0 836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1712256841
transform 1 0 812 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1712256841
transform 1 0 532 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4028
timestamp 1712256841
transform 1 0 500 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4029
timestamp 1712256841
transform 1 0 484 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1712256841
transform 1 0 468 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1712256841
transform 1 0 468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1712256841
transform 1 0 1340 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1712256841
transform 1 0 1308 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1712256841
transform 1 0 1284 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1712256841
transform 1 0 1260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1712256841
transform 1 0 1620 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_4037
timestamp 1712256841
transform 1 0 1612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1712256841
transform 1 0 3156 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4039
timestamp 1712256841
transform 1 0 1596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4040
timestamp 1712256841
transform 1 0 1580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4041
timestamp 1712256841
transform 1 0 1412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1712256841
transform 1 0 1356 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1712256841
transform 1 0 1732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1712256841
transform 1 0 1716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1712256841
transform 1 0 1660 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1712256841
transform 1 0 1292 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1712256841
transform 1 0 1252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1712256841
transform 1 0 1236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1712256841
transform 1 0 1228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1712256841
transform 1 0 1164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1712256841
transform 1 0 1164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1712256841
transform 1 0 1268 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4053
timestamp 1712256841
transform 1 0 1220 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1712256841
transform 1 0 1148 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1712256841
transform 1 0 828 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4056
timestamp 1712256841
transform 1 0 1428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1712256841
transform 1 0 1372 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1712256841
transform 1 0 1204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1712256841
transform 1 0 1228 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1712256841
transform 1 0 1188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1712256841
transform 1 0 1156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1712256841
transform 1 0 1068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1712256841
transform 1 0 748 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1712256841
transform 1 0 500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1712256841
transform 1 0 1276 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1712256841
transform 1 0 1116 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1712256841
transform 1 0 1372 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1712256841
transform 1 0 1244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4069
timestamp 1712256841
transform 1 0 1228 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1712256841
transform 1 0 1228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1712256841
transform 1 0 1084 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1712256841
transform 1 0 1044 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1712256841
transform 1 0 924 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1712256841
transform 1 0 636 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1712256841
transform 1 0 348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1712256841
transform 1 0 300 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4077
timestamp 1712256841
transform 1 0 284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4078
timestamp 1712256841
transform 1 0 1188 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4079
timestamp 1712256841
transform 1 0 1060 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1712256841
transform 1 0 1036 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1712256841
transform 1 0 1012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4082
timestamp 1712256841
transform 1 0 1428 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1712256841
transform 1 0 1428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4084
timestamp 1712256841
transform 1 0 956 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4085
timestamp 1712256841
transform 1 0 948 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1712256841
transform 1 0 916 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4087
timestamp 1712256841
transform 1 0 900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1712256841
transform 1 0 812 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1712256841
transform 1 0 1124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4090
timestamp 1712256841
transform 1 0 820 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1712256841
transform 1 0 1340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1712256841
transform 1 0 1084 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4093
timestamp 1712256841
transform 1 0 1156 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4094
timestamp 1712256841
transform 1 0 1092 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1712256841
transform 1 0 1156 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1712256841
transform 1 0 1148 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1712256841
transform 1 0 1092 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1712256841
transform 1 0 1084 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1712256841
transform 1 0 980 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1712256841
transform 1 0 660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1712256841
transform 1 0 380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4102
timestamp 1712256841
transform 1 0 316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1712256841
transform 1 0 244 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1712256841
transform 1 0 1188 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1712256841
transform 1 0 1140 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4106
timestamp 1712256841
transform 1 0 1124 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1712256841
transform 1 0 1100 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1712256841
transform 1 0 1100 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1712256841
transform 1 0 1372 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1712256841
transform 1 0 1340 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1712256841
transform 1 0 3164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4112
timestamp 1712256841
transform 1 0 3132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1712256841
transform 1 0 3044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1712256841
transform 1 0 2996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1712256841
transform 1 0 2972 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1712256841
transform 1 0 1028 0 1 2285
box -2 -2 2 2
use M2_M1  M2_M1_4117
timestamp 1712256841
transform 1 0 764 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1712256841
transform 1 0 1356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1712256841
transform 1 0 988 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4120
timestamp 1712256841
transform 1 0 1004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1712256841
transform 1 0 1004 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1712256841
transform 1 0 1028 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1712256841
transform 1 0 996 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4124
timestamp 1712256841
transform 1 0 1012 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4125
timestamp 1712256841
transform 1 0 940 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4126
timestamp 1712256841
transform 1 0 1380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1712256841
transform 1 0 1340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4128
timestamp 1712256841
transform 1 0 1140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4129
timestamp 1712256841
transform 1 0 1060 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1712256841
transform 1 0 1036 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4131
timestamp 1712256841
transform 1 0 1036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4132
timestamp 1712256841
transform 1 0 1036 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4133
timestamp 1712256841
transform 1 0 892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4134
timestamp 1712256841
transform 1 0 1292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1712256841
transform 1 0 1188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1712256841
transform 1 0 1212 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4137
timestamp 1712256841
transform 1 0 1148 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4138
timestamp 1712256841
transform 1 0 2884 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4139
timestamp 1712256841
transform 1 0 2724 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4140
timestamp 1712256841
transform 1 0 2228 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1712256841
transform 1 0 1468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1712256841
transform 1 0 1372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4143
timestamp 1712256841
transform 1 0 1348 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4144
timestamp 1712256841
transform 1 0 1332 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4145
timestamp 1712256841
transform 1 0 1300 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4146
timestamp 1712256841
transform 1 0 1268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4147
timestamp 1712256841
transform 1 0 2828 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4148
timestamp 1712256841
transform 1 0 2828 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1712256841
transform 1 0 1716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4150
timestamp 1712256841
transform 1 0 1348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4151
timestamp 1712256841
transform 1 0 1348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4152
timestamp 1712256841
transform 1 0 1348 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1712256841
transform 1 0 1332 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4154
timestamp 1712256841
transform 1 0 1260 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4155
timestamp 1712256841
transform 1 0 1348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4156
timestamp 1712256841
transform 1 0 1316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4157
timestamp 1712256841
transform 1 0 1372 0 1 1895
box -2 -2 2 2
use M2_M1  M2_M1_4158
timestamp 1712256841
transform 1 0 1372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4159
timestamp 1712256841
transform 1 0 1476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4160
timestamp 1712256841
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4161
timestamp 1712256841
transform 1 0 1412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1712256841
transform 1 0 1332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4163
timestamp 1712256841
transform 1 0 1300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4164
timestamp 1712256841
transform 1 0 1132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4165
timestamp 1712256841
transform 1 0 1044 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4166
timestamp 1712256841
transform 1 0 1004 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4167
timestamp 1712256841
transform 1 0 996 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4168
timestamp 1712256841
transform 1 0 956 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4169
timestamp 1712256841
transform 1 0 1580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4170
timestamp 1712256841
transform 1 0 1484 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4171
timestamp 1712256841
transform 1 0 564 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4172
timestamp 1712256841
transform 1 0 524 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4173
timestamp 1712256841
transform 1 0 532 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1712256841
transform 1 0 532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4175
timestamp 1712256841
transform 1 0 764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4176
timestamp 1712256841
transform 1 0 540 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4177
timestamp 1712256841
transform 1 0 956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4178
timestamp 1712256841
transform 1 0 788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4179
timestamp 1712256841
transform 1 0 804 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4180
timestamp 1712256841
transform 1 0 740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4181
timestamp 1712256841
transform 1 0 1148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4182
timestamp 1712256841
transform 1 0 1092 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4183
timestamp 1712256841
transform 1 0 924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4184
timestamp 1712256841
transform 1 0 828 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4185
timestamp 1712256841
transform 1 0 780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4186
timestamp 1712256841
transform 1 0 764 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4187
timestamp 1712256841
transform 1 0 764 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4188
timestamp 1712256841
transform 1 0 316 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4189
timestamp 1712256841
transform 1 0 308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4190
timestamp 1712256841
transform 1 0 284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4191
timestamp 1712256841
transform 1 0 908 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4192
timestamp 1712256841
transform 1 0 804 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4193
timestamp 1712256841
transform 1 0 788 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1712256841
transform 1 0 1228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4195
timestamp 1712256841
transform 1 0 1084 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4196
timestamp 1712256841
transform 1 0 1140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1712256841
transform 1 0 1100 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1712256841
transform 1 0 1596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4199
timestamp 1712256841
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1712256841
transform 1 0 1276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1712256841
transform 1 0 1196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4202
timestamp 1712256841
transform 1 0 868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4203
timestamp 1712256841
transform 1 0 1220 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4204
timestamp 1712256841
transform 1 0 1188 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4205
timestamp 1712256841
transform 1 0 2772 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1712256841
transform 1 0 2772 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4207
timestamp 1712256841
transform 1 0 2580 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4208
timestamp 1712256841
transform 1 0 1636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4209
timestamp 1712256841
transform 1 0 1628 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4210
timestamp 1712256841
transform 1 0 1292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4211
timestamp 1712256841
transform 1 0 1260 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4212
timestamp 1712256841
transform 1 0 1044 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4213
timestamp 1712256841
transform 1 0 596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1712256841
transform 1 0 516 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4215
timestamp 1712256841
transform 1 0 596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4216
timestamp 1712256841
transform 1 0 572 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4217
timestamp 1712256841
transform 1 0 2924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1712256841
transform 1 0 2492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4219
timestamp 1712256841
transform 1 0 1172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4220
timestamp 1712256841
transform 1 0 884 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4221
timestamp 1712256841
transform 1 0 772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1712256841
transform 1 0 1124 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1712256841
transform 1 0 1124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4224
timestamp 1712256841
transform 1 0 844 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4225
timestamp 1712256841
transform 1 0 1556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4226
timestamp 1712256841
transform 1 0 1548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1712256841
transform 1 0 1100 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1712256841
transform 1 0 948 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4229
timestamp 1712256841
transform 1 0 1220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1712256841
transform 1 0 1108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4231
timestamp 1712256841
transform 1 0 420 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1712256841
transform 1 0 412 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4233
timestamp 1712256841
transform 1 0 388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1712256841
transform 1 0 372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1712256841
transform 1 0 572 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4236
timestamp 1712256841
transform 1 0 420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1712256841
transform 1 0 436 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1712256841
transform 1 0 436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4239
timestamp 1712256841
transform 1 0 1276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4240
timestamp 1712256841
transform 1 0 636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4241
timestamp 1712256841
transform 1 0 636 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4242
timestamp 1712256841
transform 1 0 572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4243
timestamp 1712256841
transform 1 0 500 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4244
timestamp 1712256841
transform 1 0 444 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4245
timestamp 1712256841
transform 1 0 348 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4246
timestamp 1712256841
transform 1 0 332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4247
timestamp 1712256841
transform 1 0 300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1712256841
transform 1 0 716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1712256841
transform 1 0 548 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1712256841
transform 1 0 548 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4251
timestamp 1712256841
transform 1 0 676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4252
timestamp 1712256841
transform 1 0 460 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1712256841
transform 1 0 460 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4254
timestamp 1712256841
transform 1 0 340 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4255
timestamp 1712256841
transform 1 0 340 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4256
timestamp 1712256841
transform 1 0 804 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4257
timestamp 1712256841
transform 1 0 628 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4258
timestamp 1712256841
transform 1 0 676 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4259
timestamp 1712256841
transform 1 0 644 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1712256841
transform 1 0 308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4261
timestamp 1712256841
transform 1 0 204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1712256841
transform 1 0 1884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1712256841
transform 1 0 1204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4264
timestamp 1712256841
transform 1 0 780 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4265
timestamp 1712256841
transform 1 0 764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4266
timestamp 1712256841
transform 1 0 2852 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4267
timestamp 1712256841
transform 1 0 2772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4268
timestamp 1712256841
transform 1 0 1852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1712256841
transform 1 0 1780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4270
timestamp 1712256841
transform 1 0 1468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4271
timestamp 1712256841
transform 1 0 972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4272
timestamp 1712256841
transform 1 0 908 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4273
timestamp 1712256841
transform 1 0 276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4274
timestamp 1712256841
transform 1 0 252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1712256841
transform 1 0 364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4276
timestamp 1712256841
transform 1 0 364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1712256841
transform 1 0 2860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4278
timestamp 1712256841
transform 1 0 2316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4279
timestamp 1712256841
transform 1 0 1276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1712256841
transform 1 0 692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4281
timestamp 1712256841
transform 1 0 676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4282
timestamp 1712256841
transform 1 0 1972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1712256841
transform 1 0 1364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4284
timestamp 1712256841
transform 1 0 628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4285
timestamp 1712256841
transform 1 0 596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1712256841
transform 1 0 1052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4287
timestamp 1712256841
transform 1 0 1052 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_4288
timestamp 1712256841
transform 1 0 1020 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_4289
timestamp 1712256841
transform 1 0 1020 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4290
timestamp 1712256841
transform 1 0 940 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4291
timestamp 1712256841
transform 1 0 868 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4292
timestamp 1712256841
transform 1 0 764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1712256841
transform 1 0 716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4294
timestamp 1712256841
transform 1 0 2764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1712256841
transform 1 0 1300 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1712256841
transform 1 0 1268 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4297
timestamp 1712256841
transform 1 0 1268 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4298
timestamp 1712256841
transform 1 0 1236 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4299
timestamp 1712256841
transform 1 0 1236 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1712256841
transform 1 0 1220 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4301
timestamp 1712256841
transform 1 0 1212 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1712256841
transform 1 0 1204 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4303
timestamp 1712256841
transform 1 0 1188 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1712256841
transform 1 0 1116 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1712256841
transform 1 0 1100 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1712256841
transform 1 0 364 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4307
timestamp 1712256841
transform 1 0 292 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1712256841
transform 1 0 220 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4309
timestamp 1712256841
transform 1 0 196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4310
timestamp 1712256841
transform 1 0 268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1712256841
transform 1 0 236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4312
timestamp 1712256841
transform 1 0 564 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1712256841
transform 1 0 300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1712256841
transform 1 0 364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1712256841
transform 1 0 332 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4316
timestamp 1712256841
transform 1 0 740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1712256841
transform 1 0 340 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4318
timestamp 1712256841
transform 1 0 324 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4319
timestamp 1712256841
transform 1 0 844 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4320
timestamp 1712256841
transform 1 0 300 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1712256841
transform 1 0 268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4322
timestamp 1712256841
transform 1 0 252 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4323
timestamp 1712256841
transform 1 0 220 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4324
timestamp 1712256841
transform 1 0 212 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4325
timestamp 1712256841
transform 1 0 148 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4326
timestamp 1712256841
transform 1 0 996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4327
timestamp 1712256841
transform 1 0 596 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4328
timestamp 1712256841
transform 1 0 588 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1712256841
transform 1 0 572 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1712256841
transform 1 0 180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4331
timestamp 1712256841
transform 1 0 132 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1712256841
transform 1 0 108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1712256841
transform 1 0 1932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4334
timestamp 1712256841
transform 1 0 1492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1712256841
transform 1 0 972 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1712256841
transform 1 0 956 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1712256841
transform 1 0 1028 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4338
timestamp 1712256841
transform 1 0 1004 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1712256841
transform 1 0 148 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1712256841
transform 1 0 108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4341
timestamp 1712256841
transform 1 0 188 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4342
timestamp 1712256841
transform 1 0 188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4343
timestamp 1712256841
transform 1 0 2772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4344
timestamp 1712256841
transform 1 0 2340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4345
timestamp 1712256841
transform 1 0 1564 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4346
timestamp 1712256841
transform 1 0 892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4347
timestamp 1712256841
transform 1 0 708 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4348
timestamp 1712256841
transform 1 0 2028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4349
timestamp 1712256841
transform 1 0 1732 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1712256841
transform 1 0 828 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4351
timestamp 1712256841
transform 1 0 828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4352
timestamp 1712256841
transform 1 0 1124 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4353
timestamp 1712256841
transform 1 0 1060 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1712256841
transform 1 0 964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4355
timestamp 1712256841
transform 1 0 900 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4356
timestamp 1712256841
transform 1 0 628 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_4357
timestamp 1712256841
transform 1 0 612 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4358
timestamp 1712256841
transform 1 0 284 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4359
timestamp 1712256841
transform 1 0 276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4360
timestamp 1712256841
transform 1 0 212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4361
timestamp 1712256841
transform 1 0 212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4362
timestamp 1712256841
transform 1 0 428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4363
timestamp 1712256841
transform 1 0 228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4364
timestamp 1712256841
transform 1 0 572 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4365
timestamp 1712256841
transform 1 0 388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4366
timestamp 1712256841
transform 1 0 436 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_4367
timestamp 1712256841
transform 1 0 436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4368
timestamp 1712256841
transform 1 0 1076 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1712256841
transform 1 0 812 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1712256841
transform 1 0 516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1712256841
transform 1 0 372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4372
timestamp 1712256841
transform 1 0 372 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1712256841
transform 1 0 340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4374
timestamp 1712256841
transform 1 0 316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4375
timestamp 1712256841
transform 1 0 292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1712256841
transform 1 0 292 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1712256841
transform 1 0 260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4378
timestamp 1712256841
transform 1 0 252 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4379
timestamp 1712256841
transform 1 0 948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1712256841
transform 1 0 356 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1712256841
transform 1 0 348 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4382
timestamp 1712256841
transform 1 0 1092 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4383
timestamp 1712256841
transform 1 0 388 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_4384
timestamp 1712256841
transform 1 0 340 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_4385
timestamp 1712256841
transform 1 0 268 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4386
timestamp 1712256841
transform 1 0 196 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4387
timestamp 1712256841
transform 1 0 188 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4388
timestamp 1712256841
transform 1 0 988 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4389
timestamp 1712256841
transform 1 0 500 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4390
timestamp 1712256841
transform 1 0 516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4391
timestamp 1712256841
transform 1 0 492 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4392
timestamp 1712256841
transform 1 0 180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4393
timestamp 1712256841
transform 1 0 164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4394
timestamp 1712256841
transform 1 0 996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4395
timestamp 1712256841
transform 1 0 980 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1712256841
transform 1 0 196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4397
timestamp 1712256841
transform 1 0 108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4398
timestamp 1712256841
transform 1 0 220 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4399
timestamp 1712256841
transform 1 0 212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4400
timestamp 1712256841
transform 1 0 1180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1712256841
transform 1 0 924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1712256841
transform 1 0 1268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1712256841
transform 1 0 1196 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4404
timestamp 1712256841
transform 1 0 1116 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1712256841
transform 1 0 1092 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4406
timestamp 1712256841
transform 1 0 1012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4407
timestamp 1712256841
transform 1 0 900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4408
timestamp 1712256841
transform 1 0 788 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4409
timestamp 1712256841
transform 1 0 1212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4410
timestamp 1712256841
transform 1 0 1068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4411
timestamp 1712256841
transform 1 0 1172 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4412
timestamp 1712256841
transform 1 0 1076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4413
timestamp 1712256841
transform 1 0 1124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4414
timestamp 1712256841
transform 1 0 1124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4415
timestamp 1712256841
transform 1 0 940 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4416
timestamp 1712256841
transform 1 0 932 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4417
timestamp 1712256841
transform 1 0 916 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4418
timestamp 1712256841
transform 1 0 884 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4419
timestamp 1712256841
transform 1 0 884 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4420
timestamp 1712256841
transform 1 0 676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4421
timestamp 1712256841
transform 1 0 1108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1712256841
transform 1 0 1084 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4423
timestamp 1712256841
transform 1 0 1740 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4424
timestamp 1712256841
transform 1 0 1340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1712256841
transform 1 0 1156 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4426
timestamp 1712256841
transform 1 0 1156 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1712256841
transform 1 0 244 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4428
timestamp 1712256841
transform 1 0 244 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1712256841
transform 1 0 244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4430
timestamp 1712256841
transform 1 0 220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4431
timestamp 1712256841
transform 1 0 212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4432
timestamp 1712256841
transform 1 0 212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1712256841
transform 1 0 356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4434
timestamp 1712256841
transform 1 0 220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4435
timestamp 1712256841
transform 1 0 572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4436
timestamp 1712256841
transform 1 0 388 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1712256841
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4438
timestamp 1712256841
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4439
timestamp 1712256841
transform 1 0 740 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4440
timestamp 1712256841
transform 1 0 500 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4441
timestamp 1712256841
transform 1 0 452 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4442
timestamp 1712256841
transform 1 0 444 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4443
timestamp 1712256841
transform 1 0 1220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1712256841
transform 1 0 708 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1712256841
transform 1 0 652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4446
timestamp 1712256841
transform 1 0 468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4447
timestamp 1712256841
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1712256841
transform 1 0 420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4449
timestamp 1712256841
transform 1 0 324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4450
timestamp 1712256841
transform 1 0 324 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4451
timestamp 1712256841
transform 1 0 276 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1712256841
transform 1 0 228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4453
timestamp 1712256841
transform 1 0 748 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1712256841
transform 1 0 644 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4455
timestamp 1712256841
transform 1 0 860 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1712256841
transform 1 0 796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4457
timestamp 1712256841
transform 1 0 756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4458
timestamp 1712256841
transform 1 0 708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4459
timestamp 1712256841
transform 1 0 204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4460
timestamp 1712256841
transform 1 0 108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4461
timestamp 1712256841
transform 1 0 292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4462
timestamp 1712256841
transform 1 0 252 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1712256841
transform 1 0 772 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1712256841
transform 1 0 740 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1712256841
transform 1 0 844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4466
timestamp 1712256841
transform 1 0 324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4467
timestamp 1712256841
transform 1 0 940 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4468
timestamp 1712256841
transform 1 0 812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4469
timestamp 1712256841
transform 1 0 860 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4470
timestamp 1712256841
transform 1 0 844 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4471
timestamp 1712256841
transform 1 0 852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1712256841
transform 1 0 836 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1712256841
transform 1 0 1004 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4474
timestamp 1712256841
transform 1 0 908 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1712256841
transform 1 0 852 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4476
timestamp 1712256841
transform 1 0 652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1712256841
transform 1 0 988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4478
timestamp 1712256841
transform 1 0 964 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_4479
timestamp 1712256841
transform 1 0 2788 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4480
timestamp 1712256841
transform 1 0 2764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1712256841
transform 1 0 1884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4482
timestamp 1712256841
transform 1 0 1844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4483
timestamp 1712256841
transform 1 0 1588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1712256841
transform 1 0 1372 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4485
timestamp 1712256841
transform 1 0 1315 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1712256841
transform 1 0 1292 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1712256841
transform 1 0 148 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4488
timestamp 1712256841
transform 1 0 132 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4489
timestamp 1712256841
transform 1 0 132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1712256841
transform 1 0 84 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1712256841
transform 1 0 420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4492
timestamp 1712256841
transform 1 0 108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4493
timestamp 1712256841
transform 1 0 516 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4494
timestamp 1712256841
transform 1 0 444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1712256841
transform 1 0 476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1712256841
transform 1 0 468 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4497
timestamp 1712256841
transform 1 0 668 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4498
timestamp 1712256841
transform 1 0 580 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4499
timestamp 1712256841
transform 1 0 724 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1712256841
transform 1 0 724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1712256841
transform 1 0 676 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4502
timestamp 1712256841
transform 1 0 596 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1712256841
transform 1 0 132 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4504
timestamp 1712256841
transform 1 0 108 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4505
timestamp 1712256841
transform 1 0 228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4506
timestamp 1712256841
transform 1 0 196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4507
timestamp 1712256841
transform 1 0 620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4508
timestamp 1712256841
transform 1 0 452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4509
timestamp 1712256841
transform 1 0 708 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4510
timestamp 1712256841
transform 1 0 644 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4511
timestamp 1712256841
transform 1 0 780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4512
timestamp 1712256841
transform 1 0 180 0 1 1095
box -2 -2 2 2
use M2_M1  M2_M1_4513
timestamp 1712256841
transform 1 0 180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1712256841
transform 1 0 164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4515
timestamp 1712256841
transform 1 0 164 0 1 1095
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1712256841
transform 1 0 860 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1712256841
transform 1 0 756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4518
timestamp 1712256841
transform 1 0 868 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4519
timestamp 1712256841
transform 1 0 796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4520
timestamp 1712256841
transform 1 0 884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1712256841
transform 1 0 860 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1712256841
transform 1 0 932 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1712256841
transform 1 0 796 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4524
timestamp 1712256841
transform 1 0 740 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4525
timestamp 1712256841
transform 1 0 740 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1712256841
transform 1 0 988 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1712256841
transform 1 0 868 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1712256841
transform 1 0 180 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4529
timestamp 1712256841
transform 1 0 116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4530
timestamp 1712256841
transform 1 0 84 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4531
timestamp 1712256841
transform 1 0 84 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1712256841
transform 1 0 380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1712256841
transform 1 0 84 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1712256841
transform 1 0 516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4535
timestamp 1712256841
transform 1 0 404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4536
timestamp 1712256841
transform 1 0 452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4537
timestamp 1712256841
transform 1 0 444 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4538
timestamp 1712256841
transform 1 0 668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4539
timestamp 1712256841
transform 1 0 468 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4540
timestamp 1712256841
transform 1 0 452 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4541
timestamp 1712256841
transform 1 0 1060 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1712256841
transform 1 0 1052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4543
timestamp 1712256841
transform 1 0 1044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4544
timestamp 1712256841
transform 1 0 988 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4545
timestamp 1712256841
transform 1 0 884 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1712256841
transform 1 0 580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4547
timestamp 1712256841
transform 1 0 276 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4548
timestamp 1712256841
transform 1 0 228 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1712256841
transform 1 0 228 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4550
timestamp 1712256841
transform 1 0 700 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1712256841
transform 1 0 564 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4552
timestamp 1712256841
transform 1 0 732 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4553
timestamp 1712256841
transform 1 0 628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4554
timestamp 1712256841
transform 1 0 628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4555
timestamp 1712256841
transform 1 0 108 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4556
timestamp 1712256841
transform 1 0 84 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4557
timestamp 1712256841
transform 1 0 164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4558
timestamp 1712256841
transform 1 0 140 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4559
timestamp 1712256841
transform 1 0 724 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4560
timestamp 1712256841
transform 1 0 692 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4561
timestamp 1712256841
transform 1 0 796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4562
timestamp 1712256841
transform 1 0 212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4563
timestamp 1712256841
transform 1 0 844 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1712256841
transform 1 0 756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4565
timestamp 1712256841
transform 1 0 860 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4566
timestamp 1712256841
transform 1 0 820 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1712256841
transform 1 0 868 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4568
timestamp 1712256841
transform 1 0 836 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1712256841
transform 1 0 1308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4570
timestamp 1712256841
transform 1 0 1284 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1712256841
transform 1 0 1124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4572
timestamp 1712256841
transform 1 0 1060 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1712256841
transform 1 0 1004 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4574
timestamp 1712256841
transform 1 0 988 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4575
timestamp 1712256841
transform 1 0 980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4576
timestamp 1712256841
transform 1 0 900 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4577
timestamp 1712256841
transform 1 0 860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1712256841
transform 1 0 972 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1712256841
transform 1 0 844 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1712256841
transform 1 0 2956 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1712256841
transform 1 0 2916 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4582
timestamp 1712256841
transform 1 0 2572 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1712256841
transform 1 0 2412 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4584
timestamp 1712256841
transform 1 0 1276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4585
timestamp 1712256841
transform 1 0 1236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4586
timestamp 1712256841
transform 1 0 1068 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4587
timestamp 1712256841
transform 1 0 644 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4588
timestamp 1712256841
transform 1 0 284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4589
timestamp 1712256841
transform 1 0 228 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4590
timestamp 1712256841
transform 1 0 132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4591
timestamp 1712256841
transform 1 0 340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1712256841
transform 1 0 236 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4593
timestamp 1712256841
transform 1 0 620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4594
timestamp 1712256841
transform 1 0 316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4595
timestamp 1712256841
transform 1 0 412 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4596
timestamp 1712256841
transform 1 0 380 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4597
timestamp 1712256841
transform 1 0 1268 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1712256841
transform 1 0 1244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4599
timestamp 1712256841
transform 1 0 1188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1712256841
transform 1 0 1060 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4601
timestamp 1712256841
transform 1 0 676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4602
timestamp 1712256841
transform 1 0 460 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4603
timestamp 1712256841
transform 1 0 444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4604
timestamp 1712256841
transform 1 0 412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1712256841
transform 1 0 284 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4606
timestamp 1712256841
transform 1 0 596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4607
timestamp 1712256841
transform 1 0 460 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1712256841
transform 1 0 316 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4609
timestamp 1712256841
transform 1 0 964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4610
timestamp 1712256841
transform 1 0 516 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1712256841
transform 1 0 252 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_4612
timestamp 1712256841
transform 1 0 180 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1712256841
transform 1 0 180 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4614
timestamp 1712256841
transform 1 0 932 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4615
timestamp 1712256841
transform 1 0 676 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4616
timestamp 1712256841
transform 1 0 908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4617
timestamp 1712256841
transform 1 0 908 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1712256841
transform 1 0 108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4619
timestamp 1712256841
transform 1 0 100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1712256841
transform 1 0 220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1712256841
transform 1 0 140 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4622
timestamp 1712256841
transform 1 0 1156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4623
timestamp 1712256841
transform 1 0 628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4624
timestamp 1712256841
transform 1 0 1388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4625
timestamp 1712256841
transform 1 0 1388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4626
timestamp 1712256841
transform 1 0 1172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4627
timestamp 1712256841
transform 1 0 1076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4628
timestamp 1712256841
transform 1 0 1068 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1712256841
transform 1 0 1036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4630
timestamp 1712256841
transform 1 0 1276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4631
timestamp 1712256841
transform 1 0 940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4632
timestamp 1712256841
transform 1 0 996 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1712256841
transform 1 0 948 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4634
timestamp 1712256841
transform 1 0 1060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4635
timestamp 1712256841
transform 1 0 980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4636
timestamp 1712256841
transform 1 0 1684 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4637
timestamp 1712256841
transform 1 0 1596 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1712256841
transform 1 0 1380 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4639
timestamp 1712256841
transform 1 0 1020 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4640
timestamp 1712256841
transform 1 0 1084 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4641
timestamp 1712256841
transform 1 0 1076 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4642
timestamp 1712256841
transform 1 0 2980 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4643
timestamp 1712256841
transform 1 0 2956 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1712256841
transform 1 0 2476 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1712256841
transform 1 0 1772 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4646
timestamp 1712256841
transform 1 0 1404 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4647
timestamp 1712256841
transform 1 0 1388 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4648
timestamp 1712256841
transform 1 0 1388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4649
timestamp 1712256841
transform 1 0 1148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4650
timestamp 1712256841
transform 1 0 1076 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4651
timestamp 1712256841
transform 1 0 2708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4652
timestamp 1712256841
transform 1 0 2540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4653
timestamp 1712256841
transform 1 0 1740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1712256841
transform 1 0 1500 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1712256841
transform 1 0 1348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1712256841
transform 1 0 1036 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4657
timestamp 1712256841
transform 1 0 252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1712256841
transform 1 0 204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4659
timestamp 1712256841
transform 1 0 204 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1712256841
transform 1 0 252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4661
timestamp 1712256841
transform 1 0 236 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4662
timestamp 1712256841
transform 1 0 788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4663
timestamp 1712256841
transform 1 0 260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4664
timestamp 1712256841
transform 1 0 412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1712256841
transform 1 0 324 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4666
timestamp 1712256841
transform 1 0 788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4667
timestamp 1712256841
transform 1 0 396 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4668
timestamp 1712256841
transform 1 0 300 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1712256841
transform 1 0 1020 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4670
timestamp 1712256841
transform 1 0 580 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4671
timestamp 1712256841
transform 1 0 284 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_4672
timestamp 1712256841
transform 1 0 236 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1712256841
transform 1 0 156 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1712256841
transform 1 0 1060 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4675
timestamp 1712256841
transform 1 0 1012 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4676
timestamp 1712256841
transform 1 0 804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4677
timestamp 1712256841
transform 1 0 804 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1712256841
transform 1 0 796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4679
timestamp 1712256841
transform 1 0 908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4680
timestamp 1712256841
transform 1 0 756 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1712256841
transform 1 0 900 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4682
timestamp 1712256841
transform 1 0 860 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4683
timestamp 1712256841
transform 1 0 156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4684
timestamp 1712256841
transform 1 0 156 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_4685
timestamp 1712256841
transform 1 0 252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1712256841
transform 1 0 236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1712256841
transform 1 0 1204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4688
timestamp 1712256841
transform 1 0 988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4689
timestamp 1712256841
transform 1 0 1188 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1712256841
transform 1 0 1164 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4691
timestamp 1712256841
transform 1 0 2908 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4692
timestamp 1712256841
transform 1 0 2844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4693
timestamp 1712256841
transform 1 0 2508 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4694
timestamp 1712256841
transform 1 0 1844 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4695
timestamp 1712256841
transform 1 0 1804 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1712256841
transform 1 0 1572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1712256841
transform 1 0 1412 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1712256841
transform 1 0 1092 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4699
timestamp 1712256841
transform 1 0 1148 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4700
timestamp 1712256841
transform 1 0 644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4701
timestamp 1712256841
transform 1 0 620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4702
timestamp 1712256841
transform 1 0 412 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4703
timestamp 1712256841
transform 1 0 636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1712256841
transform 1 0 596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1712256841
transform 1 0 612 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1712256841
transform 1 0 492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4707
timestamp 1712256841
transform 1 0 692 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1712256841
transform 1 0 540 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4709
timestamp 1712256841
transform 1 0 516 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1712256841
transform 1 0 636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4711
timestamp 1712256841
transform 1 0 588 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4712
timestamp 1712256841
transform 1 0 532 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1712256841
transform 1 0 388 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1712256841
transform 1 0 372 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1712256841
transform 1 0 1204 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4716
timestamp 1712256841
transform 1 0 732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4717
timestamp 1712256841
transform 1 0 692 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1712256841
transform 1 0 644 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1712256841
transform 1 0 644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4720
timestamp 1712256841
transform 1 0 812 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1712256841
transform 1 0 692 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1712256841
transform 1 0 796 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1712256841
transform 1 0 756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4724
timestamp 1712256841
transform 1 0 516 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4725
timestamp 1712256841
transform 1 0 404 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1712256841
transform 1 0 420 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1712256841
transform 1 0 340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1712256841
transform 1 0 1588 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1712256841
transform 1 0 1524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1712256841
transform 1 0 1484 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4731
timestamp 1712256841
transform 1 0 1268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4732
timestamp 1712256841
transform 1 0 1268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4733
timestamp 1712256841
transform 1 0 1172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1712256841
transform 1 0 2748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4735
timestamp 1712256841
transform 1 0 2460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4736
timestamp 1712256841
transform 1 0 1268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1712256841
transform 1 0 1244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4738
timestamp 1712256841
transform 1 0 1204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4739
timestamp 1712256841
transform 1 0 1068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1712256841
transform 1 0 1060 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4741
timestamp 1712256841
transform 1 0 1060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1712256841
transform 1 0 1028 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1712256841
transform 1 0 1028 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4744
timestamp 1712256841
transform 1 0 1004 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4745
timestamp 1712256841
transform 1 0 1388 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1712256841
transform 1 0 892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4747
timestamp 1712256841
transform 1 0 868 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4748
timestamp 1712256841
transform 1 0 868 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4749
timestamp 1712256841
transform 1 0 900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4750
timestamp 1712256841
transform 1 0 868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1712256841
transform 1 0 940 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4752
timestamp 1712256841
transform 1 0 900 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1712256841
transform 1 0 980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1712256841
transform 1 0 948 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1712256841
transform 1 0 2444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4756
timestamp 1712256841
transform 1 0 2428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4757
timestamp 1712256841
transform 1 0 2404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1712256841
transform 1 0 2260 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4759
timestamp 1712256841
transform 1 0 1492 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4760
timestamp 1712256841
transform 1 0 956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4761
timestamp 1712256841
transform 1 0 956 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1712256841
transform 1 0 916 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4763
timestamp 1712256841
transform 1 0 916 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4764
timestamp 1712256841
transform 1 0 876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1712256841
transform 1 0 812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4766
timestamp 1712256841
transform 1 0 932 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4767
timestamp 1712256841
transform 1 0 924 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4768
timestamp 1712256841
transform 1 0 916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4769
timestamp 1712256841
transform 1 0 948 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4770
timestamp 1712256841
transform 1 0 932 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4771
timestamp 1712256841
transform 1 0 852 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1712256841
transform 1 0 844 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4773
timestamp 1712256841
transform 1 0 828 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1712256841
transform 1 0 1252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4775
timestamp 1712256841
transform 1 0 1124 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4776
timestamp 1712256841
transform 1 0 948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4777
timestamp 1712256841
transform 1 0 908 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1712256841
transform 1 0 884 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4779
timestamp 1712256841
transform 1 0 980 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4780
timestamp 1712256841
transform 1 0 956 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4781
timestamp 1712256841
transform 1 0 844 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4782
timestamp 1712256841
transform 1 0 828 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1712256841
transform 1 0 940 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4784
timestamp 1712256841
transform 1 0 916 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1712256841
transform 1 0 1796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4786
timestamp 1712256841
transform 1 0 1740 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4787
timestamp 1712256841
transform 1 0 1620 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4788
timestamp 1712256841
transform 1 0 1324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1712256841
transform 1 0 1316 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4790
timestamp 1712256841
transform 1 0 1228 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4791
timestamp 1712256841
transform 1 0 1444 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4792
timestamp 1712256841
transform 1 0 1220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4793
timestamp 1712256841
transform 1 0 1196 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1712256841
transform 1 0 1180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4795
timestamp 1712256841
transform 1 0 1172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4796
timestamp 1712256841
transform 1 0 1172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1712256841
transform 1 0 1116 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1712256841
transform 1 0 1116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4799
timestamp 1712256841
transform 1 0 1140 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4800
timestamp 1712256841
transform 1 0 1116 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4801
timestamp 1712256841
transform 1 0 1140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4802
timestamp 1712256841
transform 1 0 1092 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4803
timestamp 1712256841
transform 1 0 1076 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4804
timestamp 1712256841
transform 1 0 1228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4805
timestamp 1712256841
transform 1 0 1140 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_4806
timestamp 1712256841
transform 1 0 1092 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4807
timestamp 1712256841
transform 1 0 1052 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_4808
timestamp 1712256841
transform 1 0 1052 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4809
timestamp 1712256841
transform 1 0 1108 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4810
timestamp 1712256841
transform 1 0 1044 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4811
timestamp 1712256841
transform 1 0 1084 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4812
timestamp 1712256841
transform 1 0 1068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4813
timestamp 1712256841
transform 1 0 1156 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4814
timestamp 1712256841
transform 1 0 1140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4815
timestamp 1712256841
transform 1 0 1204 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4816
timestamp 1712256841
transform 1 0 1188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1712256841
transform 1 0 1180 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4818
timestamp 1712256841
transform 1 0 1156 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4819
timestamp 1712256841
transform 1 0 1764 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1712256841
transform 1 0 1668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4821
timestamp 1712256841
transform 1 0 1532 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4822
timestamp 1712256841
transform 1 0 1420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4823
timestamp 1712256841
transform 1 0 1412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4824
timestamp 1712256841
transform 1 0 1196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4825
timestamp 1712256841
transform 1 0 1132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4826
timestamp 1712256841
transform 1 0 1196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4827
timestamp 1712256841
transform 1 0 1188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4828
timestamp 1712256841
transform 1 0 2004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4829
timestamp 1712256841
transform 1 0 1844 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4830
timestamp 1712256841
transform 1 0 1724 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1712256841
transform 1 0 1652 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1712256841
transform 1 0 1652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4833
timestamp 1712256841
transform 1 0 1516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4834
timestamp 1712256841
transform 1 0 1452 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4835
timestamp 1712256841
transform 1 0 1436 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1712256841
transform 1 0 1084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1712256841
transform 1 0 1060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4838
timestamp 1712256841
transform 1 0 1548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4839
timestamp 1712256841
transform 1 0 1524 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4840
timestamp 1712256841
transform 1 0 1484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4841
timestamp 1712256841
transform 1 0 1484 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4842
timestamp 1712256841
transform 1 0 1468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4843
timestamp 1712256841
transform 1 0 1444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4844
timestamp 1712256841
transform 1 0 1468 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4845
timestamp 1712256841
transform 1 0 1316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4846
timestamp 1712256841
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4847
timestamp 1712256841
transform 1 0 1332 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_4848
timestamp 1712256841
transform 1 0 1332 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_4849
timestamp 1712256841
transform 1 0 1516 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4850
timestamp 1712256841
transform 1 0 1516 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1712256841
transform 1 0 1444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4852
timestamp 1712256841
transform 1 0 1332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4853
timestamp 1712256841
transform 1 0 1332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4854
timestamp 1712256841
transform 1 0 1252 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4855
timestamp 1712256841
transform 1 0 1516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1712256841
transform 1 0 1508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4857
timestamp 1712256841
transform 1 0 1532 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4858
timestamp 1712256841
transform 1 0 1460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1712256841
transform 1 0 1372 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4860
timestamp 1712256841
transform 1 0 1340 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1712256841
transform 1 0 1396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4862
timestamp 1712256841
transform 1 0 1364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4863
timestamp 1712256841
transform 1 0 1364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4864
timestamp 1712256841
transform 1 0 1412 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4865
timestamp 1712256841
transform 1 0 1396 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4866
timestamp 1712256841
transform 1 0 1500 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4867
timestamp 1712256841
transform 1 0 1404 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1712256841
transform 1 0 1620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1712256841
transform 1 0 1620 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4870
timestamp 1712256841
transform 1 0 1532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4871
timestamp 1712256841
transform 1 0 1300 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4872
timestamp 1712256841
transform 1 0 1292 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4873
timestamp 1712256841
transform 1 0 1908 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4874
timestamp 1712256841
transform 1 0 1884 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4875
timestamp 1712256841
transform 1 0 1820 0 1 455
box -2 -2 2 2
use M2_M1  M2_M1_4876
timestamp 1712256841
transform 1 0 1820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4877
timestamp 1712256841
transform 1 0 1804 0 1 455
box -2 -2 2 2
use M2_M1  M2_M1_4878
timestamp 1712256841
transform 1 0 1708 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4879
timestamp 1712256841
transform 1 0 1700 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4880
timestamp 1712256841
transform 1 0 1700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1712256841
transform 1 0 1772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1712256841
transform 1 0 1772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4883
timestamp 1712256841
transform 1 0 1796 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1712256841
transform 1 0 1780 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4885
timestamp 1712256841
transform 1 0 1828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4886
timestamp 1712256841
transform 1 0 1828 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1712256841
transform 1 0 1868 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1712256841
transform 1 0 1868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4889
timestamp 1712256841
transform 1 0 1788 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1712256841
transform 1 0 1764 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4891
timestamp 1712256841
transform 1 0 1708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4892
timestamp 1712256841
transform 1 0 1652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1712256841
transform 1 0 1612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4894
timestamp 1712256841
transform 1 0 1612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1712256841
transform 1 0 1756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4896
timestamp 1712256841
transform 1 0 1740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1712256841
transform 1 0 1804 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4898
timestamp 1712256841
transform 1 0 1780 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4899
timestamp 1712256841
transform 1 0 1660 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4900
timestamp 1712256841
transform 1 0 1652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1712256841
transform 1 0 1644 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4902
timestamp 1712256841
transform 1 0 1636 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4903
timestamp 1712256841
transform 1 0 1708 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4904
timestamp 1712256841
transform 1 0 1700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1712256841
transform 1 0 1700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4906
timestamp 1712256841
transform 1 0 1684 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1712256841
transform 1 0 1772 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4908
timestamp 1712256841
transform 1 0 1716 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4909
timestamp 1712256841
transform 1 0 1764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4910
timestamp 1712256841
transform 1 0 1764 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1712256841
transform 1 0 1900 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1712256841
transform 1 0 1852 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4913
timestamp 1712256841
transform 1 0 1780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1712256841
transform 1 0 1780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4915
timestamp 1712256841
transform 1 0 1780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4916
timestamp 1712256841
transform 1 0 1700 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4917
timestamp 1712256841
transform 1 0 1372 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1712256841
transform 1 0 2060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4919
timestamp 1712256841
transform 1 0 1828 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4920
timestamp 1712256841
transform 1 0 1516 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1712256841
transform 1 0 1508 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4922
timestamp 1712256841
transform 1 0 1500 0 1 1895
box -2 -2 2 2
use M2_M1  M2_M1_4923
timestamp 1712256841
transform 1 0 1500 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4924
timestamp 1712256841
transform 1 0 2188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4925
timestamp 1712256841
transform 1 0 2036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4926
timestamp 1712256841
transform 1 0 2060 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4927
timestamp 1712256841
transform 1 0 2044 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4928
timestamp 1712256841
transform 1 0 2068 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4929
timestamp 1712256841
transform 1 0 2060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4930
timestamp 1712256841
transform 1 0 2140 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1712256841
transform 1 0 2140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1712256841
transform 1 0 1908 0 1 695
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1712256841
transform 1 0 1876 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4934
timestamp 1712256841
transform 1 0 2044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1712256841
transform 1 0 1852 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_4936
timestamp 1712256841
transform 1 0 836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1712256841
transform 1 0 636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4938
timestamp 1712256841
transform 1 0 2004 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4939
timestamp 1712256841
transform 1 0 1932 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4940
timestamp 1712256841
transform 1 0 1924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4941
timestamp 1712256841
transform 1 0 1924 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4942
timestamp 1712256841
transform 1 0 2180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1712256841
transform 1 0 2164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4944
timestamp 1712256841
transform 1 0 2332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4945
timestamp 1712256841
transform 1 0 2276 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4946
timestamp 1712256841
transform 1 0 2068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4947
timestamp 1712256841
transform 1 0 2068 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1712256841
transform 1 0 2044 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4949
timestamp 1712256841
transform 1 0 2028 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4950
timestamp 1712256841
transform 1 0 2020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4951
timestamp 1712256841
transform 1 0 2012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4952
timestamp 1712256841
transform 1 0 2012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4953
timestamp 1712256841
transform 1 0 1924 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4954
timestamp 1712256841
transform 1 0 1884 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4955
timestamp 1712256841
transform 1 0 1988 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4956
timestamp 1712256841
transform 1 0 1956 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1712256841
transform 1 0 1884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1712256841
transform 1 0 1884 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1712256841
transform 1 0 2188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4960
timestamp 1712256841
transform 1 0 1972 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1712256841
transform 1 0 1908 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4962
timestamp 1712256841
transform 1 0 1876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1712256841
transform 1 0 1876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4964
timestamp 1712256841
transform 1 0 1868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4965
timestamp 1712256841
transform 1 0 1860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4966
timestamp 1712256841
transform 1 0 1860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4967
timestamp 1712256841
transform 1 0 1844 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4968
timestamp 1712256841
transform 1 0 1564 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4969
timestamp 1712256841
transform 1 0 2380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1712256841
transform 1 0 1924 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4971
timestamp 1712256841
transform 1 0 2332 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4972
timestamp 1712256841
transform 1 0 2308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4973
timestamp 1712256841
transform 1 0 2388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4974
timestamp 1712256841
transform 1 0 2300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1712256841
transform 1 0 2500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4976
timestamp 1712256841
transform 1 0 2412 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4977
timestamp 1712256841
transform 1 0 2436 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4978
timestamp 1712256841
transform 1 0 2396 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4979
timestamp 1712256841
transform 1 0 2180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4980
timestamp 1712256841
transform 1 0 2404 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1712256841
transform 1 0 2388 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4982
timestamp 1712256841
transform 1 0 2340 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4983
timestamp 1712256841
transform 1 0 2140 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4984
timestamp 1712256841
transform 1 0 2092 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4985
timestamp 1712256841
transform 1 0 1804 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4986
timestamp 1712256841
transform 1 0 2020 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4987
timestamp 1712256841
transform 1 0 1948 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4988
timestamp 1712256841
transform 1 0 1900 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4989
timestamp 1712256841
transform 1 0 1796 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1712256841
transform 1 0 2220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4991
timestamp 1712256841
transform 1 0 2220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4992
timestamp 1712256841
transform 1 0 2308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4993
timestamp 1712256841
transform 1 0 2292 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4994
timestamp 1712256841
transform 1 0 2140 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1712256841
transform 1 0 2052 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4996
timestamp 1712256841
transform 1 0 2420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1712256841
transform 1 0 2204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4998
timestamp 1712256841
transform 1 0 2068 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4999
timestamp 1712256841
transform 1 0 2020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5000
timestamp 1712256841
transform 1 0 2020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5001
timestamp 1712256841
transform 1 0 1940 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1712256841
transform 1 0 1748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5003
timestamp 1712256841
transform 1 0 1724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5004
timestamp 1712256841
transform 1 0 1684 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5005
timestamp 1712256841
transform 1 0 1668 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5006
timestamp 1712256841
transform 1 0 1684 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_5007
timestamp 1712256841
transform 1 0 1604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1712256841
transform 1 0 1724 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5009
timestamp 1712256841
transform 1 0 1716 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5010
timestamp 1712256841
transform 1 0 1692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5011
timestamp 1712256841
transform 1 0 1692 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5012
timestamp 1712256841
transform 1 0 1516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5013
timestamp 1712256841
transform 1 0 1476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5014
timestamp 1712256841
transform 1 0 2332 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5015
timestamp 1712256841
transform 1 0 2156 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5016
timestamp 1712256841
transform 1 0 2300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5017
timestamp 1712256841
transform 1 0 2292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5018
timestamp 1712256841
transform 1 0 2436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5019
timestamp 1712256841
transform 1 0 2300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5020
timestamp 1712256841
transform 1 0 2444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5021
timestamp 1712256841
transform 1 0 2364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5022
timestamp 1712256841
transform 1 0 2524 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5023
timestamp 1712256841
transform 1 0 2500 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1712256841
transform 1 0 2564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5025
timestamp 1712256841
transform 1 0 2564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5026
timestamp 1712256841
transform 1 0 2404 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5027
timestamp 1712256841
transform 1 0 2340 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5028
timestamp 1712256841
transform 1 0 2284 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5029
timestamp 1712256841
transform 1 0 2260 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1712256841
transform 1 0 2220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1712256841
transform 1 0 2052 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_5032
timestamp 1712256841
transform 1 0 2028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1712256841
transform 1 0 1988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5034
timestamp 1712256841
transform 1 0 2588 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5035
timestamp 1712256841
transform 1 0 2532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5036
timestamp 1712256841
transform 1 0 2532 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5037
timestamp 1712256841
transform 1 0 2388 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5038
timestamp 1712256841
transform 1 0 2340 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5039
timestamp 1712256841
transform 1 0 2204 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1712256841
transform 1 0 2172 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5041
timestamp 1712256841
transform 1 0 1604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1712256841
transform 1 0 2084 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1712256841
transform 1 0 1660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5044
timestamp 1712256841
transform 1 0 1644 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5045
timestamp 1712256841
transform 1 0 1620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5046
timestamp 1712256841
transform 1 0 2292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5047
timestamp 1712256841
transform 1 0 2236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1712256841
transform 1 0 2404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5049
timestamp 1712256841
transform 1 0 2340 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5050
timestamp 1712256841
transform 1 0 1500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5051
timestamp 1712256841
transform 1 0 1468 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5052
timestamp 1712256841
transform 1 0 1556 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1712256841
transform 1 0 1468 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5054
timestamp 1712256841
transform 1 0 1692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5055
timestamp 1712256841
transform 1 0 1556 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1712256841
transform 1 0 1604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1712256841
transform 1 0 1444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5058
timestamp 1712256841
transform 1 0 3052 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5059
timestamp 1712256841
transform 1 0 2972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5060
timestamp 1712256841
transform 1 0 2884 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5061
timestamp 1712256841
transform 1 0 2716 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5062
timestamp 1712256841
transform 1 0 2668 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1712256841
transform 1 0 2564 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1712256841
transform 1 0 1652 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1712256841
transform 1 0 1612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5066
timestamp 1712256841
transform 1 0 1604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5067
timestamp 1712256841
transform 1 0 2276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1712256841
transform 1 0 2268 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5069
timestamp 1712256841
transform 1 0 2220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1712256841
transform 1 0 2180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5071
timestamp 1712256841
transform 1 0 2500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1712256841
transform 1 0 2260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5073
timestamp 1712256841
transform 1 0 2516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5074
timestamp 1712256841
transform 1 0 2388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1712256841
transform 1 0 2548 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5076
timestamp 1712256841
transform 1 0 2476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1712256841
transform 1 0 2348 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5078
timestamp 1712256841
transform 1 0 2340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5079
timestamp 1712256841
transform 1 0 2308 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5080
timestamp 1712256841
transform 1 0 2228 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5081
timestamp 1712256841
transform 1 0 2228 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1712256841
transform 1 0 2196 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5083
timestamp 1712256841
transform 1 0 2140 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5084
timestamp 1712256841
transform 1 0 2052 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5085
timestamp 1712256841
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5086
timestamp 1712256841
transform 1 0 2396 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5087
timestamp 1712256841
transform 1 0 2348 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1712256841
transform 1 0 2292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1712256841
transform 1 0 2004 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1712256841
transform 1 0 1964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1712256841
transform 1 0 2052 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1712256841
transform 1 0 1948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5093
timestamp 1712256841
transform 1 0 1948 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5094
timestamp 1712256841
transform 1 0 1940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5095
timestamp 1712256841
transform 1 0 2108 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1712256841
transform 1 0 2100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1712256841
transform 1 0 2180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5098
timestamp 1712256841
transform 1 0 2172 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1712256841
transform 1 0 2540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5100
timestamp 1712256841
transform 1 0 2436 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1712256841
transform 1 0 2412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1712256841
transform 1 0 2356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1712256841
transform 1 0 2244 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5104
timestamp 1712256841
transform 1 0 2116 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1712256841
transform 1 0 1428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5106
timestamp 1712256841
transform 1 0 1348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5107
timestamp 1712256841
transform 1 0 2708 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1712256841
transform 1 0 1796 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1712256841
transform 1 0 1388 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1712256841
transform 1 0 1468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1712256841
transform 1 0 1468 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5112
timestamp 1712256841
transform 1 0 2716 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5113
timestamp 1712256841
transform 1 0 2604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1712256841
transform 1 0 2572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5115
timestamp 1712256841
transform 1 0 2468 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5116
timestamp 1712256841
transform 1 0 2444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5117
timestamp 1712256841
transform 1 0 2308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5118
timestamp 1712256841
transform 1 0 2260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5119
timestamp 1712256841
transform 1 0 1572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5120
timestamp 1712256841
transform 1 0 1404 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5121
timestamp 1712256841
transform 1 0 2396 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5122
timestamp 1712256841
transform 1 0 2356 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5123
timestamp 1712256841
transform 1 0 2300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5124
timestamp 1712256841
transform 1 0 2244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5125
timestamp 1712256841
transform 1 0 2444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5126
timestamp 1712256841
transform 1 0 2340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5127
timestamp 1712256841
transform 1 0 2492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5128
timestamp 1712256841
transform 1 0 2420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5129
timestamp 1712256841
transform 1 0 2612 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5130
timestamp 1712256841
transform 1 0 2524 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5131
timestamp 1712256841
transform 1 0 2548 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5132
timestamp 1712256841
transform 1 0 2356 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5133
timestamp 1712256841
transform 1 0 2316 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5134
timestamp 1712256841
transform 1 0 2172 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1712256841
transform 1 0 2100 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5136
timestamp 1712256841
transform 1 0 2084 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5137
timestamp 1712256841
transform 1 0 2052 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5138
timestamp 1712256841
transform 1 0 2428 0 1 1136
box -2 -2 2 2
use M2_M1  M2_M1_5139
timestamp 1712256841
transform 1 0 2364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5140
timestamp 1712256841
transform 1 0 2356 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5141
timestamp 1712256841
transform 1 0 2084 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5142
timestamp 1712256841
transform 1 0 2052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5143
timestamp 1712256841
transform 1 0 1980 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5144
timestamp 1712256841
transform 1 0 1972 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5145
timestamp 1712256841
transform 1 0 1980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5146
timestamp 1712256841
transform 1 0 1980 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1712256841
transform 1 0 2172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5148
timestamp 1712256841
transform 1 0 2148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5149
timestamp 1712256841
transform 1 0 2268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5150
timestamp 1712256841
transform 1 0 2236 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5151
timestamp 1712256841
transform 1 0 2468 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5152
timestamp 1712256841
transform 1 0 2436 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5153
timestamp 1712256841
transform 1 0 2428 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5154
timestamp 1712256841
transform 1 0 2380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5155
timestamp 1712256841
transform 1 0 2300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5156
timestamp 1712256841
transform 1 0 2604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1712256841
transform 1 0 1860 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5158
timestamp 1712256841
transform 1 0 1764 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5159
timestamp 1712256841
transform 1 0 1652 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5160
timestamp 1712256841
transform 1 0 1572 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5161
timestamp 1712256841
transform 1 0 1620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5162
timestamp 1712256841
transform 1 0 1588 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1712256841
transform 1 0 2012 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5164
timestamp 1712256841
transform 1 0 1892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1712256841
transform 1 0 1828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5166
timestamp 1712256841
transform 1 0 1804 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5167
timestamp 1712256841
transform 1 0 1820 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5168
timestamp 1712256841
transform 1 0 1820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5169
timestamp 1712256841
transform 1 0 1740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5170
timestamp 1712256841
transform 1 0 1684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5171
timestamp 1712256841
transform 1 0 1788 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5172
timestamp 1712256841
transform 1 0 1740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1712256841
transform 1 0 1844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5174
timestamp 1712256841
transform 1 0 1788 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5175
timestamp 1712256841
transform 1 0 1756 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5176
timestamp 1712256841
transform 1 0 1860 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5177
timestamp 1712256841
transform 1 0 1852 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5178
timestamp 1712256841
transform 1 0 1836 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5179
timestamp 1712256841
transform 1 0 1820 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5180
timestamp 1712256841
transform 1 0 1820 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5181
timestamp 1712256841
transform 1 0 1772 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5182
timestamp 1712256841
transform 1 0 1932 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5183
timestamp 1712256841
transform 1 0 1724 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1712256841
transform 1 0 1892 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5185
timestamp 1712256841
transform 1 0 1892 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1712256841
transform 1 0 1812 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5187
timestamp 1712256841
transform 1 0 1796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1712256841
transform 1 0 1836 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5189
timestamp 1712256841
transform 1 0 1828 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5190
timestamp 1712256841
transform 1 0 1868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5191
timestamp 1712256841
transform 1 0 1844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5192
timestamp 1712256841
transform 1 0 2980 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5193
timestamp 1712256841
transform 1 0 2892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5194
timestamp 1712256841
transform 1 0 2876 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5195
timestamp 1712256841
transform 1 0 2820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5196
timestamp 1712256841
transform 1 0 2692 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5197
timestamp 1712256841
transform 1 0 2644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5198
timestamp 1712256841
transform 1 0 2068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5199
timestamp 1712256841
transform 1 0 1884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1712256841
transform 1 0 1700 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5201
timestamp 1712256841
transform 1 0 1748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5202
timestamp 1712256841
transform 1 0 1748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5203
timestamp 1712256841
transform 1 0 2876 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5204
timestamp 1712256841
transform 1 0 2740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5205
timestamp 1712256841
transform 1 0 2724 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_5206
timestamp 1712256841
transform 1 0 2628 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5207
timestamp 1712256841
transform 1 0 2596 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5208
timestamp 1712256841
transform 1 0 2516 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5209
timestamp 1712256841
transform 1 0 2508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1712256841
transform 1 0 2028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5211
timestamp 1712256841
transform 1 0 1788 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5212
timestamp 1712256841
transform 1 0 1716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5213
timestamp 1712256841
transform 1 0 1444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5214
timestamp 1712256841
transform 1 0 1348 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5215
timestamp 1712256841
transform 1 0 2084 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1712256841
transform 1 0 1980 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1712256841
transform 1 0 1908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1712256841
transform 1 0 1900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5219
timestamp 1712256841
transform 1 0 1940 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5220
timestamp 1712256841
transform 1 0 1940 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5221
timestamp 1712256841
transform 1 0 2004 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5222
timestamp 1712256841
transform 1 0 1956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5223
timestamp 1712256841
transform 1 0 1972 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5224
timestamp 1712256841
transform 1 0 1916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1712256841
transform 1 0 2340 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1712256841
transform 1 0 2164 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1712256841
transform 1 0 2244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1712256841
transform 1 0 2212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5229
timestamp 1712256841
transform 1 0 2052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5230
timestamp 1712256841
transform 1 0 2044 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1712256841
transform 1 0 1884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5232
timestamp 1712256841
transform 1 0 1828 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5233
timestamp 1712256841
transform 1 0 1908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1712256841
transform 1 0 1884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5235
timestamp 1712256841
transform 1 0 2068 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5236
timestamp 1712256841
transform 1 0 1940 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1712256841
transform 1 0 2124 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5238
timestamp 1712256841
transform 1 0 2108 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1712256841
transform 1 0 2092 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1712256841
transform 1 0 2092 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5241
timestamp 1712256841
transform 1 0 2228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1712256841
transform 1 0 2140 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1712256841
transform 1 0 2236 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5244
timestamp 1712256841
transform 1 0 2236 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1712256841
transform 1 0 2444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5246
timestamp 1712256841
transform 1 0 2180 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_5247
timestamp 1712256841
transform 1 0 3068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1712256841
transform 1 0 3004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1712256841
transform 1 0 2820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5250
timestamp 1712256841
transform 1 0 2708 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1712256841
transform 1 0 2492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1712256841
transform 1 0 2420 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5253
timestamp 1712256841
transform 1 0 2196 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5254
timestamp 1712256841
transform 1 0 2140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1712256841
transform 1 0 2444 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5256
timestamp 1712256841
transform 1 0 2236 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5257
timestamp 1712256841
transform 1 0 2180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5258
timestamp 1712256841
transform 1 0 2140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1712256841
transform 1 0 2244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5260
timestamp 1712256841
transform 1 0 2188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5261
timestamp 1712256841
transform 1 0 2260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5262
timestamp 1712256841
transform 1 0 2252 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5263
timestamp 1712256841
transform 1 0 2276 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1712256841
transform 1 0 2220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5265
timestamp 1712256841
transform 1 0 2452 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1712256841
transform 1 0 2236 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1712256841
transform 1 0 2380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5268
timestamp 1712256841
transform 1 0 2300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1712256841
transform 1 0 2300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5270
timestamp 1712256841
transform 1 0 2164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5271
timestamp 1712256841
transform 1 0 2148 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1712256841
transform 1 0 2188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5273
timestamp 1712256841
transform 1 0 2164 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1712256841
transform 1 0 2340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5275
timestamp 1712256841
transform 1 0 2300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5276
timestamp 1712256841
transform 1 0 2380 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5277
timestamp 1712256841
transform 1 0 2364 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5278
timestamp 1712256841
transform 1 0 2372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1712256841
transform 1 0 2260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1712256841
transform 1 0 2420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5281
timestamp 1712256841
transform 1 0 2340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5282
timestamp 1712256841
transform 1 0 2476 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1712256841
transform 1 0 2404 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5284
timestamp 1712256841
transform 1 0 2476 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5285
timestamp 1712256841
transform 1 0 2460 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1712256841
transform 1 0 2812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5287
timestamp 1712256841
transform 1 0 2748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5288
timestamp 1712256841
transform 1 0 2524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1712256841
transform 1 0 2492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1712256841
transform 1 0 2476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1712256841
transform 1 0 2420 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5292
timestamp 1712256841
transform 1 0 2404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5293
timestamp 1712256841
transform 1 0 2508 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5294
timestamp 1712256841
transform 1 0 2412 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1712256841
transform 1 0 2388 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1712256841
transform 1 0 2364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5297
timestamp 1712256841
transform 1 0 2364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5298
timestamp 1712256841
transform 1 0 2364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1712256841
transform 1 0 2364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5300
timestamp 1712256841
transform 1 0 2356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1712256841
transform 1 0 2372 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5302
timestamp 1712256841
transform 1 0 2332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5303
timestamp 1712256841
transform 1 0 2932 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5304
timestamp 1712256841
transform 1 0 2916 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1712256841
transform 1 0 2692 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1712256841
transform 1 0 2692 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_5307
timestamp 1712256841
transform 1 0 2524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1712256841
transform 1 0 2460 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5309
timestamp 1712256841
transform 1 0 2452 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5310
timestamp 1712256841
transform 1 0 2436 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5311
timestamp 1712256841
transform 1 0 2404 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5312
timestamp 1712256841
transform 1 0 2684 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1712256841
transform 1 0 2452 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5314
timestamp 1712256841
transform 1 0 2604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5315
timestamp 1712256841
transform 1 0 2588 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1712256841
transform 1 0 2588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5317
timestamp 1712256841
transform 1 0 2572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5318
timestamp 1712256841
transform 1 0 2364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5319
timestamp 1712256841
transform 1 0 2308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5320
timestamp 1712256841
transform 1 0 2412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5321
timestamp 1712256841
transform 1 0 2388 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5322
timestamp 1712256841
transform 1 0 2588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5323
timestamp 1712256841
transform 1 0 2556 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5324
timestamp 1712256841
transform 1 0 2588 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5325
timestamp 1712256841
transform 1 0 2556 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5326
timestamp 1712256841
transform 1 0 2604 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5327
timestamp 1712256841
transform 1 0 2460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5328
timestamp 1712256841
transform 1 0 2564 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5329
timestamp 1712256841
transform 1 0 2564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5330
timestamp 1712256841
transform 1 0 2692 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5331
timestamp 1712256841
transform 1 0 2628 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1712256841
transform 1 0 2700 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5333
timestamp 1712256841
transform 1 0 2684 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5334
timestamp 1712256841
transform 1 0 2756 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1712256841
transform 1 0 2756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5336
timestamp 1712256841
transform 1 0 2740 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1712256841
transform 1 0 2636 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5338
timestamp 1712256841
transform 1 0 2564 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5339
timestamp 1712256841
transform 1 0 2524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5340
timestamp 1712256841
transform 1 0 2628 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1712256841
transform 1 0 2588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1712256841
transform 1 0 2540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5343
timestamp 1712256841
transform 1 0 2108 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5344
timestamp 1712256841
transform 1 0 2532 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1712256841
transform 1 0 2532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1712256841
transform 1 0 2540 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5347
timestamp 1712256841
transform 1 0 2492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5348
timestamp 1712256841
transform 1 0 2692 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5349
timestamp 1712256841
transform 1 0 2540 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5350
timestamp 1712256841
transform 1 0 2708 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1712256841
transform 1 0 2676 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1712256841
transform 1 0 2676 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5353
timestamp 1712256841
transform 1 0 2668 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5354
timestamp 1712256841
transform 1 0 2628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5355
timestamp 1712256841
transform 1 0 2572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5356
timestamp 1712256841
transform 1 0 2548 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5357
timestamp 1712256841
transform 1 0 2620 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5358
timestamp 1712256841
transform 1 0 2620 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5359
timestamp 1712256841
transform 1 0 2844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5360
timestamp 1712256841
transform 1 0 2716 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5361
timestamp 1712256841
transform 1 0 2716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5362
timestamp 1712256841
transform 1 0 2716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5363
timestamp 1712256841
transform 1 0 2676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5364
timestamp 1712256841
transform 1 0 2652 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1712256841
transform 1 0 2604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1712256841
transform 1 0 2092 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1712256841
transform 1 0 2084 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1712256841
transform 1 0 2100 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5369
timestamp 1712256841
transform 1 0 2028 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5370
timestamp 1712256841
transform 1 0 3316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1712256841
transform 1 0 3156 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5372
timestamp 1712256841
transform 1 0 3140 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5373
timestamp 1712256841
transform 1 0 2676 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5374
timestamp 1712256841
transform 1 0 2724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5375
timestamp 1712256841
transform 1 0 2540 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1712256841
transform 1 0 2044 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5377
timestamp 1712256841
transform 1 0 1980 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5378
timestamp 1712256841
transform 1 0 1980 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1712256841
transform 1 0 1668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5380
timestamp 1712256841
transform 1 0 1652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5381
timestamp 1712256841
transform 1 0 3196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5382
timestamp 1712256841
transform 1 0 3196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5383
timestamp 1712256841
transform 1 0 3132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5384
timestamp 1712256841
transform 1 0 3284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5385
timestamp 1712256841
transform 1 0 3196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5386
timestamp 1712256841
transform 1 0 3180 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5387
timestamp 1712256841
transform 1 0 3180 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1712256841
transform 1 0 2732 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5389
timestamp 1712256841
transform 1 0 2684 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5390
timestamp 1712256841
transform 1 0 2676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5391
timestamp 1712256841
transform 1 0 2668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5392
timestamp 1712256841
transform 1 0 2780 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5393
timestamp 1712256841
transform 1 0 2780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5394
timestamp 1712256841
transform 1 0 2748 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1712256841
transform 1 0 2748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5396
timestamp 1712256841
transform 1 0 2676 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5397
timestamp 1712256841
transform 1 0 2636 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5398
timestamp 1712256841
transform 1 0 2708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5399
timestamp 1712256841
transform 1 0 2708 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5400
timestamp 1712256841
transform 1 0 2676 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5401
timestamp 1712256841
transform 1 0 2668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5402
timestamp 1712256841
transform 1 0 2932 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5403
timestamp 1712256841
transform 1 0 2860 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5404
timestamp 1712256841
transform 1 0 2916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5405
timestamp 1712256841
transform 1 0 2900 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5406
timestamp 1712256841
transform 1 0 2996 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5407
timestamp 1712256841
transform 1 0 2908 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1712256841
transform 1 0 3020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1712256841
transform 1 0 3004 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1712256841
transform 1 0 3036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1712256841
transform 1 0 2996 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5412
timestamp 1712256841
transform 1 0 2972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5413
timestamp 1712256841
transform 1 0 2940 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5414
timestamp 1712256841
transform 1 0 3260 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5415
timestamp 1712256841
transform 1 0 3108 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_5416
timestamp 1712256841
transform 1 0 3076 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1712256841
transform 1 0 2956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5418
timestamp 1712256841
transform 1 0 2940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5419
timestamp 1712256841
transform 1 0 3036 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5420
timestamp 1712256841
transform 1 0 3036 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1712256841
transform 1 0 2996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5422
timestamp 1712256841
transform 1 0 2996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5423
timestamp 1712256841
transform 1 0 3044 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5424
timestamp 1712256841
transform 1 0 2980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5425
timestamp 1712256841
transform 1 0 2972 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1712256841
transform 1 0 2956 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5427
timestamp 1712256841
transform 1 0 2932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1712256841
transform 1 0 2908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5429
timestamp 1712256841
transform 1 0 3092 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5430
timestamp 1712256841
transform 1 0 3020 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5431
timestamp 1712256841
transform 1 0 3036 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5432
timestamp 1712256841
transform 1 0 2804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5433
timestamp 1712256841
transform 1 0 2636 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5434
timestamp 1712256841
transform 1 0 2628 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5435
timestamp 1712256841
transform 1 0 3092 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_5436
timestamp 1712256841
transform 1 0 2916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5437
timestamp 1712256841
transform 1 0 3012 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5438
timestamp 1712256841
transform 1 0 2996 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5439
timestamp 1712256841
transform 1 0 2940 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5440
timestamp 1712256841
transform 1 0 2940 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_5441
timestamp 1712256841
transform 1 0 2964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1712256841
transform 1 0 2932 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5443
timestamp 1712256841
transform 1 0 2988 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5444
timestamp 1712256841
transform 1 0 2924 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5445
timestamp 1712256841
transform 1 0 3092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5446
timestamp 1712256841
transform 1 0 2972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5447
timestamp 1712256841
transform 1 0 2860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5448
timestamp 1712256841
transform 1 0 2860 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1712256841
transform 1 0 2988 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1712256841
transform 1 0 2972 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5451
timestamp 1712256841
transform 1 0 3276 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5452
timestamp 1712256841
transform 1 0 3268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1712256841
transform 1 0 3236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1712256841
transform 1 0 2948 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5455
timestamp 1712256841
transform 1 0 2876 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1712256841
transform 1 0 2844 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1712256841
transform 1 0 2996 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5458
timestamp 1712256841
transform 1 0 2980 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1712256841
transform 1 0 3068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1712256841
transform 1 0 3036 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5461
timestamp 1712256841
transform 1 0 3164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5462
timestamp 1712256841
transform 1 0 3028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5463
timestamp 1712256841
transform 1 0 3100 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5464
timestamp 1712256841
transform 1 0 3052 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1712256841
transform 1 0 3172 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5466
timestamp 1712256841
transform 1 0 3100 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1712256841
transform 1 0 3116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5468
timestamp 1712256841
transform 1 0 3116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1712256841
transform 1 0 3108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5470
timestamp 1712256841
transform 1 0 3084 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5471
timestamp 1712256841
transform 1 0 2724 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1712256841
transform 1 0 2668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1712256841
transform 1 0 2604 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5474
timestamp 1712256841
transform 1 0 2604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1712256841
transform 1 0 2524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5476
timestamp 1712256841
transform 1 0 2524 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1712256841
transform 1 0 2524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5478
timestamp 1712256841
transform 1 0 2508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1712256841
transform 1 0 2476 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5480
timestamp 1712256841
transform 1 0 2476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1712256841
transform 1 0 2780 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1712256841
transform 1 0 2740 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5483
timestamp 1712256841
transform 1 0 3108 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1712256841
transform 1 0 3100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1712256841
transform 1 0 3084 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1712256841
transform 1 0 3084 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1712256841
transform 1 0 3060 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1712256841
transform 1 0 3060 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1712256841
transform 1 0 3068 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5490
timestamp 1712256841
transform 1 0 3052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5491
timestamp 1712256841
transform 1 0 3060 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5492
timestamp 1712256841
transform 1 0 2812 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5493
timestamp 1712256841
transform 1 0 2996 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1712256841
transform 1 0 2932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5495
timestamp 1712256841
transform 1 0 3108 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5496
timestamp 1712256841
transform 1 0 3028 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5497
timestamp 1712256841
transform 1 0 2964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1712256841
transform 1 0 2964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1712256841
transform 1 0 3164 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1712256841
transform 1 0 3084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5501
timestamp 1712256841
transform 1 0 3092 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5502
timestamp 1712256841
transform 1 0 3044 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1712256841
transform 1 0 2620 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1712256841
transform 1 0 2548 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5505
timestamp 1712256841
transform 1 0 3108 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5506
timestamp 1712256841
transform 1 0 3068 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5507
timestamp 1712256841
transform 1 0 3060 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_5508
timestamp 1712256841
transform 1 0 2916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1712256841
transform 1 0 3108 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5510
timestamp 1712256841
transform 1 0 3092 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1712256841
transform 1 0 2892 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5512
timestamp 1712256841
transform 1 0 2892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5513
timestamp 1712256841
transform 1 0 2884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5514
timestamp 1712256841
transform 1 0 2860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5515
timestamp 1712256841
transform 1 0 3036 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5516
timestamp 1712256841
transform 1 0 2868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1712256841
transform 1 0 3044 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5518
timestamp 1712256841
transform 1 0 3036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5519
timestamp 1712256841
transform 1 0 3004 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1712256841
transform 1 0 3004 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5521
timestamp 1712256841
transform 1 0 3060 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1712256841
transform 1 0 3012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5523
timestamp 1712256841
transform 1 0 2612 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1712256841
transform 1 0 2532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1712256841
transform 1 0 2996 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1712256841
transform 1 0 2972 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1712256841
transform 1 0 2956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1712256841
transform 1 0 2868 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1712256841
transform 1 0 3068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5530
timestamp 1712256841
transform 1 0 2924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1712256841
transform 1 0 2844 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5532
timestamp 1712256841
transform 1 0 3172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5533
timestamp 1712256841
transform 1 0 2884 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1712256841
transform 1 0 2868 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5535
timestamp 1712256841
transform 1 0 2908 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5536
timestamp 1712256841
transform 1 0 2852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5537
timestamp 1712256841
transform 1 0 2876 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1712256841
transform 1 0 2748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5539
timestamp 1712256841
transform 1 0 2788 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5540
timestamp 1712256841
transform 1 0 2748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5541
timestamp 1712256841
transform 1 0 2908 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5542
timestamp 1712256841
transform 1 0 2852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1712256841
transform 1 0 2868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5544
timestamp 1712256841
transform 1 0 2868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5545
timestamp 1712256841
transform 1 0 2844 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1712256841
transform 1 0 2804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5547
timestamp 1712256841
transform 1 0 2860 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5548
timestamp 1712256841
transform 1 0 2852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5549
timestamp 1712256841
transform 1 0 2916 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5550
timestamp 1712256841
transform 1 0 2836 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5551
timestamp 1712256841
transform 1 0 2716 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5552
timestamp 1712256841
transform 1 0 2620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1712256841
transform 1 0 2876 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5554
timestamp 1712256841
transform 1 0 2844 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5555
timestamp 1712256841
transform 1 0 2908 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5556
timestamp 1712256841
transform 1 0 2844 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5557
timestamp 1712256841
transform 1 0 2844 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5558
timestamp 1712256841
transform 1 0 2828 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5559
timestamp 1712256841
transform 1 0 2772 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1712256841
transform 1 0 2740 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5561
timestamp 1712256841
transform 1 0 2788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5562
timestamp 1712256841
transform 1 0 2748 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5563
timestamp 1712256841
transform 1 0 2740 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5564
timestamp 1712256841
transform 1 0 2732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5565
timestamp 1712256841
transform 1 0 2884 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5566
timestamp 1712256841
transform 1 0 2732 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5567
timestamp 1712256841
transform 1 0 2900 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5568
timestamp 1712256841
transform 1 0 2852 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5569
timestamp 1712256841
transform 1 0 2924 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1712256841
transform 1 0 2868 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5571
timestamp 1712256841
transform 1 0 3236 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5572
timestamp 1712256841
transform 1 0 3228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5573
timestamp 1712256841
transform 1 0 3204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5574
timestamp 1712256841
transform 1 0 2732 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5575
timestamp 1712256841
transform 1 0 2604 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5576
timestamp 1712256841
transform 1 0 2900 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1712256841
transform 1 0 2772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5578
timestamp 1712256841
transform 1 0 2780 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5579
timestamp 1712256841
transform 1 0 2756 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5580
timestamp 1712256841
transform 1 0 2820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5581
timestamp 1712256841
transform 1 0 2636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5582
timestamp 1712256841
transform 1 0 2628 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5583
timestamp 1712256841
transform 1 0 2628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5584
timestamp 1712256841
transform 1 0 2820 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5585
timestamp 1712256841
transform 1 0 2788 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5586
timestamp 1712256841
transform 1 0 2756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5587
timestamp 1712256841
transform 1 0 2748 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5588
timestamp 1712256841
transform 1 0 2740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1712256841
transform 1 0 2828 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5590
timestamp 1712256841
transform 1 0 2812 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5591
timestamp 1712256841
transform 1 0 2764 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5592
timestamp 1712256841
transform 1 0 2764 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5593
timestamp 1712256841
transform 1 0 2788 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5594
timestamp 1712256841
transform 1 0 2756 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5595
timestamp 1712256841
transform 1 0 2772 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5596
timestamp 1712256841
transform 1 0 2748 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5597
timestamp 1712256841
transform 1 0 2772 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1712256841
transform 1 0 2740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5599
timestamp 1712256841
transform 1 0 2684 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5600
timestamp 1712256841
transform 1 0 2492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5601
timestamp 1712256841
transform 1 0 2588 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5602
timestamp 1712256841
transform 1 0 2540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5603
timestamp 1712256841
transform 1 0 2652 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5604
timestamp 1712256841
transform 1 0 2644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1712256841
transform 1 0 3244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5606
timestamp 1712256841
transform 1 0 3212 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5607
timestamp 1712256841
transform 1 0 3188 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5608
timestamp 1712256841
transform 1 0 3164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5609
timestamp 1712256841
transform 1 0 3164 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5610
timestamp 1712256841
transform 1 0 3356 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5611
timestamp 1712256841
transform 1 0 3332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5612
timestamp 1712256841
transform 1 0 2780 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5613
timestamp 1712256841
transform 1 0 2740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1712256841
transform 1 0 2932 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1712256841
transform 1 0 2932 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5616
timestamp 1712256841
transform 1 0 3108 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5617
timestamp 1712256841
transform 1 0 3068 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5618
timestamp 1712256841
transform 1 0 3212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5619
timestamp 1712256841
transform 1 0 3204 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5620
timestamp 1712256841
transform 1 0 3180 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5621
timestamp 1712256841
transform 1 0 3092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5622
timestamp 1712256841
transform 1 0 3332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5623
timestamp 1712256841
transform 1 0 3196 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_5624
timestamp 1712256841
transform 1 0 3436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1712256841
transform 1 0 3324 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_5626
timestamp 1712256841
transform 1 0 3340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1712256841
transform 1 0 3324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5628
timestamp 1712256841
transform 1 0 3076 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5629
timestamp 1712256841
transform 1 0 2892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5630
timestamp 1712256841
transform 1 0 3404 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5631
timestamp 1712256841
transform 1 0 3364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1712256841
transform 1 0 3292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1712256841
transform 1 0 3276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5634
timestamp 1712256841
transform 1 0 3268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5635
timestamp 1712256841
transform 1 0 3244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5636
timestamp 1712256841
transform 1 0 3244 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5637
timestamp 1712256841
transform 1 0 3340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5638
timestamp 1712256841
transform 1 0 3340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5639
timestamp 1712256841
transform 1 0 3332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1712256841
transform 1 0 3316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1712256841
transform 1 0 3316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5642
timestamp 1712256841
transform 1 0 3396 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5643
timestamp 1712256841
transform 1 0 3372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1712256841
transform 1 0 3348 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5645
timestamp 1712256841
transform 1 0 3324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1712256841
transform 1 0 3324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1712256841
transform 1 0 3428 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1712256841
transform 1 0 3396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5649
timestamp 1712256841
transform 1 0 3412 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5650
timestamp 1712256841
transform 1 0 3404 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1712256841
transform 1 0 3404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1712256841
transform 1 0 2964 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5653
timestamp 1712256841
transform 1 0 2924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5654
timestamp 1712256841
transform 1 0 3348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5655
timestamp 1712256841
transform 1 0 3308 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5656
timestamp 1712256841
transform 1 0 3308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1712256841
transform 1 0 3140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1712256841
transform 1 0 2956 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1712256841
transform 1 0 2916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1712256841
transform 1 0 3412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5661
timestamp 1712256841
transform 1 0 3348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1712256841
transform 1 0 3292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5663
timestamp 1712256841
transform 1 0 3180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5664
timestamp 1712256841
transform 1 0 2996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5665
timestamp 1712256841
transform 1 0 2964 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1712256841
transform 1 0 3044 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1712256841
transform 1 0 2988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5668
timestamp 1712256841
transform 1 0 3172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5669
timestamp 1712256841
transform 1 0 3148 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5670
timestamp 1712256841
transform 1 0 3340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5671
timestamp 1712256841
transform 1 0 3300 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1712256841
transform 1 0 3428 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5673
timestamp 1712256841
transform 1 0 3388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1712256841
transform 1 0 3244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5675
timestamp 1712256841
transform 1 0 3228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1712256841
transform 1 0 3180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5677
timestamp 1712256841
transform 1 0 3356 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5678
timestamp 1712256841
transform 1 0 3300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5679
timestamp 1712256841
transform 1 0 3300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5680
timestamp 1712256841
transform 1 0 3348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1712256841
transform 1 0 3348 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1712256841
transform 1 0 3228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5683
timestamp 1712256841
transform 1 0 3260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5684
timestamp 1712256841
transform 1 0 3236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5685
timestamp 1712256841
transform 1 0 3396 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5686
timestamp 1712256841
transform 1 0 3340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5687
timestamp 1712256841
transform 1 0 3340 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5688
timestamp 1712256841
transform 1 0 3316 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5689
timestamp 1712256841
transform 1 0 3316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1712256841
transform 1 0 3428 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5691
timestamp 1712256841
transform 1 0 3428 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1712256841
transform 1 0 3412 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1712256841
transform 1 0 3412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1712256841
transform 1 0 3412 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1712256841
transform 1 0 3388 0 1 1045
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1712256841
transform 1 0 3388 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_5697
timestamp 1712256841
transform 1 0 3252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5698
timestamp 1712256841
transform 1 0 3276 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5699
timestamp 1712256841
transform 1 0 3268 0 1 1085
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1712256841
transform 1 0 3228 0 1 1085
box -2 -2 2 2
use M2_M1  M2_M1_5701
timestamp 1712256841
transform 1 0 3228 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5702
timestamp 1712256841
transform 1 0 3300 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_5703
timestamp 1712256841
transform 1 0 3244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5704
timestamp 1712256841
transform 1 0 3244 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_5705
timestamp 1712256841
transform 1 0 3196 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5706
timestamp 1712256841
transform 1 0 3132 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1712256841
transform 1 0 3156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5708
timestamp 1712256841
transform 1 0 3140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5709
timestamp 1712256841
transform 1 0 3212 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5710
timestamp 1712256841
transform 1 0 3180 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5711
timestamp 1712256841
transform 1 0 3268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1712256841
transform 1 0 3188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5713
timestamp 1712256841
transform 1 0 3196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5714
timestamp 1712256841
transform 1 0 3052 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5715
timestamp 1712256841
transform 1 0 3052 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5716
timestamp 1712256841
transform 1 0 2948 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5717
timestamp 1712256841
transform 1 0 2932 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5718
timestamp 1712256841
transform 1 0 2716 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5719
timestamp 1712256841
transform 1 0 2716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5720
timestamp 1712256841
transform 1 0 2956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1712256841
transform 1 0 2940 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5722
timestamp 1712256841
transform 1 0 2980 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5723
timestamp 1712256841
transform 1 0 2948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5724
timestamp 1712256841
transform 1 0 2804 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5725
timestamp 1712256841
transform 1 0 2804 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5726
timestamp 1712256841
transform 1 0 2572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5727
timestamp 1712256841
transform 1 0 2572 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5728
timestamp 1712256841
transform 1 0 2684 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5729
timestamp 1712256841
transform 1 0 2684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5730
timestamp 1712256841
transform 1 0 2604 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5731
timestamp 1712256841
transform 1 0 2468 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5732
timestamp 1712256841
transform 1 0 2356 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5733
timestamp 1712256841
transform 1 0 2316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5734
timestamp 1712256841
transform 1 0 1988 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5735
timestamp 1712256841
transform 1 0 1964 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5736
timestamp 1712256841
transform 1 0 2252 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5737
timestamp 1712256841
transform 1 0 2252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5738
timestamp 1712256841
transform 1 0 2140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5739
timestamp 1712256841
transform 1 0 2100 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5740
timestamp 1712256841
transform 1 0 2092 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5741
timestamp 1712256841
transform 1 0 2052 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5742
timestamp 1712256841
transform 1 0 1884 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5743
timestamp 1712256841
transform 1 0 1860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5744
timestamp 1712256841
transform 1 0 1892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5745
timestamp 1712256841
transform 1 0 1804 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5746
timestamp 1712256841
transform 1 0 1732 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5747
timestamp 1712256841
transform 1 0 1684 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5748
timestamp 1712256841
transform 1 0 1572 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5749
timestamp 1712256841
transform 1 0 1572 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5750
timestamp 1712256841
transform 1 0 1484 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5751
timestamp 1712256841
transform 1 0 1484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5752
timestamp 1712256841
transform 1 0 1404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5753
timestamp 1712256841
transform 1 0 1380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5754
timestamp 1712256841
transform 1 0 1252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5755
timestamp 1712256841
transform 1 0 1244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5756
timestamp 1712256841
transform 1 0 1148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1712256841
transform 1 0 1044 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5758
timestamp 1712256841
transform 1 0 1068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5759
timestamp 1712256841
transform 1 0 940 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5760
timestamp 1712256841
transform 1 0 172 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5761
timestamp 1712256841
transform 1 0 156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5762
timestamp 1712256841
transform 1 0 108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5763
timestamp 1712256841
transform 1 0 108 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5764
timestamp 1712256841
transform 1 0 220 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5765
timestamp 1712256841
transform 1 0 220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5766
timestamp 1712256841
transform 1 0 332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5767
timestamp 1712256841
transform 1 0 332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5768
timestamp 1712256841
transform 1 0 444 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5769
timestamp 1712256841
transform 1 0 348 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5770
timestamp 1712256841
transform 1 0 444 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5771
timestamp 1712256841
transform 1 0 436 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5772
timestamp 1712256841
transform 1 0 460 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5773
timestamp 1712256841
transform 1 0 460 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5774
timestamp 1712256841
transform 1 0 604 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5775
timestamp 1712256841
transform 1 0 604 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5776
timestamp 1712256841
transform 1 0 700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5777
timestamp 1712256841
transform 1 0 548 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5778
timestamp 1712256841
transform 1 0 836 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5779
timestamp 1712256841
transform 1 0 836 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5780
timestamp 1712256841
transform 1 0 1140 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5781
timestamp 1712256841
transform 1 0 1140 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5782
timestamp 1712256841
transform 1 0 3076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5783
timestamp 1712256841
transform 1 0 3076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1712256841
transform 1 0 3044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5785
timestamp 1712256841
transform 1 0 3028 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5786
timestamp 1712256841
transform 1 0 3044 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5787
timestamp 1712256841
transform 1 0 3044 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5788
timestamp 1712256841
transform 1 0 3180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5789
timestamp 1712256841
transform 1 0 2972 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1712256841
transform 1 0 2940 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5791
timestamp 1712256841
transform 1 0 2996 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5792
timestamp 1712256841
transform 1 0 2972 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5793
timestamp 1712256841
transform 1 0 2916 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5794
timestamp 1712256841
transform 1 0 2796 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5795
timestamp 1712256841
transform 1 0 2972 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5796
timestamp 1712256841
transform 1 0 2940 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5797
timestamp 1712256841
transform 1 0 2884 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1712256841
transform 1 0 2876 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5799
timestamp 1712256841
transform 1 0 2788 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5800
timestamp 1712256841
transform 1 0 2764 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5801
timestamp 1712256841
transform 1 0 2788 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1712256841
transform 1 0 2764 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1712256841
transform 1 0 2740 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5804
timestamp 1712256841
transform 1 0 2428 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5805
timestamp 1712256841
transform 1 0 2284 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5806
timestamp 1712256841
transform 1 0 2180 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5807
timestamp 1712256841
transform 1 0 2132 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5808
timestamp 1712256841
transform 1 0 2044 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5809
timestamp 1712256841
transform 1 0 2140 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5810
timestamp 1712256841
transform 1 0 1300 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5811
timestamp 1712256841
transform 1 0 2332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1712256841
transform 1 0 2180 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5813
timestamp 1712256841
transform 1 0 1852 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5814
timestamp 1712256841
transform 1 0 1644 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5815
timestamp 1712256841
transform 1 0 1364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1712256841
transform 1 0 1252 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5817
timestamp 1712256841
transform 1 0 1068 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5818
timestamp 1712256841
transform 1 0 1292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5819
timestamp 1712256841
transform 1 0 1188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5820
timestamp 1712256841
transform 1 0 948 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5821
timestamp 1712256841
transform 1 0 932 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5822
timestamp 1712256841
transform 1 0 868 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5823
timestamp 1712256841
transform 1 0 1316 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5824
timestamp 1712256841
transform 1 0 1220 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5825
timestamp 1712256841
transform 1 0 1356 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5826
timestamp 1712256841
transform 1 0 1308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5827
timestamp 1712256841
transform 1 0 972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5828
timestamp 1712256841
transform 1 0 804 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5829
timestamp 1712256841
transform 1 0 772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5830
timestamp 1712256841
transform 1 0 732 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5831
timestamp 1712256841
transform 1 0 1996 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5832
timestamp 1712256841
transform 1 0 1972 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5833
timestamp 1712256841
transform 1 0 1764 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5834
timestamp 1712256841
transform 1 0 2004 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5835
timestamp 1712256841
transform 1 0 1972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5836
timestamp 1712256841
transform 1 0 1924 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_5837
timestamp 1712256841
transform 1 0 1844 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5838
timestamp 1712256841
transform 1 0 1556 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5839
timestamp 1712256841
transform 1 0 1508 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5840
timestamp 1712256841
transform 1 0 1476 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5841
timestamp 1712256841
transform 1 0 2076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5842
timestamp 1712256841
transform 1 0 2052 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1712256841
transform 1 0 2108 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5844
timestamp 1712256841
transform 1 0 2052 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5845
timestamp 1712256841
transform 1 0 2452 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5846
timestamp 1712256841
transform 1 0 2364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5847
timestamp 1712256841
transform 1 0 2060 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1712256841
transform 1 0 2036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5849
timestamp 1712256841
transform 1 0 1956 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5850
timestamp 1712256841
transform 1 0 3164 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5851
timestamp 1712256841
transform 1 0 3068 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5852
timestamp 1712256841
transform 1 0 3020 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_5853
timestamp 1712256841
transform 1 0 2556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5854
timestamp 1712256841
transform 1 0 2532 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5855
timestamp 1712256841
transform 1 0 2460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1712256841
transform 1 0 2380 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5857
timestamp 1712256841
transform 1 0 3052 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5858
timestamp 1712256841
transform 1 0 2852 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5859
timestamp 1712256841
transform 1 0 972 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5860
timestamp 1712256841
transform 1 0 860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5861
timestamp 1712256841
transform 1 0 620 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5862
timestamp 1712256841
transform 1 0 500 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5863
timestamp 1712256841
transform 1 0 468 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1712256841
transform 1 0 436 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5865
timestamp 1712256841
transform 1 0 348 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5866
timestamp 1712256841
transform 1 0 284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5867
timestamp 1712256841
transform 1 0 276 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5868
timestamp 1712256841
transform 1 0 260 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5869
timestamp 1712256841
transform 1 0 228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5870
timestamp 1712256841
transform 1 0 196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5871
timestamp 1712256841
transform 1 0 2916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5872
timestamp 1712256841
transform 1 0 2868 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5873
timestamp 1712256841
transform 1 0 2868 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5874
timestamp 1712256841
transform 1 0 2764 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5875
timestamp 1712256841
transform 1 0 2644 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5876
timestamp 1712256841
transform 1 0 3092 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5877
timestamp 1712256841
transform 1 0 3092 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1712256841
transform 1 0 3076 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5879
timestamp 1712256841
transform 1 0 3148 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5880
timestamp 1712256841
transform 1 0 3124 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1712256841
transform 1 0 3060 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5882
timestamp 1712256841
transform 1 0 2972 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1712256841
transform 1 0 3068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1712256841
transform 1 0 3020 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1712256841
transform 1 0 2556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5886
timestamp 1712256841
transform 1 0 2540 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1712256841
transform 1 0 2636 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5888
timestamp 1712256841
transform 1 0 2572 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5889
timestamp 1712256841
transform 1 0 2540 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5890
timestamp 1712256841
transform 1 0 2484 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5891
timestamp 1712256841
transform 1 0 2420 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5892
timestamp 1712256841
transform 1 0 2900 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5893
timestamp 1712256841
transform 1 0 2796 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5894
timestamp 1712256841
transform 1 0 2748 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5895
timestamp 1712256841
transform 1 0 2692 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5896
timestamp 1712256841
transform 1 0 2716 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5897
timestamp 1712256841
transform 1 0 2596 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5898
timestamp 1712256841
transform 1 0 2556 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5899
timestamp 1712256841
transform 1 0 2556 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_5900
timestamp 1712256841
transform 1 0 2532 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1712256841
transform 1 0 2508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5902
timestamp 1712256841
transform 1 0 2524 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5903
timestamp 1712256841
transform 1 0 2492 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5904
timestamp 1712256841
transform 1 0 2476 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5905
timestamp 1712256841
transform 1 0 2212 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5906
timestamp 1712256841
transform 1 0 2772 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5907
timestamp 1712256841
transform 1 0 2684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5908
timestamp 1712256841
transform 1 0 2652 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_5909
timestamp 1712256841
transform 1 0 2628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5910
timestamp 1712256841
transform 1 0 2604 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5911
timestamp 1712256841
transform 1 0 2524 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5912
timestamp 1712256841
transform 1 0 2412 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1712256841
transform 1 0 2412 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_5914
timestamp 1712256841
transform 1 0 2428 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5915
timestamp 1712256841
transform 1 0 2396 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1712256841
transform 1 0 2180 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5917
timestamp 1712256841
transform 1 0 2044 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5918
timestamp 1712256841
transform 1 0 1988 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5919
timestamp 1712256841
transform 1 0 2372 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5920
timestamp 1712256841
transform 1 0 2332 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5921
timestamp 1712256841
transform 1 0 2276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5922
timestamp 1712256841
transform 1 0 2220 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5923
timestamp 1712256841
transform 1 0 2180 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5924
timestamp 1712256841
transform 1 0 2028 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1712256841
transform 1 0 2420 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5926
timestamp 1712256841
transform 1 0 2340 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1712256841
transform 1 0 2268 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5928
timestamp 1712256841
transform 1 0 2028 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5929
timestamp 1712256841
transform 1 0 2004 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1712256841
transform 1 0 2148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5931
timestamp 1712256841
transform 1 0 2020 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5932
timestamp 1712256841
transform 1 0 2260 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5933
timestamp 1712256841
transform 1 0 2236 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5934
timestamp 1712256841
transform 1 0 2116 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5935
timestamp 1712256841
transform 1 0 2084 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5936
timestamp 1712256841
transform 1 0 2060 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1712256841
transform 1 0 1916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5938
timestamp 1712256841
transform 1 0 2348 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5939
timestamp 1712256841
transform 1 0 2164 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5940
timestamp 1712256841
transform 1 0 2340 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5941
timestamp 1712256841
transform 1 0 2284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5942
timestamp 1712256841
transform 1 0 2236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5943
timestamp 1712256841
transform 1 0 2132 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5944
timestamp 1712256841
transform 1 0 1988 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1712256841
transform 1 0 2308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5946
timestamp 1712256841
transform 1 0 2236 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_5947
timestamp 1712256841
transform 1 0 2324 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1712256841
transform 1 0 2300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5949
timestamp 1712256841
transform 1 0 2324 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5950
timestamp 1712256841
transform 1 0 2324 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5951
timestamp 1712256841
transform 1 0 2228 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5952
timestamp 1712256841
transform 1 0 2180 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5953
timestamp 1712256841
transform 1 0 2260 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5954
timestamp 1712256841
transform 1 0 2220 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1712256841
transform 1 0 2268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5956
timestamp 1712256841
transform 1 0 2260 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5957
timestamp 1712256841
transform 1 0 2092 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5958
timestamp 1712256841
transform 1 0 2068 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_5959
timestamp 1712256841
transform 1 0 2124 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5960
timestamp 1712256841
transform 1 0 2084 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5961
timestamp 1712256841
transform 1 0 2172 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5962
timestamp 1712256841
transform 1 0 2148 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5963
timestamp 1712256841
transform 1 0 1964 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5964
timestamp 1712256841
transform 1 0 1932 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5965
timestamp 1712256841
transform 1 0 1884 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1712256841
transform 1 0 2020 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5967
timestamp 1712256841
transform 1 0 1868 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5968
timestamp 1712256841
transform 1 0 1852 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5969
timestamp 1712256841
transform 1 0 2228 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5970
timestamp 1712256841
transform 1 0 2116 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5971
timestamp 1712256841
transform 1 0 1932 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5972
timestamp 1712256841
transform 1 0 1916 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5973
timestamp 1712256841
transform 1 0 1908 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5974
timestamp 1712256841
transform 1 0 1980 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5975
timestamp 1712256841
transform 1 0 1924 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5976
timestamp 1712256841
transform 1 0 1836 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5977
timestamp 1712256841
transform 1 0 1780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5978
timestamp 1712256841
transform 1 0 1724 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5979
timestamp 1712256841
transform 1 0 1708 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5980
timestamp 1712256841
transform 1 0 1812 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5981
timestamp 1712256841
transform 1 0 1788 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5982
timestamp 1712256841
transform 1 0 1860 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5983
timestamp 1712256841
transform 1 0 1804 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5984
timestamp 1712256841
transform 1 0 1860 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1712256841
transform 1 0 1812 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5986
timestamp 1712256841
transform 1 0 1884 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_5987
timestamp 1712256841
transform 1 0 1868 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5988
timestamp 1712256841
transform 1 0 1772 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5989
timestamp 1712256841
transform 1 0 1668 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5990
timestamp 1712256841
transform 1 0 1660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1712256841
transform 1 0 1644 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_5992
timestamp 1712256841
transform 1 0 1916 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_5993
timestamp 1712256841
transform 1 0 1908 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5994
timestamp 1712256841
transform 1 0 1956 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5995
timestamp 1712256841
transform 1 0 1900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5996
timestamp 1712256841
transform 1 0 1964 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5997
timestamp 1712256841
transform 1 0 1916 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1712256841
transform 1 0 1668 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5999
timestamp 1712256841
transform 1 0 1660 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6000
timestamp 1712256841
transform 1 0 1756 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6001
timestamp 1712256841
transform 1 0 1660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6002
timestamp 1712256841
transform 1 0 1756 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6003
timestamp 1712256841
transform 1 0 1708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6004
timestamp 1712256841
transform 1 0 1612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6005
timestamp 1712256841
transform 1 0 1588 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6006
timestamp 1712256841
transform 1 0 1732 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6007
timestamp 1712256841
transform 1 0 1604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6008
timestamp 1712256841
transform 1 0 1756 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6009
timestamp 1712256841
transform 1 0 1708 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6010
timestamp 1712256841
transform 1 0 1964 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6011
timestamp 1712256841
transform 1 0 1836 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6012
timestamp 1712256841
transform 1 0 1828 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6013
timestamp 1712256841
transform 1 0 1804 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6014
timestamp 1712256841
transform 1 0 1828 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6015
timestamp 1712256841
transform 1 0 1652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6016
timestamp 1712256841
transform 1 0 1620 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6017
timestamp 1712256841
transform 1 0 1612 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6018
timestamp 1712256841
transform 1 0 1548 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6019
timestamp 1712256841
transform 1 0 1548 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6020
timestamp 1712256841
transform 1 0 1780 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6021
timestamp 1712256841
transform 1 0 1620 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6022
timestamp 1712256841
transform 1 0 1596 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6023
timestamp 1712256841
transform 1 0 1564 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6024
timestamp 1712256841
transform 1 0 1556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6025
timestamp 1712256841
transform 1 0 1524 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6026
timestamp 1712256841
transform 1 0 1516 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6027
timestamp 1712256841
transform 1 0 1460 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6028
timestamp 1712256841
transform 1 0 1452 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6029
timestamp 1712256841
transform 1 0 1548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6030
timestamp 1712256841
transform 1 0 1444 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6031
timestamp 1712256841
transform 1 0 1636 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6032
timestamp 1712256841
transform 1 0 1524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1712256841
transform 1 0 1420 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6034
timestamp 1712256841
transform 1 0 1412 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6035
timestamp 1712256841
transform 1 0 1380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6036
timestamp 1712256841
transform 1 0 1380 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6037
timestamp 1712256841
transform 1 0 1644 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1712256841
transform 1 0 1580 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6039
timestamp 1712256841
transform 1 0 1428 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6040
timestamp 1712256841
transform 1 0 1348 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1712256841
transform 1 0 1420 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1712256841
transform 1 0 1340 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6043
timestamp 1712256841
transform 1 0 1604 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6044
timestamp 1712256841
transform 1 0 1428 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6045
timestamp 1712256841
transform 1 0 1324 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6046
timestamp 1712256841
transform 1 0 1308 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6047
timestamp 1712256841
transform 1 0 1404 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6048
timestamp 1712256841
transform 1 0 1316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6049
timestamp 1712256841
transform 1 0 1612 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6050
timestamp 1712256841
transform 1 0 1404 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6051
timestamp 1712256841
transform 1 0 1252 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6052
timestamp 1712256841
transform 1 0 1244 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6053
timestamp 1712256841
transform 1 0 1436 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6054
timestamp 1712256841
transform 1 0 1236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6055
timestamp 1712256841
transform 1 0 1540 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6056
timestamp 1712256841
transform 1 0 1476 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6057
timestamp 1712256841
transform 1 0 1588 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6058
timestamp 1712256841
transform 1 0 1500 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6059
timestamp 1712256841
transform 1 0 1484 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6060
timestamp 1712256841
transform 1 0 1404 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1712256841
transform 1 0 1196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6062
timestamp 1712256841
transform 1 0 1172 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6063
timestamp 1712256841
transform 1 0 1092 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6064
timestamp 1712256841
transform 1 0 1092 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6065
timestamp 1712256841
transform 1 0 1092 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6066
timestamp 1712256841
transform 1 0 1220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6067
timestamp 1712256841
transform 1 0 1196 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6068
timestamp 1712256841
transform 1 0 1236 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6069
timestamp 1712256841
transform 1 0 1212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1712256841
transform 1 0 1236 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6071
timestamp 1712256841
transform 1 0 1188 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6072
timestamp 1712256841
transform 1 0 1428 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6073
timestamp 1712256841
transform 1 0 1148 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6074
timestamp 1712256841
transform 1 0 1148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6075
timestamp 1712256841
transform 1 0 1076 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6076
timestamp 1712256841
transform 1 0 1052 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6077
timestamp 1712256841
transform 1 0 1036 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6078
timestamp 1712256841
transform 1 0 1036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6079
timestamp 1712256841
transform 1 0 1020 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1712256841
transform 1 0 236 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1712256841
transform 1 0 1132 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6082
timestamp 1712256841
transform 1 0 1012 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6083
timestamp 1712256841
transform 1 0 1132 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6084
timestamp 1712256841
transform 1 0 1084 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6085
timestamp 1712256841
transform 1 0 628 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6086
timestamp 1712256841
transform 1 0 276 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6087
timestamp 1712256841
transform 1 0 1140 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6088
timestamp 1712256841
transform 1 0 620 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6089
timestamp 1712256841
transform 1 0 1164 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6090
timestamp 1712256841
transform 1 0 1140 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1712256841
transform 1 0 756 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6092
timestamp 1712256841
transform 1 0 324 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6093
timestamp 1712256841
transform 1 0 1012 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6094
timestamp 1712256841
transform 1 0 748 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6095
timestamp 1712256841
transform 1 0 1060 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6096
timestamp 1712256841
transform 1 0 1036 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6097
timestamp 1712256841
transform 1 0 1092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6098
timestamp 1712256841
transform 1 0 1076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6099
timestamp 1712256841
transform 1 0 1052 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6100
timestamp 1712256841
transform 1 0 1012 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6101
timestamp 1712256841
transform 1 0 996 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1712256841
transform 1 0 1100 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6103
timestamp 1712256841
transform 1 0 908 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1712256841
transform 1 0 732 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6105
timestamp 1712256841
transform 1 0 1140 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6106
timestamp 1712256841
transform 1 0 892 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6107
timestamp 1712256841
transform 1 0 604 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6108
timestamp 1712256841
transform 1 0 572 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6109
timestamp 1712256841
transform 1 0 564 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1712256841
transform 1 0 532 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6111
timestamp 1712256841
transform 1 0 604 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6112
timestamp 1712256841
transform 1 0 300 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6113
timestamp 1712256841
transform 1 0 628 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6114
timestamp 1712256841
transform 1 0 596 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6115
timestamp 1712256841
transform 1 0 740 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6116
timestamp 1712256841
transform 1 0 644 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6117
timestamp 1712256841
transform 1 0 996 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6118
timestamp 1712256841
transform 1 0 844 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6119
timestamp 1712256841
transform 1 0 804 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6120
timestamp 1712256841
transform 1 0 732 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1712256841
transform 1 0 676 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6122
timestamp 1712256841
transform 1 0 660 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6123
timestamp 1712256841
transform 1 0 628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6124
timestamp 1712256841
transform 1 0 532 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6125
timestamp 1712256841
transform 1 0 508 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6126
timestamp 1712256841
transform 1 0 596 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6127
timestamp 1712256841
transform 1 0 524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6128
timestamp 1712256841
transform 1 0 668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6129
timestamp 1712256841
transform 1 0 596 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6130
timestamp 1712256841
transform 1 0 524 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6131
timestamp 1712256841
transform 1 0 412 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1712256841
transform 1 0 556 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6133
timestamp 1712256841
transform 1 0 516 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6134
timestamp 1712256841
transform 1 0 636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6135
timestamp 1712256841
transform 1 0 556 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6136
timestamp 1712256841
transform 1 0 564 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6137
timestamp 1712256841
transform 1 0 500 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6138
timestamp 1712256841
transform 1 0 588 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6139
timestamp 1712256841
transform 1 0 556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6140
timestamp 1712256841
transform 1 0 684 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1712256841
transform 1 0 612 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6142
timestamp 1712256841
transform 1 0 884 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6143
timestamp 1712256841
transform 1 0 876 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6144
timestamp 1712256841
transform 1 0 876 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6145
timestamp 1712256841
transform 1 0 908 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6146
timestamp 1712256841
transform 1 0 860 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6147
timestamp 1712256841
transform 1 0 828 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6148
timestamp 1712256841
transform 1 0 828 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6149
timestamp 1712256841
transform 1 0 788 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6150
timestamp 1712256841
transform 1 0 788 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6151
timestamp 1712256841
transform 1 0 892 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6152
timestamp 1712256841
transform 1 0 828 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1712256841
transform 1 0 796 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6154
timestamp 1712256841
transform 1 0 796 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6155
timestamp 1712256841
transform 1 0 780 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6156
timestamp 1712256841
transform 1 0 756 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6157
timestamp 1712256841
transform 1 0 724 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6158
timestamp 1712256841
transform 1 0 740 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6159
timestamp 1712256841
transform 1 0 668 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6160
timestamp 1712256841
transform 1 0 836 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6161
timestamp 1712256841
transform 1 0 732 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6162
timestamp 1712256841
transform 1 0 956 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6163
timestamp 1712256841
transform 1 0 852 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6164
timestamp 1712256841
transform 1 0 836 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6165
timestamp 1712256841
transform 1 0 804 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6166
timestamp 1712256841
transform 1 0 692 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6167
timestamp 1712256841
transform 1 0 836 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6168
timestamp 1712256841
transform 1 0 812 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6169
timestamp 1712256841
transform 1 0 644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6170
timestamp 1712256841
transform 1 0 524 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1712256841
transform 1 0 716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6172
timestamp 1712256841
transform 1 0 636 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6173
timestamp 1712256841
transform 1 0 740 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6174
timestamp 1712256841
transform 1 0 716 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1712256841
transform 1 0 900 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6176
timestamp 1712256841
transform 1 0 900 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6177
timestamp 1712256841
transform 1 0 860 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6178
timestamp 1712256841
transform 1 0 804 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6179
timestamp 1712256841
transform 1 0 1044 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6180
timestamp 1712256841
transform 1 0 988 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6181
timestamp 1712256841
transform 1 0 996 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6182
timestamp 1712256841
transform 1 0 980 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6183
timestamp 1712256841
transform 1 0 996 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6184
timestamp 1712256841
transform 1 0 844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6185
timestamp 1712256841
transform 1 0 1204 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6186
timestamp 1712256841
transform 1 0 964 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6187
timestamp 1712256841
transform 1 0 964 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6188
timestamp 1712256841
transform 1 0 860 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6189
timestamp 1712256841
transform 1 0 772 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6190
timestamp 1712256841
transform 1 0 756 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6191
timestamp 1712256841
transform 1 0 1668 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6192
timestamp 1712256841
transform 1 0 1660 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6193
timestamp 1712256841
transform 1 0 1844 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6194
timestamp 1712256841
transform 1 0 1828 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6195
timestamp 1712256841
transform 1 0 1876 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6196
timestamp 1712256841
transform 1 0 1796 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6197
timestamp 1712256841
transform 1 0 1692 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6198
timestamp 1712256841
transform 1 0 1332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6199
timestamp 1712256841
transform 1 0 1948 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6200
timestamp 1712256841
transform 1 0 1908 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6201
timestamp 1712256841
transform 1 0 3116 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6202
timestamp 1712256841
transform 1 0 2964 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6203
timestamp 1712256841
transform 1 0 2828 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6204
timestamp 1712256841
transform 1 0 2676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6205
timestamp 1712256841
transform 1 0 2396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6206
timestamp 1712256841
transform 1 0 2236 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6207
timestamp 1712256841
transform 1 0 2068 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6208
timestamp 1712256841
transform 1 0 2044 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6209
timestamp 1712256841
transform 1 0 1844 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6210
timestamp 1712256841
transform 1 0 1116 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6211
timestamp 1712256841
transform 1 0 868 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6212
timestamp 1712256841
transform 1 0 636 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6213
timestamp 1712256841
transform 1 0 556 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6214
timestamp 1712256841
transform 1 0 484 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6215
timestamp 1712256841
transform 1 0 460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6216
timestamp 1712256841
transform 1 0 436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6217
timestamp 1712256841
transform 1 0 3108 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6218
timestamp 1712256841
transform 1 0 3092 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6219
timestamp 1712256841
transform 1 0 3212 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6220
timestamp 1712256841
transform 1 0 3172 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6221
timestamp 1712256841
transform 1 0 3148 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6222
timestamp 1712256841
transform 1 0 3116 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6223
timestamp 1712256841
transform 1 0 3100 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6224
timestamp 1712256841
transform 1 0 3084 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6225
timestamp 1712256841
transform 1 0 2844 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6226
timestamp 1712256841
transform 1 0 2628 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6227
timestamp 1712256841
transform 1 0 2428 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6228
timestamp 1712256841
transform 1 0 2300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6229
timestamp 1712256841
transform 1 0 2036 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6230
timestamp 1712256841
transform 1 0 1908 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6231
timestamp 1712256841
transform 1 0 1716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6232
timestamp 1712256841
transform 1 0 1588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6233
timestamp 1712256841
transform 1 0 1292 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6234
timestamp 1712256841
transform 1 0 2412 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6235
timestamp 1712256841
transform 1 0 2396 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6236
timestamp 1712256841
transform 1 0 1924 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6237
timestamp 1712256841
transform 1 0 1820 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1712256841
transform 1 0 716 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6239
timestamp 1712256841
transform 1 0 716 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6240
timestamp 1712256841
transform 1 0 932 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6241
timestamp 1712256841
transform 1 0 932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6242
timestamp 1712256841
transform 1 0 900 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6243
timestamp 1712256841
transform 1 0 900 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6244
timestamp 1712256841
transform 1 0 2156 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6245
timestamp 1712256841
transform 1 0 1956 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6246
timestamp 1712256841
transform 1 0 1276 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6247
timestamp 1712256841
transform 1 0 1244 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_6248
timestamp 1712256841
transform 1 0 1516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6249
timestamp 1712256841
transform 1 0 1500 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6250
timestamp 1712256841
transform 1 0 2220 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_6251
timestamp 1712256841
transform 1 0 2220 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6252
timestamp 1712256841
transform 1 0 3140 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6253
timestamp 1712256841
transform 1 0 3044 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6254
timestamp 1712256841
transform 1 0 2748 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6255
timestamp 1712256841
transform 1 0 2748 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6256
timestamp 1712256841
transform 1 0 3172 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6257
timestamp 1712256841
transform 1 0 3172 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6258
timestamp 1712256841
transform 1 0 2852 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6259
timestamp 1712256841
transform 1 0 2852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6260
timestamp 1712256841
transform 1 0 2620 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6261
timestamp 1712256841
transform 1 0 2540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6262
timestamp 1712256841
transform 1 0 2708 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6263
timestamp 1712256841
transform 1 0 2636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6264
timestamp 1712256841
transform 1 0 2764 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6265
timestamp 1712256841
transform 1 0 2764 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6266
timestamp 1712256841
transform 1 0 2500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1712256841
transform 1 0 2412 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6268
timestamp 1712256841
transform 1 0 2084 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6269
timestamp 1712256841
transform 1 0 2004 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6270
timestamp 1712256841
transform 1 0 2308 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6271
timestamp 1712256841
transform 1 0 2236 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6272
timestamp 1712256841
transform 1 0 2180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6273
timestamp 1712256841
transform 1 0 2164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6274
timestamp 1712256841
transform 1 0 2068 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6275
timestamp 1712256841
transform 1 0 1988 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6276
timestamp 1712256841
transform 1 0 1788 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6277
timestamp 1712256841
transform 1 0 1724 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1712256841
transform 1 0 1916 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6279
timestamp 1712256841
transform 1 0 1852 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6280
timestamp 1712256841
transform 1 0 1660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6281
timestamp 1712256841
transform 1 0 1636 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6282
timestamp 1712256841
transform 1 0 1564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6283
timestamp 1712256841
transform 1 0 1564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6284
timestamp 1712256841
transform 1 0 1460 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6285
timestamp 1712256841
transform 1 0 1396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6286
timestamp 1712256841
transform 1 0 1420 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6287
timestamp 1712256841
transform 1 0 1340 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6288
timestamp 1712256841
transform 1 0 1340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6289
timestamp 1712256841
transform 1 0 1308 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6290
timestamp 1712256841
transform 1 0 1252 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1712256841
transform 1 0 1164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6292
timestamp 1712256841
transform 1 0 1196 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6293
timestamp 1712256841
transform 1 0 1108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6294
timestamp 1712256841
transform 1 0 220 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6295
timestamp 1712256841
transform 1 0 140 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6296
timestamp 1712256841
transform 1 0 252 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6297
timestamp 1712256841
transform 1 0 140 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6298
timestamp 1712256841
transform 1 0 308 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6299
timestamp 1712256841
transform 1 0 220 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6300
timestamp 1712256841
transform 1 0 300 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6301
timestamp 1712256841
transform 1 0 300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6302
timestamp 1712256841
transform 1 0 492 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6303
timestamp 1712256841
transform 1 0 404 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1712256841
transform 1 0 372 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1712256841
transform 1 0 356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6306
timestamp 1712256841
transform 1 0 460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6307
timestamp 1712256841
transform 1 0 460 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6308
timestamp 1712256841
transform 1 0 668 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6309
timestamp 1712256841
transform 1 0 580 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6310
timestamp 1712256841
transform 1 0 524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6311
timestamp 1712256841
transform 1 0 420 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6312
timestamp 1712256841
transform 1 0 892 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6313
timestamp 1712256841
transform 1 0 788 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6314
timestamp 1712256841
transform 1 0 1044 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6315
timestamp 1712256841
transform 1 0 980 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6316
timestamp 1712256841
transform 1 0 3364 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6317
timestamp 1712256841
transform 1 0 3364 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6318
timestamp 1712256841
transform 1 0 3276 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6319
timestamp 1712256841
transform 1 0 3276 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6320
timestamp 1712256841
transform 1 0 3380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6321
timestamp 1712256841
transform 1 0 3316 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1712256841
transform 1 0 3412 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1712256841
transform 1 0 3372 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6324
timestamp 1712256841
transform 1 0 3420 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1712256841
transform 1 0 3420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1712256841
transform 1 0 3364 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6327
timestamp 1712256841
transform 1 0 3364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6328
timestamp 1712256841
transform 1 0 3364 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6329
timestamp 1712256841
transform 1 0 3316 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1712256841
transform 1 0 3092 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1712256841
transform 1 0 3092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6332
timestamp 1712256841
transform 1 0 3188 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6333
timestamp 1712256841
transform 1 0 3036 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6334
timestamp 1712256841
transform 1 0 3196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1712256841
transform 1 0 3076 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6336
timestamp 1712256841
transform 1 0 3268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6337
timestamp 1712256841
transform 1 0 3236 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6338
timestamp 1712256841
transform 1 0 3308 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1712256841
transform 1 0 3284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6340
timestamp 1712256841
transform 1 0 3404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6341
timestamp 1712256841
transform 1 0 3324 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6342
timestamp 1712256841
transform 1 0 3308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6343
timestamp 1712256841
transform 1 0 3308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6344
timestamp 1712256841
transform 1 0 3340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6345
timestamp 1712256841
transform 1 0 3244 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6346
timestamp 1712256841
transform 1 0 3164 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6347
timestamp 1712256841
transform 1 0 3164 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6348
timestamp 1712256841
transform 1 0 3356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6349
timestamp 1712256841
transform 1 0 3340 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_6350
timestamp 1712256841
transform 1 0 3340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6351
timestamp 1712256841
transform 1 0 3340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6352
timestamp 1712256841
transform 1 0 3332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6353
timestamp 1712256841
transform 1 0 3396 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6354
timestamp 1712256841
transform 1 0 3356 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6355
timestamp 1712256841
transform 1 0 3348 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6356
timestamp 1712256841
transform 1 0 3316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6357
timestamp 1712256841
transform 1 0 3364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6358
timestamp 1712256841
transform 1 0 3324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6359
timestamp 1712256841
transform 1 0 3324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6360
timestamp 1712256841
transform 1 0 3380 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1712256841
transform 1 0 3356 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6362
timestamp 1712256841
transform 1 0 3428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6363
timestamp 1712256841
transform 1 0 3428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1712256841
transform 1 0 3404 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6365
timestamp 1712256841
transform 1 0 3364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6366
timestamp 1712256841
transform 1 0 3428 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6367
timestamp 1712256841
transform 1 0 3396 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6368
timestamp 1712256841
transform 1 0 3348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6369
timestamp 1712256841
transform 1 0 3308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6370
timestamp 1712256841
transform 1 0 3308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6371
timestamp 1712256841
transform 1 0 3252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6372
timestamp 1712256841
transform 1 0 3212 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6373
timestamp 1712256841
transform 1 0 3068 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6374
timestamp 1712256841
transform 1 0 2940 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6375
timestamp 1712256841
transform 1 0 2884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6376
timestamp 1712256841
transform 1 0 2364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6377
timestamp 1712256841
transform 1 0 2332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6378
timestamp 1712256841
transform 1 0 2324 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6379
timestamp 1712256841
transform 1 0 2308 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1712256841
transform 1 0 2308 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6381
timestamp 1712256841
transform 1 0 2284 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6382
timestamp 1712256841
transform 1 0 3052 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6383
timestamp 1712256841
transform 1 0 2716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6384
timestamp 1712256841
transform 1 0 2556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6385
timestamp 1712256841
transform 1 0 2516 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1712256841
transform 1 0 2372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1712256841
transform 1 0 2212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6388
timestamp 1712256841
transform 1 0 2116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6389
timestamp 1712256841
transform 1 0 1812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6390
timestamp 1712256841
transform 1 0 1636 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6391
timestamp 1712256841
transform 1 0 1428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6392
timestamp 1712256841
transform 1 0 1060 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6393
timestamp 1712256841
transform 1 0 916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6394
timestamp 1712256841
transform 1 0 2124 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6395
timestamp 1712256841
transform 1 0 2044 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1712256841
transform 1 0 2028 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6397
timestamp 1712256841
transform 1 0 1996 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6398
timestamp 1712256841
transform 1 0 1996 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1712256841
transform 1 0 2204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6400
timestamp 1712256841
transform 1 0 2188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6401
timestamp 1712256841
transform 1 0 2076 0 1 2255
box -2 -2 2 2
use M2_M1  M2_M1_6402
timestamp 1712256841
transform 1 0 2076 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6403
timestamp 1712256841
transform 1 0 2060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6404
timestamp 1712256841
transform 1 0 2060 0 1 2255
box -2 -2 2 2
use M2_M1  M2_M1_6405
timestamp 1712256841
transform 1 0 1716 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6406
timestamp 1712256841
transform 1 0 2428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6407
timestamp 1712256841
transform 1 0 2420 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6408
timestamp 1712256841
transform 1 0 2396 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6409
timestamp 1712256841
transform 1 0 2396 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6410
timestamp 1712256841
transform 1 0 2380 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6411
timestamp 1712256841
transform 1 0 1740 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6412
timestamp 1712256841
transform 1 0 2508 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6413
timestamp 1712256841
transform 1 0 2500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6414
timestamp 1712256841
transform 1 0 2492 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6415
timestamp 1712256841
transform 1 0 2452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6416
timestamp 1712256841
transform 1 0 2356 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6417
timestamp 1712256841
transform 1 0 2228 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6418
timestamp 1712256841
transform 1 0 1940 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6419
timestamp 1712256841
transform 1 0 2636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6420
timestamp 1712256841
transform 1 0 2620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6421
timestamp 1712256841
transform 1 0 2612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6422
timestamp 1712256841
transform 1 0 2460 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6423
timestamp 1712256841
transform 1 0 2196 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6424
timestamp 1712256841
transform 1 0 1844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6425
timestamp 1712256841
transform 1 0 2860 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6426
timestamp 1712256841
transform 1 0 2828 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6427
timestamp 1712256841
transform 1 0 2828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6428
timestamp 1712256841
transform 1 0 2796 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6429
timestamp 1712256841
transform 1 0 2796 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6430
timestamp 1712256841
transform 1 0 2468 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6431
timestamp 1712256841
transform 1 0 2444 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6432
timestamp 1712256841
transform 1 0 1292 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6433
timestamp 1712256841
transform 1 0 1220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6434
timestamp 1712256841
transform 1 0 1196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6435
timestamp 1712256841
transform 1 0 1004 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6436
timestamp 1712256841
transform 1 0 972 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6437
timestamp 1712256841
transform 1 0 1044 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1712256841
transform 1 0 956 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6439
timestamp 1712256841
transform 1 0 844 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6440
timestamp 1712256841
transform 1 0 812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6441
timestamp 1712256841
transform 1 0 812 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6442
timestamp 1712256841
transform 1 0 3020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6443
timestamp 1712256841
transform 1 0 2980 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6444
timestamp 1712256841
transform 1 0 2932 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6445
timestamp 1712256841
transform 1 0 2876 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6446
timestamp 1712256841
transform 1 0 2852 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6447
timestamp 1712256841
transform 1 0 2852 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6448
timestamp 1712256841
transform 1 0 940 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1712256841
transform 1 0 852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6450
timestamp 1712256841
transform 1 0 732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6451
timestamp 1712256841
transform 1 0 724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6452
timestamp 1712256841
transform 1 0 684 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6453
timestamp 1712256841
transform 1 0 676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6454
timestamp 1712256841
transform 1 0 964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6455
timestamp 1712256841
transform 1 0 900 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_6456
timestamp 1712256841
transform 1 0 796 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6457
timestamp 1712256841
transform 1 0 780 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6458
timestamp 1712256841
transform 1 0 700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1712256841
transform 1 0 628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6460
timestamp 1712256841
transform 1 0 892 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6461
timestamp 1712256841
transform 1 0 676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6462
timestamp 1712256841
transform 1 0 532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6463
timestamp 1712256841
transform 1 0 476 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6464
timestamp 1712256841
transform 1 0 708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6465
timestamp 1712256841
transform 1 0 524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6466
timestamp 1712256841
transform 1 0 444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6467
timestamp 1712256841
transform 1 0 404 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6468
timestamp 1712256841
transform 1 0 620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6469
timestamp 1712256841
transform 1 0 524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6470
timestamp 1712256841
transform 1 0 380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6471
timestamp 1712256841
transform 1 0 348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6472
timestamp 1712256841
transform 1 0 684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6473
timestamp 1712256841
transform 1 0 564 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6474
timestamp 1712256841
transform 1 0 308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6475
timestamp 1712256841
transform 1 0 244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6476
timestamp 1712256841
transform 1 0 772 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6477
timestamp 1712256841
transform 1 0 772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6478
timestamp 1712256841
transform 1 0 572 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6479
timestamp 1712256841
transform 1 0 244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6480
timestamp 1712256841
transform 1 0 228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6481
timestamp 1712256841
transform 1 0 644 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6482
timestamp 1712256841
transform 1 0 644 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1712256841
transform 1 0 508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6484
timestamp 1712256841
transform 1 0 100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6485
timestamp 1712256841
transform 1 0 84 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_6486
timestamp 1712256841
transform 1 0 68 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6487
timestamp 1712256841
transform 1 0 68 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_6488
timestamp 1712256841
transform 1 0 932 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6489
timestamp 1712256841
transform 1 0 908 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6490
timestamp 1712256841
transform 1 0 732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6491
timestamp 1712256841
transform 1 0 564 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6492
timestamp 1712256841
transform 1 0 172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6493
timestamp 1712256841
transform 1 0 164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6494
timestamp 1712256841
transform 1 0 116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6495
timestamp 1712256841
transform 1 0 916 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6496
timestamp 1712256841
transform 1 0 876 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6497
timestamp 1712256841
transform 1 0 876 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6498
timestamp 1712256841
transform 1 0 804 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1712256841
transform 1 0 804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6500
timestamp 1712256841
transform 1 0 788 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_6501
timestamp 1712256841
transform 1 0 612 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6502
timestamp 1712256841
transform 1 0 596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6503
timestamp 1712256841
transform 1 0 564 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6504
timestamp 1712256841
transform 1 0 3044 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6505
timestamp 1712256841
transform 1 0 2876 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6506
timestamp 1712256841
transform 1 0 2876 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6507
timestamp 1712256841
transform 1 0 2876 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6508
timestamp 1712256841
transform 1 0 2844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6509
timestamp 1712256841
transform 1 0 2836 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6510
timestamp 1712256841
transform 1 0 2724 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6511
timestamp 1712256841
transform 1 0 2452 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6512
timestamp 1712256841
transform 1 0 2444 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6513
timestamp 1712256841
transform 1 0 1412 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6514
timestamp 1712256841
transform 1 0 1052 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6515
timestamp 1712256841
transform 1 0 1052 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_6516
timestamp 1712256841
transform 1 0 1052 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6517
timestamp 1712256841
transform 1 0 1036 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_6518
timestamp 1712256841
transform 1 0 1020 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_6519
timestamp 1712256841
transform 1 0 1020 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6520
timestamp 1712256841
transform 1 0 1012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6521
timestamp 1712256841
transform 1 0 988 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6522
timestamp 1712256841
transform 1 0 972 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6523
timestamp 1712256841
transform 1 0 1372 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6524
timestamp 1712256841
transform 1 0 1268 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6525
timestamp 1712256841
transform 1 0 1268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6526
timestamp 1712256841
transform 1 0 1164 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6527
timestamp 1712256841
transform 1 0 1164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6528
timestamp 1712256841
transform 1 0 1140 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6529
timestamp 1712256841
transform 1 0 1132 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6530
timestamp 1712256841
transform 1 0 1124 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6531
timestamp 1712256841
transform 1 0 1420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6532
timestamp 1712256841
transform 1 0 1372 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6533
timestamp 1712256841
transform 1 0 1372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6534
timestamp 1712256841
transform 1 0 1284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6535
timestamp 1712256841
transform 1 0 1260 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6536
timestamp 1712256841
transform 1 0 1220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6537
timestamp 1712256841
transform 1 0 1116 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6538
timestamp 1712256841
transform 1 0 1580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1712256841
transform 1 0 1532 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6540
timestamp 1712256841
transform 1 0 1476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6541
timestamp 1712256841
transform 1 0 1428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6542
timestamp 1712256841
transform 1 0 1284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1712256841
transform 1 0 1268 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6544
timestamp 1712256841
transform 1 0 1236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6545
timestamp 1712256841
transform 1 0 1220 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1712256841
transform 1 0 1628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6547
timestamp 1712256841
transform 1 0 1508 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6548
timestamp 1712256841
transform 1 0 1476 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1712256841
transform 1 0 1460 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_6550
timestamp 1712256841
transform 1 0 1452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6551
timestamp 1712256841
transform 1 0 1436 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1712256841
transform 1 0 1732 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6553
timestamp 1712256841
transform 1 0 1708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6554
timestamp 1712256841
transform 1 0 1676 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1712256841
transform 1 0 1644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6556
timestamp 1712256841
transform 1 0 1812 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6557
timestamp 1712256841
transform 1 0 1812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6558
timestamp 1712256841
transform 1 0 1804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6559
timestamp 1712256841
transform 1 0 1796 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6560
timestamp 1712256841
transform 1 0 1788 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1712256841
transform 1 0 1900 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1712256841
transform 1 0 1900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6563
timestamp 1712256841
transform 1 0 1876 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1712256841
transform 1 0 1852 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6565
timestamp 1712256841
transform 1 0 1844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6566
timestamp 1712256841
transform 1 0 2188 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6567
timestamp 1712256841
transform 1 0 2124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6568
timestamp 1712256841
transform 1 0 2108 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6569
timestamp 1712256841
transform 1 0 2108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6570
timestamp 1712256841
transform 1 0 2068 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6571
timestamp 1712256841
transform 1 0 2004 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6572
timestamp 1712256841
transform 1 0 2004 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1712256841
transform 1 0 2004 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6574
timestamp 1712256841
transform 1 0 2292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6575
timestamp 1712256841
transform 1 0 2260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6576
timestamp 1712256841
transform 1 0 2252 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6577
timestamp 1712256841
transform 1 0 2244 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6578
timestamp 1712256841
transform 1 0 2236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1712256841
transform 1 0 2220 0 1 1655
box -2 -2 2 2
use M2_M1  M2_M1_6580
timestamp 1712256841
transform 1 0 2212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1712256841
transform 1 0 2172 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1712256841
transform 1 0 2812 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6583
timestamp 1712256841
transform 1 0 2756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1712256841
transform 1 0 2708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1712256841
transform 1 0 2708 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6586
timestamp 1712256841
transform 1 0 2532 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1712256841
transform 1 0 2436 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6588
timestamp 1712256841
transform 1 0 2428 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1712256841
transform 1 0 3268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6590
timestamp 1712256841
transform 1 0 3140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6591
timestamp 1712256841
transform 1 0 3140 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6592
timestamp 1712256841
transform 1 0 3100 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_6593
timestamp 1712256841
transform 1 0 3060 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6594
timestamp 1712256841
transform 1 0 2428 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6595
timestamp 1712256841
transform 1 0 2332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6596
timestamp 1712256841
transform 1 0 2460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6597
timestamp 1712256841
transform 1 0 2460 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6598
timestamp 1712256841
transform 1 0 2308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6599
timestamp 1712256841
transform 1 0 2812 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6600
timestamp 1712256841
transform 1 0 2772 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6601
timestamp 1712256841
transform 1 0 2500 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6602
timestamp 1712256841
transform 1 0 2388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6603
timestamp 1712256841
transform 1 0 2252 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6604
timestamp 1712256841
transform 1 0 2444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1712256841
transform 1 0 2380 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6606
timestamp 1712256841
transform 1 0 2156 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6607
timestamp 1712256841
transform 1 0 2572 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6608
timestamp 1712256841
transform 1 0 2460 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6609
timestamp 1712256841
transform 1 0 2412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1712256841
transform 1 0 2532 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6611
timestamp 1712256841
transform 1 0 2380 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6612
timestamp 1712256841
transform 1 0 2372 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6613
timestamp 1712256841
transform 1 0 2628 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6614
timestamp 1712256841
transform 1 0 2420 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6615
timestamp 1712256841
transform 1 0 2412 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6616
timestamp 1712256841
transform 1 0 2284 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6617
timestamp 1712256841
transform 1 0 2212 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6618
timestamp 1712256841
transform 1 0 2428 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6619
timestamp 1712256841
transform 1 0 2204 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6620
timestamp 1712256841
transform 1 0 2204 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6621
timestamp 1712256841
transform 1 0 2036 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6622
timestamp 1712256841
transform 1 0 2004 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6623
timestamp 1712256841
transform 1 0 1972 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6624
timestamp 1712256841
transform 1 0 1948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6625
timestamp 1712256841
transform 1 0 1828 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6626
timestamp 1712256841
transform 1 0 1628 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6627
timestamp 1712256841
transform 1 0 2340 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6628
timestamp 1712256841
transform 1 0 2316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6629
timestamp 1712256841
transform 1 0 1940 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6630
timestamp 1712256841
transform 1 0 1932 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6631
timestamp 1712256841
transform 1 0 1588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6632
timestamp 1712256841
transform 1 0 2276 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6633
timestamp 1712256841
transform 1 0 2236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6634
timestamp 1712256841
transform 1 0 1724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6635
timestamp 1712256841
transform 1 0 1596 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6636
timestamp 1712256841
transform 1 0 2100 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1712256841
transform 1 0 2100 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6638
timestamp 1712256841
transform 1 0 2068 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6639
timestamp 1712256841
transform 1 0 1724 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6640
timestamp 1712256841
transform 1 0 1524 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6641
timestamp 1712256841
transform 1 0 1820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6642
timestamp 1712256841
transform 1 0 1788 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6643
timestamp 1712256841
transform 1 0 1660 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6644
timestamp 1712256841
transform 1 0 1468 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6645
timestamp 1712256841
transform 1 0 1204 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6646
timestamp 1712256841
transform 1 0 1916 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6647
timestamp 1712256841
transform 1 0 1900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6648
timestamp 1712256841
transform 1 0 1876 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6649
timestamp 1712256841
transform 1 0 1764 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6650
timestamp 1712256841
transform 1 0 1620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6651
timestamp 1712256841
transform 1 0 1500 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6652
timestamp 1712256841
transform 1 0 1100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6653
timestamp 1712256841
transform 1 0 1740 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6654
timestamp 1712256841
transform 1 0 1684 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6655
timestamp 1712256841
transform 1 0 1684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6656
timestamp 1712256841
transform 1 0 1628 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6657
timestamp 1712256841
transform 1 0 1492 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6658
timestamp 1712256841
transform 1 0 1220 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6659
timestamp 1712256841
transform 1 0 1684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6660
timestamp 1712256841
transform 1 0 1620 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6661
timestamp 1712256841
transform 1 0 1556 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6662
timestamp 1712256841
transform 1 0 1500 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6663
timestamp 1712256841
transform 1 0 1484 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6664
timestamp 1712256841
transform 1 0 1116 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6665
timestamp 1712256841
transform 1 0 1460 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6666
timestamp 1712256841
transform 1 0 1292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1712256841
transform 1 0 772 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6668
timestamp 1712256841
transform 1 0 1356 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6669
timestamp 1712256841
transform 1 0 1268 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1712256841
transform 1 0 684 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6671
timestamp 1712256841
transform 1 0 1332 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6672
timestamp 1712256841
transform 1 0 1300 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6673
timestamp 1712256841
transform 1 0 1236 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6674
timestamp 1712256841
transform 1 0 652 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6675
timestamp 1712256841
transform 1 0 1252 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6676
timestamp 1712256841
transform 1 0 1228 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6677
timestamp 1712256841
transform 1 0 948 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6678
timestamp 1712256841
transform 1 0 716 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6679
timestamp 1712256841
transform 1 0 1252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6680
timestamp 1712256841
transform 1 0 1140 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6681
timestamp 1712256841
transform 1 0 924 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6682
timestamp 1712256841
transform 1 0 820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6683
timestamp 1712256841
transform 1 0 1028 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6684
timestamp 1712256841
transform 1 0 948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6685
timestamp 1712256841
transform 1 0 788 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6686
timestamp 1712256841
transform 1 0 1148 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6687
timestamp 1712256841
transform 1 0 924 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6688
timestamp 1712256841
transform 1 0 812 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6689
timestamp 1712256841
transform 1 0 652 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6690
timestamp 1712256841
transform 1 0 636 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6691
timestamp 1712256841
transform 1 0 1020 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6692
timestamp 1712256841
transform 1 0 900 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6693
timestamp 1712256841
transform 1 0 892 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6694
timestamp 1712256841
transform 1 0 788 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6695
timestamp 1712256841
transform 1 0 764 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6696
timestamp 1712256841
transform 1 0 796 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6697
timestamp 1712256841
transform 1 0 724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6698
timestamp 1712256841
transform 1 0 684 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6699
timestamp 1712256841
transform 1 0 612 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6700
timestamp 1712256841
transform 1 0 612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6701
timestamp 1712256841
transform 1 0 724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6702
timestamp 1712256841
transform 1 0 700 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6703
timestamp 1712256841
transform 1 0 636 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6704
timestamp 1712256841
transform 1 0 540 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6705
timestamp 1712256841
transform 1 0 540 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6706
timestamp 1712256841
transform 1 0 796 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6707
timestamp 1712256841
transform 1 0 716 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6708
timestamp 1712256841
transform 1 0 596 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6709
timestamp 1712256841
transform 1 0 548 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6710
timestamp 1712256841
transform 1 0 540 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6711
timestamp 1712256841
transform 1 0 836 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6712
timestamp 1712256841
transform 1 0 708 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6713
timestamp 1712256841
transform 1 0 708 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6714
timestamp 1712256841
transform 1 0 668 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6715
timestamp 1712256841
transform 1 0 660 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6716
timestamp 1712256841
transform 1 0 612 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6717
timestamp 1712256841
transform 1 0 676 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1712256841
transform 1 0 676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6719
timestamp 1712256841
transform 1 0 948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6720
timestamp 1712256841
transform 1 0 940 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6721
timestamp 1712256841
transform 1 0 1012 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6722
timestamp 1712256841
transform 1 0 996 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6723
timestamp 1712256841
transform 1 0 932 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6724
timestamp 1712256841
transform 1 0 3396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1712256841
transform 1 0 3364 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_6726
timestamp 1712256841
transform 1 0 3292 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6727
timestamp 1712256841
transform 1 0 3268 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_6728
timestamp 1712256841
transform 1 0 2156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6729
timestamp 1712256841
transform 1 0 2156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6730
timestamp 1712256841
transform 1 0 3156 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6731
timestamp 1712256841
transform 1 0 3148 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6732
timestamp 1712256841
transform 1 0 3116 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6733
timestamp 1712256841
transform 1 0 2924 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6734
timestamp 1712256841
transform 1 0 2820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6735
timestamp 1712256841
transform 1 0 2716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6736
timestamp 1712256841
transform 1 0 2596 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6737
timestamp 1712256841
transform 1 0 2588 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1712256841
transform 1 0 3268 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1712256841
transform 1 0 3108 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1712256841
transform 1 0 3148 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1712256841
transform 1 0 2908 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1712256841
transform 1 0 2924 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1712256841
transform 1 0 2844 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1712256841
transform 1 0 3132 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1712256841
transform 1 0 2948 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1712256841
transform 1 0 2868 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1712256841
transform 1 0 3140 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1712256841
transform 1 0 3004 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1712256841
transform 1 0 2916 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1712256841
transform 1 0 2836 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1712256841
transform 1 0 3092 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1712256841
transform 1 0 2988 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1712256841
transform 1 0 2812 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1712256841
transform 1 0 2772 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1712256841
transform 1 0 2716 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1712256841
transform 1 0 2716 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1712256841
transform 1 0 1492 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1712256841
transform 1 0 1492 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1712256841
transform 1 0 1428 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1712256841
transform 1 0 2804 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1712256841
transform 1 0 2732 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1712256841
transform 1 0 2732 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1712256841
transform 1 0 1532 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1712256841
transform 1 0 1444 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1712256841
transform 1 0 1404 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1712256841
transform 1 0 3212 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1712256841
transform 1 0 3076 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1712256841
transform 1 0 3076 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1712256841
transform 1 0 2900 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1712256841
transform 1 0 2892 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1712256841
transform 1 0 2860 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1712256841
transform 1 0 2716 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1712256841
transform 1 0 2572 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1712256841
transform 1 0 2572 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1712256841
transform 1 0 2516 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1712256841
transform 1 0 2508 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1712256841
transform 1 0 2508 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1712256841
transform 1 0 2396 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1712256841
transform 1 0 2396 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1712256841
transform 1 0 2364 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1712256841
transform 1 0 1980 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1712256841
transform 1 0 1652 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1712256841
transform 1 0 1652 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1712256841
transform 1 0 1620 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1712256841
transform 1 0 1620 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1712256841
transform 1 0 1604 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1712256841
transform 1 0 1604 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1712256841
transform 1 0 1436 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1712256841
transform 1 0 1436 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1712256841
transform 1 0 1372 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1712256841
transform 1 0 1364 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1712256841
transform 1 0 1340 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1712256841
transform 1 0 1316 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1712256841
transform 1 0 1316 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1712256841
transform 1 0 1260 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1712256841
transform 1 0 1084 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1712256841
transform 1 0 1012 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1712256841
transform 1 0 748 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1712256841
transform 1 0 724 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1712256841
transform 1 0 692 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1712256841
transform 1 0 692 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1712256841
transform 1 0 676 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1712256841
transform 1 0 676 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1712256841
transform 1 0 668 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1712256841
transform 1 0 668 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1712256841
transform 1 0 636 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1712256841
transform 1 0 636 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1712256841
transform 1 0 620 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1712256841
transform 1 0 620 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1712256841
transform 1 0 596 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1712256841
transform 1 0 3236 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1712256841
transform 1 0 2844 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1712256841
transform 1 0 2732 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1712256841
transform 1 0 2692 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1712256841
transform 1 0 2668 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1712256841
transform 1 0 3308 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1712256841
transform 1 0 3244 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1712256841
transform 1 0 3172 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1712256841
transform 1 0 3100 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1712256841
transform 1 0 2940 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1712256841
transform 1 0 3068 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1712256841
transform 1 0 2988 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1712256841
transform 1 0 2964 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1712256841
transform 1 0 2852 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1712256841
transform 1 0 2940 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1712256841
transform 1 0 2788 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1712256841
transform 1 0 3428 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1712256841
transform 1 0 3308 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1712256841
transform 1 0 3284 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1712256841
transform 1 0 3428 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1712256841
transform 1 0 3308 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1712256841
transform 1 0 3292 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1712256841
transform 1 0 2796 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1712256841
transform 1 0 2692 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1712256841
transform 1 0 3004 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1712256841
transform 1 0 2932 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1712256841
transform 1 0 3228 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1712256841
transform 1 0 3108 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1712256841
transform 1 0 2684 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1712256841
transform 1 0 2548 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1712256841
transform 1 0 2796 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1712256841
transform 1 0 2652 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1712256841
transform 1 0 2556 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1712256841
transform 1 0 2420 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1712256841
transform 1 0 2140 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1712256841
transform 1 0 2020 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1712256841
transform 1 0 2364 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1712256841
transform 1 0 2252 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1712256841
transform 1 0 2196 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1712256841
transform 1 0 2076 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1712256841
transform 1 0 2028 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1712256841
transform 1 0 1980 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1712256841
transform 1 0 1612 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1712256841
transform 1 0 1492 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1712256841
transform 1 0 1372 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1712256841
transform 1 0 1332 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1712256841
transform 1 0 1396 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1712256841
transform 1 0 1260 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1712256841
transform 1 0 1140 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1712256841
transform 1 0 1060 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1712256841
transform 1 0 332 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1712256841
transform 1 0 260 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1712256841
transform 1 0 388 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1712256841
transform 1 0 332 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1712256841
transform 1 0 500 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1712256841
transform 1 0 420 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1712256841
transform 1 0 3420 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1712256841
transform 1 0 3252 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1712256841
transform 1 0 3340 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1712256841
transform 1 0 3284 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1712256841
transform 1 0 3420 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1712256841
transform 1 0 3316 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1712256841
transform 1 0 3380 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1712256841
transform 1 0 3300 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1712256841
transform 1 0 2988 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1712256841
transform 1 0 2796 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1712256841
transform 1 0 3380 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1712256841
transform 1 0 3092 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1712256841
transform 1 0 2980 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1712256841
transform 1 0 2756 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1712256841
transform 1 0 2692 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1712256841
transform 1 0 2948 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1712256841
transform 1 0 2820 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1712256841
transform 1 0 3044 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1712256841
transform 1 0 2860 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1712256841
transform 1 0 2852 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1712256841
transform 1 0 2780 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1712256841
transform 1 0 2660 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1712256841
transform 1 0 2604 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1712256841
transform 1 0 2572 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1712256841
transform 1 0 2492 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1712256841
transform 1 0 2468 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1712256841
transform 1 0 2404 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1712256841
transform 1 0 220 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1712256841
transform 1 0 156 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1712256841
transform 1 0 180 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1712256841
transform 1 0 84 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1712256841
transform 1 0 748 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1712256841
transform 1 0 708 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1712256841
transform 1 0 972 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1712256841
transform 1 0 796 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1712256841
transform 1 0 1284 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1712256841
transform 1 0 1212 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1712256841
transform 1 0 2964 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1712256841
transform 1 0 2876 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1712256841
transform 1 0 2980 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1712256841
transform 1 0 2932 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1712256841
transform 1 0 2732 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1712256841
transform 1 0 2564 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1712256841
transform 1 0 2348 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1712256841
transform 1 0 2268 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1712256841
transform 1 0 2380 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1712256841
transform 1 0 2316 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1712256841
transform 1 0 2308 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1712256841
transform 1 0 2196 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1712256841
transform 1 0 1596 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1712256841
transform 1 0 1532 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1712256841
transform 1 0 3324 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1712256841
transform 1 0 3228 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1712256841
transform 1 0 3204 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1712256841
transform 1 0 3164 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1712256841
transform 1 0 3084 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1712256841
transform 1 0 3268 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1712256841
transform 1 0 3204 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1712256841
transform 1 0 3204 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1712256841
transform 1 0 3188 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1712256841
transform 1 0 3188 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1712256841
transform 1 0 3100 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1712256841
transform 1 0 3100 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1712256841
transform 1 0 3092 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1712256841
transform 1 0 3052 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1712256841
transform 1 0 3020 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1712256841
transform 1 0 2948 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1712256841
transform 1 0 2948 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1712256841
transform 1 0 2908 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1712256841
transform 1 0 2844 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1712256841
transform 1 0 2740 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1712256841
transform 1 0 2892 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1712256841
transform 1 0 2780 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1712256841
transform 1 0 3404 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1712256841
transform 1 0 3364 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1712256841
transform 1 0 3292 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1712256841
transform 1 0 3180 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1712256841
transform 1 0 3276 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1712256841
transform 1 0 3180 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1712256841
transform 1 0 3356 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1712256841
transform 1 0 3284 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1712256841
transform 1 0 3404 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1712256841
transform 1 0 3364 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1712256841
transform 1 0 3316 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1712256841
transform 1 0 3428 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1712256841
transform 1 0 3340 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1712256841
transform 1 0 3428 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1712256841
transform 1 0 3372 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1712256841
transform 1 0 3300 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1712256841
transform 1 0 3292 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1712256841
transform 1 0 3244 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1712256841
transform 1 0 3204 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1712256841
transform 1 0 3164 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1712256841
transform 1 0 3060 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1712256841
transform 1 0 3012 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1712256841
transform 1 0 2932 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1712256841
transform 1 0 2892 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1712256841
transform 1 0 2828 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1712256841
transform 1 0 3348 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1712256841
transform 1 0 3292 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1712256841
transform 1 0 3284 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1712256841
transform 1 0 3276 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1712256841
transform 1 0 3220 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1712256841
transform 1 0 3196 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1712256841
transform 1 0 3060 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1712256841
transform 1 0 3420 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1712256841
transform 1 0 3276 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1712256841
transform 1 0 3268 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1712256841
transform 1 0 3260 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1712256841
transform 1 0 3228 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1712256841
transform 1 0 3228 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1712256841
transform 1 0 3156 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1712256841
transform 1 0 3164 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1712256841
transform 1 0 3068 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1712256841
transform 1 0 2860 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1712256841
transform 1 0 3188 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1712256841
transform 1 0 3116 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1712256841
transform 1 0 3356 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1712256841
transform 1 0 3228 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1712256841
transform 1 0 2708 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1712256841
transform 1 0 2652 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1712256841
transform 1 0 2652 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1712256841
transform 1 0 2612 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1712256841
transform 1 0 2612 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1712256841
transform 1 0 2604 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1712256841
transform 1 0 2604 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1712256841
transform 1 0 2580 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1712256841
transform 1 0 2580 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1712256841
transform 1 0 2356 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1712256841
transform 1 0 1796 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1712256841
transform 1 0 1796 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1712256841
transform 1 0 1700 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1712256841
transform 1 0 1444 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1712256841
transform 1 0 1436 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1712256841
transform 1 0 1236 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1712256841
transform 1 0 3316 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1712256841
transform 1 0 3244 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1712256841
transform 1 0 3236 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1712256841
transform 1 0 3180 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1712256841
transform 1 0 3044 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1712256841
transform 1 0 3044 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1712256841
transform 1 0 2908 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1712256841
transform 1 0 3300 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1712256841
transform 1 0 3204 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1712256841
transform 1 0 3108 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1712256841
transform 1 0 3004 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1712256841
transform 1 0 2972 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1712256841
transform 1 0 2948 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1712256841
transform 1 0 2764 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1712256841
transform 1 0 2668 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1712256841
transform 1 0 2660 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1712256841
transform 1 0 2660 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1712256841
transform 1 0 2628 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1712256841
transform 1 0 2620 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1712256841
transform 1 0 2572 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1712256841
transform 1 0 2540 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1712256841
transform 1 0 2444 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1712256841
transform 1 0 2204 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1712256841
transform 1 0 1956 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1712256841
transform 1 0 1956 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1712256841
transform 1 0 1852 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1712256841
transform 1 0 1788 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1712256841
transform 1 0 1748 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1712256841
transform 1 0 1748 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1712256841
transform 1 0 1748 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1712256841
transform 1 0 1428 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1712256841
transform 1 0 1428 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1712256841
transform 1 0 1428 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1712256841
transform 1 0 1388 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1712256841
transform 1 0 1380 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1712256841
transform 1 0 1060 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1712256841
transform 1 0 1020 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1712256841
transform 1 0 852 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1712256841
transform 1 0 852 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1712256841
transform 1 0 844 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1712256841
transform 1 0 796 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1712256841
transform 1 0 796 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1712256841
transform 1 0 2580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1712256841
transform 1 0 2572 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1712256841
transform 1 0 2524 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1712256841
transform 1 0 2396 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1712256841
transform 1 0 2148 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1712256841
transform 1 0 2148 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1712256841
transform 1 0 1556 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1712256841
transform 1 0 1532 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1712256841
transform 1 0 1492 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1712256841
transform 1 0 1452 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1712256841
transform 1 0 1436 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1712256841
transform 1 0 1428 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1712256841
transform 1 0 1332 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1712256841
transform 1 0 1292 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1712256841
transform 1 0 1052 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1712256841
transform 1 0 980 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1712256841
transform 1 0 948 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1712256841
transform 1 0 1484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1712256841
transform 1 0 1452 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1712256841
transform 1 0 1172 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1712256841
transform 1 0 2876 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1712256841
transform 1 0 2780 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1712256841
transform 1 0 3028 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1712256841
transform 1 0 2916 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1712256841
transform 1 0 3092 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1712256841
transform 1 0 3060 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1712256841
transform 1 0 2972 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1712256841
transform 1 0 2948 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1712256841
transform 1 0 2932 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1712256841
transform 1 0 2836 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1712256841
transform 1 0 2836 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1712256841
transform 1 0 2820 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1712256841
transform 1 0 2812 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1712256841
transform 1 0 2756 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1712256841
transform 1 0 1476 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1712256841
transform 1 0 1452 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1712256841
transform 1 0 2524 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1712256841
transform 1 0 2492 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1712256841
transform 1 0 2492 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1712256841
transform 1 0 2444 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1712256841
transform 1 0 2444 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1712256841
transform 1 0 2340 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1712256841
transform 1 0 2316 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1712256841
transform 1 0 2300 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1712256841
transform 1 0 2260 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1712256841
transform 1 0 2060 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1712256841
transform 1 0 1956 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1712256841
transform 1 0 1924 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1712256841
transform 1 0 1836 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1712256841
transform 1 0 1700 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1712256841
transform 1 0 1700 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1712256841
transform 1 0 1668 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1712256841
transform 1 0 1628 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1712256841
transform 1 0 1612 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1712256841
transform 1 0 2964 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1712256841
transform 1 0 2892 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1712256841
transform 1 0 3012 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1712256841
transform 1 0 2916 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1712256841
transform 1 0 2860 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1712256841
transform 1 0 1012 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1712256841
transform 1 0 908 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1712256841
transform 1 0 1252 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1712256841
transform 1 0 1076 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1712256841
transform 1 0 1028 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1712256841
transform 1 0 916 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1712256841
transform 1 0 2028 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1712256841
transform 1 0 2028 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1712256841
transform 1 0 1972 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1712256841
transform 1 0 1972 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1712256841
transform 1 0 1924 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1712256841
transform 1 0 1740 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1712256841
transform 1 0 1668 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1712256841
transform 1 0 1460 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1712256841
transform 1 0 1428 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1712256841
transform 1 0 820 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1712256841
transform 1 0 692 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1712256841
transform 1 0 644 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1712256841
transform 1 0 1764 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1712256841
transform 1 0 1668 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1712256841
transform 1 0 1620 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1712256841
transform 1 0 3068 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1712256841
transform 1 0 2972 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1712256841
transform 1 0 2788 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1712256841
transform 1 0 2572 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1712256841
transform 1 0 2572 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1712256841
transform 1 0 2412 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1712256841
transform 1 0 2396 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1712256841
transform 1 0 2364 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1712256841
transform 1 0 1700 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1712256841
transform 1 0 1476 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1712256841
transform 1 0 1452 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1712256841
transform 1 0 1940 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1712256841
transform 1 0 1796 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1712256841
transform 1 0 1772 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1712256841
transform 1 0 2652 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1712256841
transform 1 0 2620 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1712256841
transform 1 0 2436 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1712256841
transform 1 0 2412 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1712256841
transform 1 0 2796 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1712256841
transform 1 0 2748 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1712256841
transform 1 0 1292 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1712256841
transform 1 0 1188 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1712256841
transform 1 0 1108 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1712256841
transform 1 0 1108 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1712256841
transform 1 0 1084 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1712256841
transform 1 0 956 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1712256841
transform 1 0 1404 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1712256841
transform 1 0 1092 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1712256841
transform 1 0 2620 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1712256841
transform 1 0 1628 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1712256841
transform 1 0 2908 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1712256841
transform 1 0 2676 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1712256841
transform 1 0 1916 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1712256841
transform 1 0 1476 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1712256841
transform 1 0 1340 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1712256841
transform 1 0 1268 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1712256841
transform 1 0 1260 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1712256841
transform 1 0 1188 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1712256841
transform 1 0 1124 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1712256841
transform 1 0 2940 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1712256841
transform 1 0 2908 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1712256841
transform 1 0 2876 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1712256841
transform 1 0 2756 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1712256841
transform 1 0 756 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1712256841
transform 1 0 732 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1712256841
transform 1 0 1604 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1712256841
transform 1 0 1532 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1712256841
transform 1 0 1500 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1712256841
transform 1 0 2332 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1712256841
transform 1 0 2300 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1712256841
transform 1 0 1564 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1712256841
transform 1 0 1540 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1712256841
transform 1 0 916 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1712256841
transform 1 0 764 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1712256841
transform 1 0 724 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1712256841
transform 1 0 1532 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1712256841
transform 1 0 1492 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1712256841
transform 1 0 1492 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1712256841
transform 1 0 1316 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1712256841
transform 1 0 2772 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1712256841
transform 1 0 2628 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1712256841
transform 1 0 2628 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1712256841
transform 1 0 1684 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1712256841
transform 1 0 3084 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1712256841
transform 1 0 2916 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1712256841
transform 1 0 2292 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1712256841
transform 1 0 2108 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1712256841
transform 1 0 1404 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1712256841
transform 1 0 1332 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1712256841
transform 1 0 1116 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1712256841
transform 1 0 1092 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1712256841
transform 1 0 1068 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1712256841
transform 1 0 1052 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1712256841
transform 1 0 1052 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1712256841
transform 1 0 1004 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1712256841
transform 1 0 1068 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1712256841
transform 1 0 972 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1712256841
transform 1 0 972 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1712256841
transform 1 0 780 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1712256841
transform 1 0 676 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1712256841
transform 1 0 1972 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1712256841
transform 1 0 1852 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1712256841
transform 1 0 1828 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1712256841
transform 1 0 2892 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1712256841
transform 1 0 2828 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1712256841
transform 1 0 2780 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1712256841
transform 1 0 2780 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1712256841
transform 1 0 2652 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1712256841
transform 1 0 2540 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1712256841
transform 1 0 1060 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1712256841
transform 1 0 908 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1712256841
transform 1 0 692 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1712256841
transform 1 0 1884 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1712256841
transform 1 0 1684 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1712256841
transform 1 0 1636 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1712256841
transform 1 0 1420 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1712256841
transform 1 0 2716 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1712256841
transform 1 0 2660 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1712256841
transform 1 0 2692 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1712256841
transform 1 0 2636 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1712256841
transform 1 0 1588 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1712256841
transform 1 0 1556 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1712256841
transform 1 0 3380 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1712256841
transform 1 0 3324 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1712256841
transform 1 0 3252 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1712256841
transform 1 0 3228 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1712256841
transform 1 0 3148 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1712256841
transform 1 0 3076 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1712256841
transform 1 0 2900 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1712256841
transform 1 0 2900 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1712256841
transform 1 0 2748 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1712256841
transform 1 0 2868 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1712256841
transform 1 0 2804 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1712256841
transform 1 0 3020 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1712256841
transform 1 0 2820 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1712256841
transform 1 0 2748 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1712256841
transform 1 0 3084 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1712256841
transform 1 0 2796 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1712256841
transform 1 0 2716 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1712256841
transform 1 0 2716 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1712256841
transform 1 0 2660 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1712256841
transform 1 0 2604 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1712256841
transform 1 0 2572 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1712256841
transform 1 0 2500 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1712256841
transform 1 0 2500 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1712256841
transform 1 0 2468 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1712256841
transform 1 0 2468 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1712256841
transform 1 0 2468 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1712256841
transform 1 0 1260 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1712256841
transform 1 0 1140 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1712256841
transform 1 0 1124 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1712256841
transform 1 0 980 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1712256841
transform 1 0 980 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1712256841
transform 1 0 980 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1712256841
transform 1 0 956 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1712256841
transform 1 0 924 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1712256841
transform 1 0 924 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1712256841
transform 1 0 892 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1712256841
transform 1 0 884 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1712256841
transform 1 0 524 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1712256841
transform 1 0 1340 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1712256841
transform 1 0 812 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1712256841
transform 1 0 580 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1712256841
transform 1 0 444 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1712256841
transform 1 0 428 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1712256841
transform 1 0 356 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1712256841
transform 1 0 356 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1712256841
transform 1 0 316 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1712256841
transform 1 0 308 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1712256841
transform 1 0 300 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1712256841
transform 1 0 292 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1712256841
transform 1 0 292 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1712256841
transform 1 0 292 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1712256841
transform 1 0 292 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1712256841
transform 1 0 260 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1712256841
transform 1 0 260 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1712256841
transform 1 0 148 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1712256841
transform 1 0 92 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1712256841
transform 1 0 1900 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1712256841
transform 1 0 1788 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1712256841
transform 1 0 1636 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1712256841
transform 1 0 1636 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1712256841
transform 1 0 1564 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1712256841
transform 1 0 1564 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1712256841
transform 1 0 1388 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1712256841
transform 1 0 2108 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1712256841
transform 1 0 2052 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1712256841
transform 1 0 2036 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1712256841
transform 1 0 1932 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1712256841
transform 1 0 2556 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1712256841
transform 1 0 2556 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1712256841
transform 1 0 2308 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1712256841
transform 1 0 1044 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1712256841
transform 1 0 1356 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1712256841
transform 1 0 700 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1712256841
transform 1 0 692 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1712256841
transform 1 0 612 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1712256841
transform 1 0 1436 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1712256841
transform 1 0 1372 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1712256841
transform 1 0 1036 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1712256841
transform 1 0 1028 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1712256841
transform 1 0 876 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1712256841
transform 1 0 876 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1712256841
transform 1 0 756 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1712256841
transform 1 0 692 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1712256841
transform 1 0 3116 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1712256841
transform 1 0 3052 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1712256841
transform 1 0 2924 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1712256841
transform 1 0 2756 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1712256841
transform 1 0 2284 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1712256841
transform 1 0 2284 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1712256841
transform 1 0 1996 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1712256841
transform 1 0 1996 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1712256841
transform 1 0 1932 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1712256841
transform 1 0 2628 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1712256841
transform 1 0 2620 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1712256841
transform 1 0 2316 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1712256841
transform 1 0 1324 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1712256841
transform 1 0 1324 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1712256841
transform 1 0 1220 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1712256841
transform 1 0 1196 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1712256841
transform 1 0 1060 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1712256841
transform 1 0 1060 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1712256841
transform 1 0 1028 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1712256841
transform 1 0 964 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1712256841
transform 1 0 940 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1712256841
transform 1 0 924 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1712256841
transform 1 0 916 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1712256841
transform 1 0 860 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1712256841
transform 1 0 604 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1712256841
transform 1 0 492 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1712256841
transform 1 0 3100 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1712256841
transform 1 0 2788 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1712256841
transform 1 0 2412 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1712256841
transform 1 0 2356 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1712256841
transform 1 0 2276 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1712256841
transform 1 0 2244 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1712256841
transform 1 0 2740 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1712256841
transform 1 0 2700 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1712256841
transform 1 0 2676 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1712256841
transform 1 0 2676 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1712256841
transform 1 0 2532 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1712256841
transform 1 0 2524 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1712256841
transform 1 0 1180 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1712256841
transform 1 0 1180 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1712256841
transform 1 0 1148 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1712256841
transform 1 0 1116 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1712256841
transform 1 0 1108 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1712256841
transform 1 0 1260 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1712256841
transform 1 0 1148 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1712256841
transform 1 0 1604 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1712256841
transform 1 0 932 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1712256841
transform 1 0 660 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1712256841
transform 1 0 356 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1712256841
transform 1 0 348 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1712256841
transform 1 0 276 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1712256841
transform 1 0 652 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1712256841
transform 1 0 580 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1712256841
transform 1 0 148 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1712256841
transform 1 0 2612 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1712256841
transform 1 0 2564 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1712256841
transform 1 0 1140 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1712256841
transform 1 0 1140 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1712256841
transform 1 0 1012 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1712256841
transform 1 0 1076 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1712256841
transform 1 0 1028 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1712256841
transform 1 0 972 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1712256841
transform 1 0 916 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1712256841
transform 1 0 1652 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1712256841
transform 1 0 1604 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1712256841
transform 1 0 1236 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1712256841
transform 1 0 1212 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1712256841
transform 1 0 1196 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1712256841
transform 1 0 1196 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1712256841
transform 1 0 1188 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1712256841
transform 1 0 132 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1712256841
transform 1 0 612 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1712256841
transform 1 0 452 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1712256841
transform 1 0 428 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1712256841
transform 1 0 420 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1712256841
transform 1 0 364 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1712256841
transform 1 0 364 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1712256841
transform 1 0 516 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1712256841
transform 1 0 508 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1712256841
transform 1 0 492 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1712256841
transform 1 0 404 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1712256841
transform 1 0 380 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1712256841
transform 1 0 380 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1712256841
transform 1 0 2028 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1712256841
transform 1 0 2028 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1712256841
transform 1 0 1964 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1712256841
transform 1 0 1940 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1712256841
transform 1 0 1812 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1712256841
transform 1 0 1804 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1712256841
transform 1 0 1588 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1712256841
transform 1 0 1548 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1712256841
transform 1 0 1324 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1712256841
transform 1 0 1284 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1712256841
transform 1 0 1252 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1712256841
transform 1 0 3068 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1712256841
transform 1 0 2980 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1712256841
transform 1 0 2404 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1712256841
transform 1 0 2164 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1712256841
transform 1 0 2076 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1712256841
transform 1 0 1996 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1712256841
transform 1 0 2612 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1712256841
transform 1 0 2588 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1712256841
transform 1 0 2588 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1712256841
transform 1 0 2508 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1712256841
transform 1 0 2356 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1712256841
transform 1 0 2356 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1712256841
transform 1 0 1412 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1712256841
transform 1 0 1404 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1712256841
transform 1 0 1244 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1712256841
transform 1 0 1564 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1712256841
transform 1 0 1532 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1712256841
transform 1 0 1172 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1712256841
transform 1 0 1172 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1712256841
transform 1 0 844 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1712256841
transform 1 0 804 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1712256841
transform 1 0 668 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1712256841
transform 1 0 700 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1712256841
transform 1 0 676 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1712256841
transform 1 0 628 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1712256841
transform 1 0 548 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1712256841
transform 1 0 540 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1712256841
transform 1 0 540 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1712256841
transform 1 0 452 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1712256841
transform 1 0 340 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1712256841
transform 1 0 220 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1712256841
transform 1 0 988 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1712256841
transform 1 0 820 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1712256841
transform 1 0 748 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1712256841
transform 1 0 748 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1712256841
transform 1 0 492 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1712256841
transform 1 0 428 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1712256841
transform 1 0 412 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1712256841
transform 1 0 380 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1712256841
transform 1 0 660 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1712256841
transform 1 0 460 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1712256841
transform 1 0 460 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1712256841
transform 1 0 356 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1712256841
transform 1 0 836 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1712256841
transform 1 0 756 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1712256841
transform 1 0 436 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1712256841
transform 1 0 276 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1712256841
transform 1 0 2620 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1712256841
transform 1 0 2596 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1712256841
transform 1 0 2372 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1712256841
transform 1 0 2260 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1712256841
transform 1 0 2956 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1712256841
transform 1 0 2620 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1712256841
transform 1 0 2572 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1712256841
transform 1 0 2572 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1712256841
transform 1 0 2500 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1712256841
transform 1 0 2388 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1712256841
transform 1 0 2556 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1712256841
transform 1 0 2540 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1712256841
transform 1 0 1596 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1712256841
transform 1 0 1572 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1712256841
transform 1 0 1572 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1712256841
transform 1 0 1108 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1712256841
transform 1 0 1100 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1712256841
transform 1 0 1092 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1712256841
transform 1 0 1084 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1712256841
transform 1 0 988 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1712256841
transform 1 0 988 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1712256841
transform 1 0 932 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1712256841
transform 1 0 932 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1712256841
transform 1 0 1364 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1712256841
transform 1 0 1332 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1712256841
transform 1 0 676 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1712256841
transform 1 0 676 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1712256841
transform 1 0 628 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1712256841
transform 1 0 508 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1712256841
transform 1 0 596 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1712256841
transform 1 0 596 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1712256841
transform 1 0 540 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1712256841
transform 1 0 524 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1712256841
transform 1 0 428 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1712256841
transform 1 0 428 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1712256841
transform 1 0 284 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1712256841
transform 1 0 284 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1712256841
transform 1 0 132 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1712256841
transform 1 0 92 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1712256841
transform 1 0 484 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1712256841
transform 1 0 460 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1712256841
transform 1 0 460 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1712256841
transform 1 0 436 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1712256841
transform 1 0 380 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1712256841
transform 1 0 1300 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1712256841
transform 1 0 524 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1712256841
transform 1 0 476 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1712256841
transform 1 0 476 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1712256841
transform 1 0 436 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1712256841
transform 1 0 412 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1712256841
transform 1 0 412 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1712256841
transform 1 0 412 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1712256841
transform 1 0 388 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1712256841
transform 1 0 388 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1712256841
transform 1 0 1244 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1712256841
transform 1 0 988 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1712256841
transform 1 0 1340 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1712256841
transform 1 0 1268 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1712256841
transform 1 0 1268 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1712256841
transform 1 0 1020 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1712256841
transform 1 0 972 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1712256841
transform 1 0 2988 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1712256841
transform 1 0 2772 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1712256841
transform 1 0 2772 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1712256841
transform 1 0 2228 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1712256841
transform 1 0 2212 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1712256841
transform 1 0 2188 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1712256841
transform 1 0 2036 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1712256841
transform 1 0 1996 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1712256841
transform 1 0 1884 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1712256841
transform 1 0 2652 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1712256841
transform 1 0 2580 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1712256841
transform 1 0 2508 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1712256841
transform 1 0 2444 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1712256841
transform 1 0 1852 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1712256841
transform 1 0 1764 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1712256841
transform 1 0 1764 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1712256841
transform 1 0 1764 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1712256841
transform 1 0 1724 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1712256841
transform 1 0 1604 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1712256841
transform 1 0 2636 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1712256841
transform 1 0 2516 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1712256841
transform 1 0 2508 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1712256841
transform 1 0 2484 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1712256841
transform 1 0 1332 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1712256841
transform 1 0 1756 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1712256841
transform 1 0 1556 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1712256841
transform 1 0 1556 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1712256841
transform 1 0 1484 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1712256841
transform 1 0 1308 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1712256841
transform 1 0 1492 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1712256841
transform 1 0 1452 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1712256841
transform 1 0 1044 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1712256841
transform 1 0 1044 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1712256841
transform 1 0 796 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1712256841
transform 1 0 820 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1712256841
transform 1 0 628 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1712256841
transform 1 0 604 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1712256841
transform 1 0 548 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1712256841
transform 1 0 228 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1712256841
transform 1 0 196 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1712256841
transform 1 0 1964 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1712256841
transform 1 0 860 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1712256841
transform 1 0 508 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1712256841
transform 1 0 404 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1712256841
transform 1 0 404 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1712256841
transform 1 0 508 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1712256841
transform 1 0 460 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1712256841
transform 1 0 364 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1712256841
transform 1 0 2796 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1712256841
transform 1 0 2796 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1712256841
transform 1 0 2724 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1712256841
transform 1 0 2724 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1712256841
transform 1 0 2692 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1712256841
transform 1 0 2692 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1712256841
transform 1 0 2660 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1712256841
transform 1 0 2652 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1712256841
transform 1 0 2580 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1712256841
transform 1 0 2572 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1712256841
transform 1 0 2484 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1712256841
transform 1 0 2364 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1712256841
transform 1 0 2300 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1712256841
transform 1 0 2260 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1712256841
transform 1 0 2500 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1712256841
transform 1 0 2420 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1712256841
transform 1 0 1956 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1712256841
transform 1 0 2652 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1712256841
transform 1 0 2652 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1712256841
transform 1 0 2540 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1712256841
transform 1 0 2540 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1712256841
transform 1 0 2492 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1712256841
transform 1 0 2476 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1712256841
transform 1 0 2868 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1712256841
transform 1 0 2188 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1712256841
transform 1 0 1572 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1712256841
transform 1 0 1468 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1712256841
transform 1 0 1084 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1712256841
transform 1 0 1060 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1712256841
transform 1 0 1028 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1712256841
transform 1 0 404 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1712256841
transform 1 0 356 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1712256841
transform 1 0 476 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1712256841
transform 1 0 452 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1712256841
transform 1 0 308 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1712256841
transform 1 0 268 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1712256841
transform 1 0 292 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1712256841
transform 1 0 196 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1712256841
transform 1 0 228 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1712256841
transform 1 0 140 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1712256841
transform 1 0 1148 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1712256841
transform 1 0 1068 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1712256841
transform 1 0 1724 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1712256841
transform 1 0 1644 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1712256841
transform 1 0 2148 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1712256841
transform 1 0 2060 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1712256841
transform 1 0 2036 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1712256841
transform 1 0 1972 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1712256841
transform 1 0 2740 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1712256841
transform 1 0 2660 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1712256841
transform 1 0 2660 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1712256841
transform 1 0 2612 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1712256841
transform 1 0 2876 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1712256841
transform 1 0 2836 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1712256841
transform 1 0 3132 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1712256841
transform 1 0 2980 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1712256841
transform 1 0 2996 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1712256841
transform 1 0 2860 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1712256841
transform 1 0 3404 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1712256841
transform 1 0 3372 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1712256841
transform 1 0 3252 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1712256841
transform 1 0 3196 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1712256841
transform 1 0 3132 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1712256841
transform 1 0 3132 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1712256841
transform 1 0 3084 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1712256841
transform 1 0 3084 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1712256841
transform 1 0 3020 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1712256841
transform 1 0 3260 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1712256841
transform 1 0 3228 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1712256841
transform 1 0 3372 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1712256841
transform 1 0 3292 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1712256841
transform 1 0 3284 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1712256841
transform 1 0 3260 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1712256841
transform 1 0 3284 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1712256841
transform 1 0 3188 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1712256841
transform 1 0 3372 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1712256841
transform 1 0 3300 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1712256841
transform 1 0 3284 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1712256841
transform 1 0 3236 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1712256841
transform 1 0 3372 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1712256841
transform 1 0 3212 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1712256841
transform 1 0 3372 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1712256841
transform 1 0 3332 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1712256841
transform 1 0 3324 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1712256841
transform 1 0 3260 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1712256841
transform 1 0 3260 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1712256841
transform 1 0 3220 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1712256841
transform 1 0 3212 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1712256841
transform 1 0 3204 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1712256841
transform 1 0 3196 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1712256841
transform 1 0 3180 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1712256841
transform 1 0 3140 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1712256841
transform 1 0 3052 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1712256841
transform 1 0 3364 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1712256841
transform 1 0 3324 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1712256841
transform 1 0 3164 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1712256841
transform 1 0 3140 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1712256841
transform 1 0 3140 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1712256841
transform 1 0 3100 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1712256841
transform 1 0 3100 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1712256841
transform 1 0 3076 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1712256841
transform 1 0 2636 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1712256841
transform 1 0 1740 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1712256841
transform 1 0 3364 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1712256841
transform 1 0 3284 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1712256841
transform 1 0 3180 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1712256841
transform 1 0 3148 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1712256841
transform 1 0 3148 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1712256841
transform 1 0 3060 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1712256841
transform 1 0 3028 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1712256841
transform 1 0 2100 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1712256841
transform 1 0 2084 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1712256841
transform 1 0 2020 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1712256841
transform 1 0 2100 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1712256841
transform 1 0 2044 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1712256841
transform 1 0 2044 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1712256841
transform 1 0 1964 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1712256841
transform 1 0 1964 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1712256841
transform 1 0 1940 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1712256841
transform 1 0 1900 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1712256841
transform 1 0 1900 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1712256841
transform 1 0 1852 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1712256841
transform 1 0 2300 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1712256841
transform 1 0 2284 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1712256841
transform 1 0 2308 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1712256841
transform 1 0 2252 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1712256841
transform 1 0 2284 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1712256841
transform 1 0 2260 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1712256841
transform 1 0 2228 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1712256841
transform 1 0 2212 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1712256841
transform 1 0 2172 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1712256841
transform 1 0 2148 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1712256841
transform 1 0 2548 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1712256841
transform 1 0 2436 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1712256841
transform 1 0 2412 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1712256841
transform 1 0 2444 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1712256841
transform 1 0 2444 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1712256841
transform 1 0 2412 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1712256841
transform 1 0 2380 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1712256841
transform 1 0 2284 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1712256841
transform 1 0 2652 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1712256841
transform 1 0 2628 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1712256841
transform 1 0 2124 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1712256841
transform 1 0 1996 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1712256841
transform 1 0 1556 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1712256841
transform 1 0 1532 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1712256841
transform 1 0 1380 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1712256841
transform 1 0 1268 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1712256841
transform 1 0 1268 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1712256841
transform 1 0 1228 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1712256841
transform 1 0 1228 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1712256841
transform 1 0 868 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1712256841
transform 1 0 1636 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1712256841
transform 1 0 1604 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1712256841
transform 1 0 1132 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1712256841
transform 1 0 1020 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1712256841
transform 1 0 940 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1712256841
transform 1 0 1444 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1712256841
transform 1 0 1420 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1712256841
transform 1 0 1156 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1712256841
transform 1 0 1084 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1712256841
transform 1 0 1748 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1712256841
transform 1 0 1716 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1712256841
transform 1 0 1276 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1712256841
transform 1 0 1188 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1712256841
transform 1 0 692 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1712256841
transform 1 0 628 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1712256841
transform 1 0 484 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1712256841
transform 1 0 1172 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1712256841
transform 1 0 1116 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1712256841
transform 1 0 836 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1712256841
transform 1 0 772 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1712256841
transform 1 0 748 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1712256841
transform 1 0 564 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1712256841
transform 1 0 796 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1712256841
transform 1 0 500 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1712256841
transform 1 0 316 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1712256841
transform 1 0 252 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1712256841
transform 1 0 196 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1712256841
transform 1 0 428 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1712256841
transform 1 0 300 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1712256841
transform 1 0 340 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1712256841
transform 1 0 260 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1712256841
transform 1 0 204 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1712256841
transform 1 0 420 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1712256841
transform 1 0 388 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1712256841
transform 1 0 692 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1712256841
transform 1 0 652 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1712256841
transform 1 0 132 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1712256841
transform 1 0 68 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1712256841
transform 1 0 268 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1712256841
transform 1 0 220 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1712256841
transform 1 0 1772 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1712256841
transform 1 0 1684 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1712256841
transform 1 0 748 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1712256841
transform 1 0 676 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1712256841
transform 1 0 724 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1712256841
transform 1 0 692 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1712256841
transform 1 0 868 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1712256841
transform 1 0 788 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1712256841
transform 1 0 740 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1712256841
transform 1 0 1044 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1712256841
transform 1 0 492 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1712256841
transform 1 0 1212 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1712256841
transform 1 0 1164 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1712256841
transform 1 0 1388 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1712256841
transform 1 0 1124 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1712256841
transform 1 0 1124 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1712256841
transform 1 0 1060 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1712256841
transform 1 0 1500 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1712256841
transform 1 0 1420 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1712256841
transform 1 0 1700 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1712256841
transform 1 0 1604 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1712256841
transform 1 0 1580 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1712256841
transform 1 0 1340 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1712256841
transform 1 0 1340 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1712256841
transform 1 0 1124 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1712256841
transform 1 0 1540 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1712256841
transform 1 0 1212 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1712256841
transform 1 0 1148 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1712256841
transform 1 0 1140 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1712256841
transform 1 0 1108 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1712256841
transform 1 0 1084 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1712256841
transform 1 0 988 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1712256841
transform 1 0 1636 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1712256841
transform 1 0 1228 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1712256841
transform 1 0 1540 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1712256841
transform 1 0 1500 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1712256841
transform 1 0 1444 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1712256841
transform 1 0 1404 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1712256841
transform 1 0 1252 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1712256841
transform 1 0 1684 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1712256841
transform 1 0 1604 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1712256841
transform 1 0 1988 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1712256841
transform 1 0 1908 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1712256841
transform 1 0 2164 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1712256841
transform 1 0 1988 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1712256841
transform 1 0 2132 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1712256841
transform 1 0 2084 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1712256841
transform 1 0 1788 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1712256841
transform 1 0 1732 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1712256841
transform 1 0 1676 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1712256841
transform 1 0 2660 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1712256841
transform 1 0 2660 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1712256841
transform 1 0 1924 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1712256841
transform 1 0 1860 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1712256841
transform 1 0 1820 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1712256841
transform 1 0 1716 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1712256841
transform 1 0 2092 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1712256841
transform 1 0 1860 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1712256841
transform 1 0 1860 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1712256841
transform 1 0 1756 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1712256841
transform 1 0 2436 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1712256841
transform 1 0 2372 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1712256841
transform 1 0 2324 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1712256841
transform 1 0 2036 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1712256841
transform 1 0 1972 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1712256841
transform 1 0 2900 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1712256841
transform 1 0 2580 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1712256841
transform 1 0 2580 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1712256841
transform 1 0 2364 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1712256841
transform 1 0 2260 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1712256841
transform 1 0 2188 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1712256841
transform 1 0 2084 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1712256841
transform 1 0 2804 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1712256841
transform 1 0 2716 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1712256841
transform 1 0 2324 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1712256841
transform 1 0 3404 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1712256841
transform 1 0 3348 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1712256841
transform 1 0 3292 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1712256841
transform 1 0 3404 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1712256841
transform 1 0 3364 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1712256841
transform 1 0 3300 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1712256841
transform 1 0 3316 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1712256841
transform 1 0 3276 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1712256841
transform 1 0 3412 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1712256841
transform 1 0 3364 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1712256841
transform 1 0 2892 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1712256841
transform 1 0 2620 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1712256841
transform 1 0 2620 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1712256841
transform 1 0 2572 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1712256841
transform 1 0 3292 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1712256841
transform 1 0 3260 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1712256841
transform 1 0 3220 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1712256841
transform 1 0 3196 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1712256841
transform 1 0 3148 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1712256841
transform 1 0 3036 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1712256841
transform 1 0 2356 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1712256841
transform 1 0 1476 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1712256841
transform 1 0 892 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1712256841
transform 1 0 3340 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1712256841
transform 1 0 3340 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1712256841
transform 1 0 3316 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1712256841
transform 1 0 3316 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1712256841
transform 1 0 2476 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1712256841
transform 1 0 2284 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1712256841
transform 1 0 2116 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1712256841
transform 1 0 2060 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1712256841
transform 1 0 1948 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1712256841
transform 1 0 1948 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1712256841
transform 1 0 1804 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1712256841
transform 1 0 1676 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1712256841
transform 1 0 1588 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1712256841
transform 1 0 1532 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1712256841
transform 1 0 1372 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1712256841
transform 1 0 1292 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1712256841
transform 1 0 1116 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1712256841
transform 1 0 3260 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1712256841
transform 1 0 3236 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1712256841
transform 1 0 3236 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1712256841
transform 1 0 3108 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1712256841
transform 1 0 3108 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1712256841
transform 1 0 3108 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1712256841
transform 1 0 3108 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1712256841
transform 1 0 3076 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1712256841
transform 1 0 3060 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1712256841
transform 1 0 1556 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1712256841
transform 1 0 1556 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1712256841
transform 1 0 1060 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1712256841
transform 1 0 1060 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1712256841
transform 1 0 964 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1712256841
transform 1 0 964 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1712256841
transform 1 0 940 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1712256841
transform 1 0 740 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1712256841
transform 1 0 532 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1712256841
transform 1 0 532 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1712256841
transform 1 0 420 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1712256841
transform 1 0 372 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1712256841
transform 1 0 356 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1712256841
transform 1 0 308 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1712256841
transform 1 0 300 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1712256841
transform 1 0 268 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1712256841
transform 1 0 252 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1712256841
transform 1 0 172 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1712256841
transform 1 0 92 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1712256841
transform 1 0 3348 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1712256841
transform 1 0 3340 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1712256841
transform 1 0 3324 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1712256841
transform 1 0 3268 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1712256841
transform 1 0 3268 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1712256841
transform 1 0 3228 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1712256841
transform 1 0 3132 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1712256841
transform 1 0 3124 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1712256841
transform 1 0 3100 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1712256841
transform 1 0 3060 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1712256841
transform 1 0 3044 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1712256841
transform 1 0 3004 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1712256841
transform 1 0 2988 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1712256841
transform 1 0 2900 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1712256841
transform 1 0 2900 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1712256841
transform 1 0 2860 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1712256841
transform 1 0 2732 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1712256841
transform 1 0 2732 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1712256841
transform 1 0 2716 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1712256841
transform 1 0 2692 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1712256841
transform 1 0 3348 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1712256841
transform 1 0 3340 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1712256841
transform 1 0 3340 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1712256841
transform 1 0 3284 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1712256841
transform 1 0 3268 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1712256841
transform 1 0 3252 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1712256841
transform 1 0 3252 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1712256841
transform 1 0 3156 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1712256841
transform 1 0 2892 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1712256841
transform 1 0 2772 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1712256841
transform 1 0 2692 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1712256841
transform 1 0 2652 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1712256841
transform 1 0 2540 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1712256841
transform 1 0 2420 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1712256841
transform 1 0 2268 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1712256841
transform 1 0 2204 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1712256841
transform 1 0 2116 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1712256841
transform 1 0 2116 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1712256841
transform 1 0 2068 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1712256841
transform 1 0 1964 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1712256841
transform 1 0 1860 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1712256841
transform 1 0 1756 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1712256841
transform 1 0 1660 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1712256841
transform 1 0 1548 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1712256841
transform 1 0 1444 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1712256841
transform 1 0 1332 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1712256841
transform 1 0 1228 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1712256841
transform 1 0 1004 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1712256841
transform 1 0 900 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1712256841
transform 1 0 3052 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1712256841
transform 1 0 2948 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1712256841
transform 1 0 2940 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1712256841
transform 1 0 2372 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1712256841
transform 1 0 2356 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1712256841
transform 1 0 1116 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1712256841
transform 1 0 1100 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1712256841
transform 1 0 788 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1712256841
transform 1 0 676 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1712256841
transform 1 0 572 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1712256841
transform 1 0 436 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1712256841
transform 1 0 420 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1712256841
transform 1 0 300 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1712256841
transform 1 0 196 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1712256841
transform 1 0 140 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1712256841
transform 1 0 2964 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1712256841
transform 1 0 2868 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1712256841
transform 1 0 2772 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1712256841
transform 1 0 2676 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1712256841
transform 1 0 2580 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1712256841
transform 1 0 2484 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1712256841
transform 1 0 2388 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1712256841
transform 1 0 2292 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1712256841
transform 1 0 2196 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1712256841
transform 1 0 2100 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1712256841
transform 1 0 2004 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1712256841
transform 1 0 2004 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1712256841
transform 1 0 1908 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1712256841
transform 1 0 1812 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1712256841
transform 1 0 1876 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1712256841
transform 1 0 1708 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1712256841
transform 1 0 1708 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1712256841
transform 1 0 1596 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1712256841
transform 1 0 1500 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1712256841
transform 1 0 1484 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1712256841
transform 1 0 1468 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1712256841
transform 1 0 1316 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1712256841
transform 1 0 1100 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1712256841
transform 1 0 940 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1712256841
transform 1 0 780 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1712256841
transform 1 0 300 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1712256841
transform 1 0 220 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1712256841
transform 1 0 140 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1712256841
transform 1 0 140 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1712256841
transform 1 0 100 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1712256841
transform 1 0 3348 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1712256841
transform 1 0 3340 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1712256841
transform 1 0 3236 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1712256841
transform 1 0 3228 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1712256841
transform 1 0 3220 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1712256841
transform 1 0 3180 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1712256841
transform 1 0 3180 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1712256841
transform 1 0 3124 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1712256841
transform 1 0 3124 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1712256841
transform 1 0 3124 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1712256841
transform 1 0 3076 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1712256841
transform 1 0 3076 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1712256841
transform 1 0 2932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1712256841
transform 1 0 2812 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1712256841
transform 1 0 1964 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1712256841
transform 1 0 1204 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1712256841
transform 1 0 1204 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1712256841
transform 1 0 892 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1712256841
transform 1 0 668 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1712256841
transform 1 0 556 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1712256841
transform 1 0 444 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1712256841
transform 1 0 332 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1712256841
transform 1 0 2348 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1712256841
transform 1 0 2180 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1712256841
transform 1 0 2172 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1712256841
transform 1 0 1972 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1712256841
transform 1 0 1916 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1712256841
transform 1 0 1868 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1712256841
transform 1 0 2628 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1712256841
transform 1 0 2564 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1712256841
transform 1 0 2644 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1712256841
transform 1 0 2372 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1712256841
transform 1 0 2284 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1712256841
transform 1 0 2444 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1712256841
transform 1 0 2052 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1712256841
transform 1 0 2052 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1712256841
transform 1 0 1892 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1712256841
transform 1 0 1748 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1712256841
transform 1 0 1668 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1712256841
transform 1 0 1612 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1712256841
transform 1 0 1556 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1712256841
transform 1 0 1412 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1712256841
transform 1 0 2780 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1712256841
transform 1 0 2524 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1712256841
transform 1 0 1252 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1712256841
transform 1 0 1252 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1712256841
transform 1 0 1028 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1712256841
transform 1 0 868 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1712256841
transform 1 0 236 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1712256841
transform 1 0 236 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1712256841
transform 1 0 124 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1712256841
transform 1 0 2812 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1712256841
transform 1 0 2620 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1712256841
transform 1 0 2596 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1712256841
transform 1 0 2588 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1712256841
transform 1 0 708 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1712256841
transform 1 0 708 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1712256841
transform 1 0 564 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1712256841
transform 1 0 460 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1712256841
transform 1 0 412 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1712256841
transform 1 0 324 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1712256841
transform 1 0 2732 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1712256841
transform 1 0 2500 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1712256841
transform 1 0 2492 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1712256841
transform 1 0 1212 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1712256841
transform 1 0 1204 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1712256841
transform 1 0 804 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1712256841
transform 1 0 2428 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1712256841
transform 1 0 2324 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1712256841
transform 1 0 2188 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1712256841
transform 1 0 2020 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1712256841
transform 1 0 2884 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1712256841
transform 1 0 2804 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1712256841
transform 1 0 2596 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1712256841
transform 1 0 2596 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1712256841
transform 1 0 2140 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1712256841
transform 1 0 2140 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1712256841
transform 1 0 1228 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1712256841
transform 1 0 820 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1712256841
transform 1 0 732 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1712256841
transform 1 0 636 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1712256841
transform 1 0 572 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1712256841
transform 1 0 452 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1712256841
transform 1 0 388 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1712256841
transform 1 0 388 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1712256841
transform 1 0 316 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1712256841
transform 1 0 252 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1712256841
transform 1 0 180 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1712256841
transform 1 0 140 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1712256841
transform 1 0 3044 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1712256841
transform 1 0 2996 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1712256841
transform 1 0 2940 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1712256841
transform 1 0 3012 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1712256841
transform 1 0 2716 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1712256841
transform 1 0 2628 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1712256841
transform 1 0 2628 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1712256841
transform 1 0 2604 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1712256841
transform 1 0 1972 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1712256841
transform 1 0 1900 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1712256841
transform 1 0 1740 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1712256841
transform 1 0 1540 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1712256841
transform 1 0 1476 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1712256841
transform 1 0 1260 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1712256841
transform 1 0 1244 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1712256841
transform 1 0 1188 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1712256841
transform 1 0 1092 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1712256841
transform 1 0 1092 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1712256841
transform 1 0 324 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1712256841
transform 1 0 324 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1712256841
transform 1 0 212 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1712256841
transform 1 0 3076 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1712256841
transform 1 0 3012 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1712256841
transform 1 0 3012 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1712256841
transform 1 0 2956 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1712256841
transform 1 0 2492 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1712256841
transform 1 0 2636 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1712256841
transform 1 0 2476 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1712256841
transform 1 0 2324 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1712256841
transform 1 0 2324 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1712256841
transform 1 0 2252 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1712256841
transform 1 0 2108 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1712256841
transform 1 0 2108 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1712256841
transform 1 0 2044 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1712256841
transform 1 0 2044 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1712256841
transform 1 0 1932 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1712256841
transform 1 0 1932 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1712256841
transform 1 0 1828 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1712256841
transform 1 0 1676 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1712256841
transform 1 0 1628 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1712256841
transform 1 0 1476 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1712256841
transform 1 0 1364 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1712256841
transform 1 0 1332 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1712256841
transform 1 0 1276 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1712256841
transform 1 0 1236 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1712256841
transform 1 0 1036 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1712256841
transform 1 0 1004 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1712256841
transform 1 0 916 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1712256841
transform 1 0 916 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1712256841
transform 1 0 756 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1712256841
transform 1 0 660 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1712256841
transform 1 0 636 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1712256841
transform 1 0 620 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1712256841
transform 1 0 580 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1712256841
transform 1 0 548 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1712256841
transform 1 0 3060 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1712256841
transform 1 0 2892 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1712256841
transform 1 0 2828 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1712256841
transform 1 0 2724 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1712256841
transform 1 0 2516 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1712256841
transform 1 0 2372 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1712256841
transform 1 0 2212 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1712256841
transform 1 0 2156 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1712256841
transform 1 0 2044 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1712256841
transform 1 0 1980 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1712256841
transform 1 0 1892 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1712256841
transform 1 0 1740 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1712256841
transform 1 0 1620 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1712256841
transform 1 0 1548 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1712256841
transform 1 0 1436 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1712256841
transform 1 0 1436 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1712256841
transform 1 0 1388 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1712256841
transform 1 0 1268 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1712256841
transform 1 0 1212 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1712256841
transform 1 0 2332 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1712256841
transform 1 0 2324 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1712256841
transform 1 0 2300 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1712256841
transform 1 0 2276 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1712256841
transform 1 0 2228 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1712256841
transform 1 0 2228 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1712256841
transform 1 0 2220 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1712256841
transform 1 0 2220 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1712256841
transform 1 0 2172 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1712256841
transform 1 0 2164 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1712256841
transform 1 0 2148 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1712256841
transform 1 0 2148 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1712256841
transform 1 0 2132 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1712256841
transform 1 0 2132 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1712256841
transform 1 0 2132 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1712256841
transform 1 0 2092 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1712256841
transform 1 0 2084 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1712256841
transform 1 0 1780 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1712256841
transform 1 0 1756 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1712256841
transform 1 0 1756 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1712256841
transform 1 0 1692 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1712256841
transform 1 0 1684 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1712256841
transform 1 0 1500 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1712256841
transform 1 0 1492 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1712256841
transform 1 0 1284 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1712256841
transform 1 0 1284 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1712256841
transform 1 0 1100 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1712256841
transform 1 0 772 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1712256841
transform 1 0 764 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1712256841
transform 1 0 612 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1712256841
transform 1 0 500 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1712256841
transform 1 0 500 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1712256841
transform 1 0 212 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1712256841
transform 1 0 212 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1712256841
transform 1 0 140 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1712256841
transform 1 0 140 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1712256841
transform 1 0 132 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1712256841
transform 1 0 132 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1712256841
transform 1 0 108 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1712256841
transform 1 0 100 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1712256841
transform 1 0 92 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1712256841
transform 1 0 92 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1712256841
transform 1 0 92 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1712256841
transform 1 0 84 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1712256841
transform 1 0 2196 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1712256841
transform 1 0 1716 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1712256841
transform 1 0 1652 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1712256841
transform 1 0 1380 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1712256841
transform 1 0 548 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1712256841
transform 1 0 380 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1712256841
transform 1 0 380 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1712256841
transform 1 0 356 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1712256841
transform 1 0 340 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1712256841
transform 1 0 340 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1712256841
transform 1 0 308 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1712256841
transform 1 0 284 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1712256841
transform 1 0 276 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1712256841
transform 1 0 268 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1712256841
transform 1 0 252 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1712256841
transform 1 0 244 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1712256841
transform 1 0 236 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1712256841
transform 1 0 236 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1712256841
transform 1 0 228 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1712256841
transform 1 0 204 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1712256841
transform 1 0 180 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1712256841
transform 1 0 2428 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1712256841
transform 1 0 2420 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1712256841
transform 1 0 2356 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1712256841
transform 1 0 2348 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1712256841
transform 1 0 2348 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1712256841
transform 1 0 2340 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1712256841
transform 1 0 2340 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1712256841
transform 1 0 2292 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1712256841
transform 1 0 2284 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1712256841
transform 1 0 2220 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1712256841
transform 1 0 2204 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1712256841
transform 1 0 2204 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1712256841
transform 1 0 1940 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1712256841
transform 1 0 1940 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1712256841
transform 1 0 1924 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1712256841
transform 1 0 1860 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1712256841
transform 1 0 1796 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1712256841
transform 1 0 1748 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1712256841
transform 1 0 1508 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1712256841
transform 1 0 1508 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1712256841
transform 1 0 1204 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1712256841
transform 1 0 1204 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1712256841
transform 1 0 956 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1712256841
transform 1 0 2148 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1712256841
transform 1 0 2060 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1712256841
transform 1 0 2020 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1712256841
transform 1 0 2020 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1712256841
transform 1 0 2020 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1712256841
transform 1 0 2012 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1712256841
transform 1 0 1916 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1712256841
transform 1 0 1916 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1712256841
transform 1 0 1908 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1712256841
transform 1 0 1732 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1712256841
transform 1 0 1732 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1712256841
transform 1 0 1308 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1712256841
transform 1 0 1308 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1712256841
transform 1 0 612 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1712256841
transform 1 0 524 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1712256841
transform 1 0 276 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1712256841
transform 1 0 268 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1712256841
transform 1 0 244 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1712256841
transform 1 0 244 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1712256841
transform 1 0 196 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1712256841
transform 1 0 196 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1712256841
transform 1 0 196 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1712256841
transform 1 0 172 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1712256841
transform 1 0 140 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1712256841
transform 1 0 140 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1712256841
transform 1 0 124 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1712256841
transform 1 0 116 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1712256841
transform 1 0 2324 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1712256841
transform 1 0 2236 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1712256841
transform 1 0 2236 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1712256841
transform 1 0 2188 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1712256841
transform 1 0 2180 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1712256841
transform 1 0 2180 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1712256841
transform 1 0 2180 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1712256841
transform 1 0 2108 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1712256841
transform 1 0 2068 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1712256841
transform 1 0 1916 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1712256841
transform 1 0 1916 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1712256841
transform 1 0 1844 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1712256841
transform 1 0 1844 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1712256841
transform 1 0 1828 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1712256841
transform 1 0 1756 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1712256841
transform 1 0 1652 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1712256841
transform 1 0 1524 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1712256841
transform 1 0 1164 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1712256841
transform 1 0 1164 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1712256841
transform 1 0 860 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1712256841
transform 1 0 2684 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1712256841
transform 1 0 2660 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1712256841
transform 1 0 3068 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1712256841
transform 1 0 3012 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1712256841
transform 1 0 2972 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1712256841
transform 1 0 2884 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1712256841
transform 1 0 2884 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1712256841
transform 1 0 2836 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1712256841
transform 1 0 2812 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1712256841
transform 1 0 2588 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1712256841
transform 1 0 2468 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1712256841
transform 1 0 1780 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1712256841
transform 1 0 1364 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1712256841
transform 1 0 1148 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1712256841
transform 1 0 2460 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1712256841
transform 1 0 2436 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1712256841
transform 1 0 2388 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1712256841
transform 1 0 2380 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1712256841
transform 1 0 2380 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1712256841
transform 1 0 2300 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1712256841
transform 1 0 2276 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1712256841
transform 1 0 2084 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1712256841
transform 1 0 2076 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1712256841
transform 1 0 2020 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1712256841
transform 1 0 1844 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1712256841
transform 1 0 1700 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1712256841
transform 1 0 1676 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1712256841
transform 1 0 1676 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1712256841
transform 1 0 1636 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1712256841
transform 1 0 1636 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1712256841
transform 1 0 1628 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1712256841
transform 1 0 1484 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1712256841
transform 1 0 1468 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1712256841
transform 1 0 1124 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1712256841
transform 1 0 1044 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1712256841
transform 1 0 972 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1712256841
transform 1 0 948 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1712256841
transform 1 0 948 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1712256841
transform 1 0 804 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1712256841
transform 1 0 804 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1712256841
transform 1 0 700 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1712256841
transform 1 0 684 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1712256841
transform 1 0 668 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1712256841
transform 1 0 668 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1712256841
transform 1 0 636 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1712256841
transform 1 0 636 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1712256841
transform 1 0 628 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1712256841
transform 1 0 628 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1712256841
transform 1 0 612 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1712256841
transform 1 0 596 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1712256841
transform 1 0 596 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1712256841
transform 1 0 588 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1712256841
transform 1 0 580 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1712256841
transform 1 0 580 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1712256841
transform 1 0 548 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1712256841
transform 1 0 548 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1712256841
transform 1 0 532 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1712256841
transform 1 0 532 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1712256841
transform 1 0 516 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1712256841
transform 1 0 508 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1712256841
transform 1 0 3140 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1712256841
transform 1 0 2796 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1712256841
transform 1 0 3148 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1712256841
transform 1 0 3108 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1712256841
transform 1 0 3012 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1712256841
transform 1 0 3012 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1712256841
transform 1 0 2876 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1712256841
transform 1 0 2588 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1712256841
transform 1 0 3188 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1712256841
transform 1 0 3116 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1712256841
transform 1 0 2876 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1712256841
transform 1 0 2844 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1712256841
transform 1 0 2596 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1712256841
transform 1 0 2364 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1712256841
transform 1 0 2364 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1712256841
transform 1 0 2348 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1712256841
transform 1 0 2340 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1712256841
transform 1 0 2316 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1712256841
transform 1 0 2316 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1712256841
transform 1 0 2276 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1712256841
transform 1 0 2252 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1712256841
transform 1 0 2252 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1712256841
transform 1 0 2036 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1712256841
transform 1 0 2036 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1712256841
transform 1 0 1812 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1712256841
transform 1 0 1812 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1712256841
transform 1 0 1668 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1712256841
transform 1 0 1620 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1712256841
transform 1 0 1620 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1712256841
transform 1 0 1500 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1712256841
transform 1 0 1500 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1712256841
transform 1 0 1500 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1712256841
transform 1 0 1452 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1712256841
transform 1 0 1172 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1712256841
transform 1 0 1172 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1712256841
transform 1 0 1100 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1712256841
transform 1 0 924 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1712256841
transform 1 0 772 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1712256841
transform 1 0 700 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1712256841
transform 1 0 700 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1712256841
transform 1 0 628 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1712256841
transform 1 0 556 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1712256841
transform 1 0 2780 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1712256841
transform 1 0 2708 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1712256841
transform 1 0 2708 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1712256841
transform 1 0 2508 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1712256841
transform 1 0 1964 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1712256841
transform 1 0 1532 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1712256841
transform 1 0 1244 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1712256841
transform 1 0 1164 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1712256841
transform 1 0 1164 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1712256841
transform 1 0 988 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1712256841
transform 1 0 980 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1712256841
transform 1 0 916 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1712256841
transform 1 0 916 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1712256841
transform 1 0 852 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1712256841
transform 1 0 852 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1712256841
transform 1 0 580 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1712256841
transform 1 0 580 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1712256841
transform 1 0 572 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1712256841
transform 1 0 548 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1712256841
transform 1 0 548 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1712256841
transform 1 0 492 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1712256841
transform 1 0 2684 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1712256841
transform 1 0 2612 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1712256841
transform 1 0 2444 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1712256841
transform 1 0 3132 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1712256841
transform 1 0 3036 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1712256841
transform 1 0 2996 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1712256841
transform 1 0 2444 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1712256841
transform 1 0 2404 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1712256841
transform 1 0 2396 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1712256841
transform 1 0 2396 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1712256841
transform 1 0 2372 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1712256841
transform 1 0 2308 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1712256841
transform 1 0 2308 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1712256841
transform 1 0 2268 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1712256841
transform 1 0 2268 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1712256841
transform 1 0 2228 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1712256841
transform 1 0 2212 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1712256841
transform 1 0 2212 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1712256841
transform 1 0 2172 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1712256841
transform 1 0 2156 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1712256841
transform 1 0 2156 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1712256841
transform 1 0 2156 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1712256841
transform 1 0 1868 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1712256841
transform 1 0 1852 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1712256841
transform 1 0 1812 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1712256841
transform 1 0 1740 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1712256841
transform 1 0 1444 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1712256841
transform 1 0 1172 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1712256841
transform 1 0 900 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1712256841
transform 1 0 900 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1712256841
transform 1 0 356 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1712256841
transform 1 0 276 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1712256841
transform 1 0 228 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1712256841
transform 1 0 2492 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1712256841
transform 1 0 2492 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1712256841
transform 1 0 2468 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1712256841
transform 1 0 2172 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1712256841
transform 1 0 2140 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1712256841
transform 1 0 2140 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1712256841
transform 1 0 2076 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1712256841
transform 1 0 2076 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1712256841
transform 1 0 1492 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1712256841
transform 1 0 1492 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1712256841
transform 1 0 1212 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1712256841
transform 1 0 1140 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1712256841
transform 1 0 1132 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1712256841
transform 1 0 956 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1712256841
transform 1 0 956 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1712256841
transform 1 0 540 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1712256841
transform 1 0 540 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1712256841
transform 1 0 236 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1712256841
transform 1 0 212 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1712256841
transform 1 0 204 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1712256841
transform 1 0 196 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1712256841
transform 1 0 148 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1712256841
transform 1 0 140 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1712256841
transform 1 0 140 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1712256841
transform 1 0 2844 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1712256841
transform 1 0 2820 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1712256841
transform 1 0 2620 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1712256841
transform 1 0 1660 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1712256841
transform 1 0 1580 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1712256841
transform 1 0 1332 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1712256841
transform 1 0 2628 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1712256841
transform 1 0 2628 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1712256841
transform 1 0 2548 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1712256841
transform 1 0 2516 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1712256841
transform 1 0 2500 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1712256841
transform 1 0 2492 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1712256841
transform 1 0 2348 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1712256841
transform 1 0 2236 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1712256841
transform 1 0 2156 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1712256841
transform 1 0 1972 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1712256841
transform 1 0 1932 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1712256841
transform 1 0 1884 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1712256841
transform 1 0 1772 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1712256841
transform 1 0 1772 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1712256841
transform 1 0 1476 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1712256841
transform 1 0 1332 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1712256841
transform 1 0 1332 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1712256841
transform 1 0 1316 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1712256841
transform 1 0 1316 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1712256841
transform 1 0 1284 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1712256841
transform 1 0 1276 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1712256841
transform 1 0 1276 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1712256841
transform 1 0 1132 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1712256841
transform 1 0 996 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1712256841
transform 1 0 932 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1712256841
transform 1 0 924 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1712256841
transform 1 0 756 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1712256841
transform 1 0 748 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1712256841
transform 1 0 684 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1712256841
transform 1 0 684 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1712256841
transform 1 0 660 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1712256841
transform 1 0 644 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1712256841
transform 1 0 580 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1712256841
transform 1 0 580 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1712256841
transform 1 0 524 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1712256841
transform 1 0 508 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1712256841
transform 1 0 500 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1712256841
transform 1 0 492 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1712256841
transform 1 0 484 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1712256841
transform 1 0 484 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1712256841
transform 1 0 476 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1712256841
transform 1 0 468 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1712256841
transform 1 0 468 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1712256841
transform 1 0 460 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1712256841
transform 1 0 452 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1712256841
transform 1 0 444 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1712256841
transform 1 0 428 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1712256841
transform 1 0 420 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1712256841
transform 1 0 380 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1712256841
transform 1 0 3156 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1712256841
transform 1 0 3124 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1712256841
transform 1 0 3124 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1712256841
transform 1 0 3068 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1712256841
transform 1 0 3012 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1712256841
transform 1 0 2988 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1712256841
transform 1 0 3276 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1712256841
transform 1 0 3196 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1712256841
transform 1 0 3196 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1712256841
transform 1 0 3020 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1712256841
transform 1 0 3012 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1712256841
transform 1 0 2868 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1712256841
transform 1 0 3068 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1712256841
transform 1 0 2980 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1712256841
transform 1 0 2908 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1712256841
transform 1 0 2908 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1712256841
transform 1 0 2780 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1712256841
transform 1 0 2564 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1712256841
transform 1 0 2388 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1712256841
transform 1 0 2388 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1712256841
transform 1 0 2356 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1712256841
transform 1 0 2316 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1712256841
transform 1 0 2300 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1712256841
transform 1 0 2300 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1712256841
transform 1 0 2228 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1712256841
transform 1 0 2228 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1712256841
transform 1 0 2076 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1712256841
transform 1 0 1956 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1712256841
transform 1 0 1956 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1712256841
transform 1 0 1852 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1712256841
transform 1 0 1852 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1712256841
transform 1 0 1804 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1712256841
transform 1 0 1788 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1712256841
transform 1 0 1772 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1712256841
transform 1 0 1764 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1712256841
transform 1 0 1732 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1712256841
transform 1 0 1724 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1712256841
transform 1 0 1612 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1712256841
transform 1 0 1564 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1712256841
transform 1 0 1564 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1712256841
transform 1 0 1516 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1712256841
transform 1 0 1268 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1712256841
transform 1 0 1188 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1712256841
transform 1 0 1108 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1712256841
transform 1 0 1020 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1712256841
transform 1 0 884 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1712256841
transform 1 0 884 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1712256841
transform 1 0 644 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1712256841
transform 1 0 556 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1712256841
transform 1 0 556 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1712256841
transform 1 0 388 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1712256841
transform 1 0 388 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1712256841
transform 1 0 300 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1712256841
transform 1 0 260 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1712256841
transform 1 0 252 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1712256841
transform 1 0 252 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1712256841
transform 1 0 252 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1712256841
transform 1 0 252 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1712256841
transform 1 0 244 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1712256841
transform 1 0 236 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1712256841
transform 1 0 228 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1712256841
transform 1 0 156 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1712256841
transform 1 0 116 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1712256841
transform 1 0 100 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1712256841
transform 1 0 100 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1712256841
transform 1 0 84 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1712256841
transform 1 0 84 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1712256841
transform 1 0 68 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1712256841
transform 1 0 68 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1712256841
transform 1 0 2852 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1712256841
transform 1 0 2828 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1712256841
transform 1 0 2700 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1712256841
transform 1 0 2676 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1712256841
transform 1 0 2660 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1712256841
transform 1 0 2628 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1712256841
transform 1 0 2620 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1712256841
transform 1 0 2476 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1712256841
transform 1 0 2476 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1712256841
transform 1 0 2460 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1712256841
transform 1 0 2044 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1712256841
transform 1 0 1868 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1712256841
transform 1 0 1580 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1712256841
transform 1 0 1284 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1712256841
transform 1 0 1284 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1712256841
transform 1 0 1188 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1712256841
transform 1 0 1164 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1712256841
transform 1 0 1164 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1712256841
transform 1 0 1132 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1712256841
transform 1 0 1132 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1712256841
transform 1 0 2564 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1712256841
transform 1 0 2460 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1712256841
transform 1 0 2284 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1712256841
transform 1 0 2276 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1712256841
transform 1 0 2164 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1712256841
transform 1 0 2164 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1712256841
transform 1 0 2116 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1712256841
transform 1 0 2044 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1712256841
transform 1 0 2044 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1712256841
transform 1 0 2036 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1712256841
transform 1 0 2004 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1712256841
transform 1 0 1804 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1712256841
transform 1 0 1804 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1712256841
transform 1 0 1636 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1712256841
transform 1 0 1604 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1712256841
transform 1 0 1580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1712256841
transform 1 0 1572 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1712256841
transform 1 0 1516 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1712256841
transform 1 0 1268 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1712256841
transform 1 0 1260 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1712256841
transform 1 0 1148 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1712256841
transform 1 0 1124 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1712256841
transform 1 0 1068 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1712256841
transform 1 0 1068 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1712256841
transform 1 0 996 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1712256841
transform 1 0 988 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1712256841
transform 1 0 3308 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1712256841
transform 1 0 3252 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1712256841
transform 1 0 3252 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1712256841
transform 1 0 3172 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1712256841
transform 1 0 1748 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1712256841
transform 1 0 1100 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1712256841
transform 1 0 1100 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1712256841
transform 1 0 1044 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1712256841
transform 1 0 980 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1712256841
transform 1 0 740 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1712256841
transform 1 0 676 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1712256841
transform 1 0 572 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1712256841
transform 1 0 428 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1712256841
transform 1 0 380 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1712256841
transform 1 0 300 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1712256841
transform 1 0 260 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1712256841
transform 1 0 204 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1712256841
transform 1 0 196 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1712256841
transform 1 0 132 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1712256841
transform 1 0 92 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1712256841
transform 1 0 2852 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1712256841
transform 1 0 2652 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1712256841
transform 1 0 2652 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1712256841
transform 1 0 2420 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1712256841
transform 1 0 2300 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1712256841
transform 1 0 2244 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1712256841
transform 1 0 2084 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1712256841
transform 1 0 2020 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1712256841
transform 1 0 1988 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1712256841
transform 1 0 1844 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1712256841
transform 1 0 1788 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1712256841
transform 1 0 1676 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1712256841
transform 1 0 1468 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1712256841
transform 1 0 1468 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1712256841
transform 1 0 1396 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1712256841
transform 1 0 1364 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1712256841
transform 1 0 3380 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1712256841
transform 1 0 3380 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1712256841
transform 1 0 3324 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1712256841
transform 1 0 3276 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1712256841
transform 1 0 3276 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1712256841
transform 1 0 3156 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1712256841
transform 1 0 3092 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1712256841
transform 1 0 3028 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1712256841
transform 1 0 3028 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1712256841
transform 1 0 2988 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1712256841
transform 1 0 2964 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1712256841
transform 1 0 2836 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1712256841
transform 1 0 2804 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1712256841
transform 1 0 2804 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1712256841
transform 1 0 2700 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1712256841
transform 1 0 2604 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1712256841
transform 1 0 2460 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1712256841
transform 1 0 1316 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1712256841
transform 1 0 1780 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1712256841
transform 1 0 1540 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1712256841
transform 1 0 1532 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1712256841
transform 1 0 1308 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1712256841
transform 1 0 1228 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1712256841
transform 1 0 1164 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1712256841
transform 1 0 1004 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1712256841
transform 1 0 740 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1712256841
transform 1 0 700 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1712256841
transform 1 0 628 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1712256841
transform 1 0 588 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1712256841
transform 1 0 588 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1712256841
transform 1 0 548 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1712256841
transform 1 0 508 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1712256841
transform 1 0 508 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1712256841
transform 1 0 2580 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1712256841
transform 1 0 2548 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1712256841
transform 1 0 2404 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1712256841
transform 1 0 2292 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1712256841
transform 1 0 2292 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1712256841
transform 1 0 2212 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1712256841
transform 1 0 2068 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1712256841
transform 1 0 2012 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1712256841
transform 1 0 2012 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1712256841
transform 1 0 1868 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1712256841
transform 1 0 1868 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1712256841
transform 1 0 1636 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1712256841
transform 1 0 1572 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1712256841
transform 1 0 1572 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1712256841
transform 1 0 1492 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1712256841
transform 1 0 1420 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1712256841
transform 1 0 1332 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1712256841
transform 1 0 1332 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1712256841
transform 1 0 972 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1712256841
transform 1 0 3348 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1712256841
transform 1 0 3292 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1712256841
transform 1 0 3284 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1712256841
transform 1 0 3268 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1712256841
transform 1 0 3244 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1712256841
transform 1 0 3228 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1712256841
transform 1 0 3228 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1712256841
transform 1 0 3188 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1712256841
transform 1 0 3188 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1712256841
transform 1 0 3180 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1712256841
transform 1 0 3140 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1712256841
transform 1 0 3036 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1712256841
transform 1 0 3036 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1712256841
transform 1 0 2884 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1712256841
transform 1 0 2700 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1712256841
transform 1 0 2700 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1712256841
transform 1 0 1628 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1712256841
transform 1 0 1436 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1712256841
transform 1 0 1404 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1712256841
transform 1 0 1404 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1712256841
transform 1 0 1364 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1712256841
transform 1 0 2876 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1712256841
transform 1 0 2804 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1712256841
transform 1 0 2620 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1712256841
transform 1 0 2532 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1712256841
transform 1 0 2412 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1712256841
transform 1 0 2148 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1712256841
transform 1 0 2076 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1712256841
transform 1 0 2076 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1712256841
transform 1 0 1612 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1712256841
transform 1 0 1572 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1712256841
transform 1 0 1572 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1712256841
transform 1 0 1492 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1712256841
transform 1 0 1476 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1712256841
transform 1 0 1460 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1712256841
transform 1 0 1380 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1712256841
transform 1 0 1300 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1712256841
transform 1 0 1252 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1712256841
transform 1 0 1252 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1712256841
transform 1 0 1204 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1712256841
transform 1 0 1204 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1712256841
transform 1 0 1084 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1712256841
transform 1 0 996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1712256841
transform 1 0 996 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1712256841
transform 1 0 2620 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1712256841
transform 1 0 2580 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1712256841
transform 1 0 2540 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1712256841
transform 1 0 2380 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1712256841
transform 1 0 2380 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1712256841
transform 1 0 2164 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1712256841
transform 1 0 2164 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1712256841
transform 1 0 1804 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1712256841
transform 1 0 1804 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1712256841
transform 1 0 1796 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1712256841
transform 1 0 1772 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1712256841
transform 1 0 1660 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1712256841
transform 1 0 1660 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1712256841
transform 1 0 1652 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1712256841
transform 1 0 1364 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1712256841
transform 1 0 1276 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1712256841
transform 1 0 1212 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1712256841
transform 1 0 1212 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1712256841
transform 1 0 1204 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1712256841
transform 1 0 1204 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1712256841
transform 1 0 1108 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1712256841
transform 1 0 1092 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1712256841
transform 1 0 1076 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1712256841
transform 1 0 1012 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1712256841
transform 1 0 996 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1712256841
transform 1 0 884 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1712256841
transform 1 0 884 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1712256841
transform 1 0 820 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1712256841
transform 1 0 812 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1712256841
transform 1 0 3100 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1712256841
transform 1 0 3092 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1712256841
transform 1 0 3092 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1712256841
transform 1 0 3060 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1712256841
transform 1 0 3060 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1712256841
transform 1 0 3028 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1712256841
transform 1 0 3020 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1712256841
transform 1 0 2948 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1712256841
transform 1 0 2948 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1712256841
transform 1 0 2484 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1712256841
transform 1 0 2476 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1712256841
transform 1 0 2444 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1712256841
transform 1 0 2188 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1712256841
transform 1 0 2188 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1712256841
transform 1 0 2164 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1712256841
transform 1 0 2052 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1712256841
transform 1 0 1980 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1712256841
transform 1 0 1956 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1712256841
transform 1 0 1924 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1712256841
transform 1 0 3100 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1712256841
transform 1 0 3100 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1712256841
transform 1 0 3060 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1712256841
transform 1 0 3060 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1712256841
transform 1 0 2972 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1712256841
transform 1 0 2972 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1712256841
transform 1 0 2948 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1712256841
transform 1 0 2940 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1712256841
transform 1 0 2708 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1712256841
transform 1 0 2116 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1712256841
transform 1 0 2092 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1712256841
transform 1 0 1980 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1712256841
transform 1 0 1980 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1712256841
transform 1 0 1956 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1712256841
transform 1 0 1956 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1712256841
transform 1 0 1884 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1712256841
transform 1 0 1876 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1712256841
transform 1 0 1764 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1712256841
transform 1 0 1764 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1712256841
transform 1 0 1740 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1712256841
transform 1 0 1716 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1712256841
transform 1 0 2428 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1712256841
transform 1 0 2412 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1712256841
transform 1 0 2388 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1712256841
transform 1 0 2380 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1712256841
transform 1 0 2372 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1712256841
transform 1 0 2308 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1712256841
transform 1 0 2276 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1712256841
transform 1 0 2276 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1712256841
transform 1 0 2212 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1712256841
transform 1 0 2204 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1712256841
transform 1 0 2156 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1712256841
transform 1 0 2084 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1712256841
transform 1 0 2228 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1712256841
transform 1 0 2172 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1712256841
transform 1 0 2132 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1712256841
transform 1 0 2108 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1712256841
transform 1 0 1916 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1712256841
transform 1 0 1916 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1712256841
transform 1 0 1884 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1712256841
transform 1 0 1836 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1712256841
transform 1 0 1828 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1712256841
transform 1 0 1748 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1712256841
transform 1 0 1628 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1712256841
transform 1 0 1628 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1712256841
transform 1 0 2340 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1712256841
transform 1 0 2276 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1712256841
transform 1 0 2276 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1712256841
transform 1 0 2244 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1712256841
transform 1 0 1668 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1712256841
transform 1 0 1628 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1712256841
transform 1 0 1532 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1712256841
transform 1 0 1460 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1712256841
transform 1 0 1452 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1712256841
transform 1 0 1356 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1712256841
transform 1 0 1212 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1712256841
transform 1 0 1060 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1712256841
transform 1 0 772 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1712256841
transform 1 0 764 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1712256841
transform 1 0 764 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1712256841
transform 1 0 764 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1712256841
transform 1 0 740 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1712256841
transform 1 0 740 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1712256841
transform 1 0 668 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1712256841
transform 1 0 1364 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1712256841
transform 1 0 1316 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1712256841
transform 1 0 1236 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1712256841
transform 1 0 980 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1712256841
transform 1 0 948 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1712256841
transform 1 0 940 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1712256841
transform 1 0 916 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1712256841
transform 1 0 884 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1712256841
transform 1 0 860 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1712256841
transform 1 0 788 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1712256841
transform 1 0 780 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1712256841
transform 1 0 764 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1712256841
transform 1 0 636 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1712256841
transform 1 0 580 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1712256841
transform 1 0 396 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1712256841
transform 1 0 396 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1712256841
transform 1 0 236 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1712256841
transform 1 0 196 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1712256841
transform 1 0 1700 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1712256841
transform 1 0 1700 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1712256841
transform 1 0 1668 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1712256841
transform 1 0 1388 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1712256841
transform 1 0 1388 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1712256841
transform 1 0 1204 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1712256841
transform 1 0 1204 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1712256841
transform 1 0 940 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1712256841
transform 1 0 940 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1712256841
transform 1 0 820 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1712256841
transform 1 0 820 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1712256841
transform 1 0 764 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1712256841
transform 1 0 372 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1712256841
transform 1 0 308 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1712256841
transform 1 0 252 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1712256841
transform 1 0 220 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1712256841
transform 1 0 908 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1712256841
transform 1 0 852 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1712256841
transform 1 0 772 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1712256841
transform 1 0 588 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1712256841
transform 1 0 460 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1712256841
transform 1 0 460 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1712256841
transform 1 0 444 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1712256841
transform 1 0 412 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1712256841
transform 1 0 412 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1712256841
transform 1 0 388 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1712256841
transform 1 0 388 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1712256841
transform 1 0 364 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1712256841
transform 1 0 324 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1712256841
transform 1 0 324 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1712256841
transform 1 0 300 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1712256841
transform 1 0 108 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1712256841
transform 1 0 1260 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1712256841
transform 1 0 1252 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1712256841
transform 1 0 1220 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1712256841
transform 1 0 724 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1712256841
transform 1 0 724 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1712256841
transform 1 0 708 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1712256841
transform 1 0 612 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1712256841
transform 1 0 508 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1712256841
transform 1 0 300 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1712256841
transform 1 0 292 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1712256841
transform 1 0 284 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1712256841
transform 1 0 236 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1712256841
transform 1 0 236 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1712256841
transform 1 0 236 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1712256841
transform 1 0 1372 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1712256841
transform 1 0 1332 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1712256841
transform 1 0 1300 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1712256841
transform 1 0 1300 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1712256841
transform 1 0 1284 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1712256841
transform 1 0 1284 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1712256841
transform 1 0 1204 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1712256841
transform 1 0 1140 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1712256841
transform 1 0 1140 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1712256841
transform 1 0 1092 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1712256841
transform 1 0 924 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1712256841
transform 1 0 924 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1712256841
transform 1 0 852 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1712256841
transform 1 0 780 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1712256841
transform 1 0 684 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1712256841
transform 1 0 3436 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1712256841
transform 1 0 3436 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1712256841
transform 1 0 3412 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1712256841
transform 1 0 3412 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1712256841
transform 1 0 3388 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1712256841
transform 1 0 3356 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1712256841
transform 1 0 3348 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1712256841
transform 1 0 3260 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1712256841
transform 1 0 3220 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1712256841
transform 1 0 3212 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1712256841
transform 1 0 3188 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1712256841
transform 1 0 3188 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1712256841
transform 1 0 3092 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1712256841
transform 1 0 3396 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1712256841
transform 1 0 3172 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1712256841
transform 1 0 3148 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1712256841
transform 1 0 3132 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1712256841
transform 1 0 3116 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1712256841
transform 1 0 3308 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1712256841
transform 1 0 2964 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1712256841
transform 1 0 2964 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1712256841
transform 1 0 2948 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1712256841
transform 1 0 2644 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1712256841
transform 1 0 2644 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1712256841
transform 1 0 1772 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1712256841
transform 1 0 3244 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1712256841
transform 1 0 3092 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1712256841
transform 1 0 2564 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1712256841
transform 1 0 2484 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1712256841
transform 1 0 2684 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1712256841
transform 1 0 2652 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1712256841
transform 1 0 2652 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1712256841
transform 1 0 2636 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1712256841
transform 1 0 2588 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1712256841
transform 1 0 1668 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1712256841
transform 1 0 1628 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1712256841
transform 1 0 1412 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1712256841
transform 1 0 1108 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1712256841
transform 1 0 1444 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1712256841
transform 1 0 1412 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1712256841
transform 1 0 1412 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1712256841
transform 1 0 1412 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1712256841
transform 1 0 1316 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1712256841
transform 1 0 1220 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1712256841
transform 1 0 1204 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1712256841
transform 1 0 2948 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1712256841
transform 1 0 2924 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1712256841
transform 1 0 2852 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1712256841
transform 1 0 2732 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1712256841
transform 1 0 2732 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1712256841
transform 1 0 2660 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1712256841
transform 1 0 2388 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1712256841
transform 1 0 1532 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1712256841
transform 1 0 1516 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1712256841
transform 1 0 1484 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1712256841
transform 1 0 1388 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1712256841
transform 1 0 3220 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1712256841
transform 1 0 3172 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1712256841
transform 1 0 3172 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1712256841
transform 1 0 3140 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1712256841
transform 1 0 3108 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1712256841
transform 1 0 3060 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1712256841
transform 1 0 3220 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1712256841
transform 1 0 2796 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1712256841
transform 1 0 1636 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1712256841
transform 1 0 3332 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1712256841
transform 1 0 3252 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1712256841
transform 1 0 3252 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1712256841
transform 1 0 3164 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1712256841
transform 1 0 3148 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1712256841
transform 1 0 3196 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1712256841
transform 1 0 2324 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1712256841
transform 1 0 3388 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1712256841
transform 1 0 3340 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1712256841
transform 1 0 1468 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1712256841
transform 1 0 1292 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1712256841
transform 1 0 1212 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1712256841
transform 1 0 1164 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1712256841
transform 1 0 1436 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1712256841
transform 1 0 1380 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1712256841
transform 1 0 1380 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1712256841
transform 1 0 852 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1712256841
transform 1 0 852 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1712256841
transform 1 0 764 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1712256841
transform 1 0 1348 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1712256841
transform 1 0 1252 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1712256841
transform 1 0 1220 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1712256841
transform 1 0 1036 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1712256841
transform 1 0 964 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1712256841
transform 1 0 868 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1712256841
transform 1 0 2332 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1712256841
transform 1 0 2244 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1712256841
transform 1 0 2244 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1712256841
transform 1 0 2084 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1712256841
transform 1 0 1908 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1712256841
transform 1 0 1604 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1712256841
transform 1 0 1604 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1712256841
transform 1 0 1532 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1712256841
transform 1 0 1452 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1712256841
transform 1 0 1412 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1712256841
transform 1 0 964 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1712256841
transform 1 0 724 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1712256841
transform 1 0 1052 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1712256841
transform 1 0 636 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1712256841
transform 1 0 564 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1712256841
transform 1 0 500 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1712256841
transform 1 0 468 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1712256841
transform 1 0 468 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1712256841
transform 1 0 468 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1712256841
transform 1 0 316 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1712256841
transform 1 0 308 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1712256841
transform 1 0 276 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1712256841
transform 1 0 236 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1712256841
transform 1 0 2996 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1712256841
transform 1 0 2852 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1712256841
transform 1 0 2836 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1712256841
transform 1 0 2684 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1712256841
transform 1 0 2676 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1712256841
transform 1 0 2636 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1712256841
transform 1 0 2116 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1712256841
transform 1 0 2116 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1712256841
transform 1 0 1956 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1712256841
transform 1 0 1028 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1712256841
transform 1 0 828 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1712256841
transform 1 0 828 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1712256841
transform 1 0 628 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1712256841
transform 1 0 628 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1712256841
transform 1 0 596 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1712256841
transform 1 0 564 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1712256841
transform 1 0 356 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1712256841
transform 1 0 316 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1712256841
transform 1 0 260 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1712256841
transform 1 0 212 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1712256841
transform 1 0 212 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1712256841
transform 1 0 2700 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1712256841
transform 1 0 2668 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1712256841
transform 1 0 2668 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1712256841
transform 1 0 2596 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1712256841
transform 1 0 2508 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1712256841
transform 1 0 2500 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1712256841
transform 1 0 2476 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1712256841
transform 1 0 2452 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1712256841
transform 1 0 2444 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1712256841
transform 1 0 2444 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1712256841
transform 1 0 2356 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1712256841
transform 1 0 2332 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1712256841
transform 1 0 2276 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1712256841
transform 1 0 2172 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1712256841
transform 1 0 2092 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1712256841
transform 1 0 2036 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1712256841
transform 1 0 1860 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1712256841
transform 1 0 1860 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1712256841
transform 1 0 1860 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1712256841
transform 1 0 1852 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1712256841
transform 1 0 1788 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1712256841
transform 1 0 1780 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1712256841
transform 1 0 1724 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1712256841
transform 1 0 1628 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1712256841
transform 1 0 1628 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1712256841
transform 1 0 1420 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1712256841
transform 1 0 1420 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1712256841
transform 1 0 1332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1712256841
transform 1 0 1300 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1712256841
transform 1 0 1300 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1712256841
transform 1 0 1100 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1712256841
transform 1 0 964 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1712256841
transform 1 0 716 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1712256841
transform 1 0 716 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1712256841
transform 1 0 460 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1712256841
transform 1 0 452 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1712256841
transform 1 0 452 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1712256841
transform 1 0 452 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1712256841
transform 1 0 444 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1712256841
transform 1 0 444 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1712256841
transform 1 0 436 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1712256841
transform 1 0 436 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1712256841
transform 1 0 420 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1712256841
transform 1 0 420 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1712256841
transform 1 0 420 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1712256841
transform 1 0 420 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1712256841
transform 1 0 420 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1712256841
transform 1 0 404 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1712256841
transform 1 0 396 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1712256841
transform 1 0 396 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1712256841
transform 1 0 396 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1712256841
transform 1 0 364 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1712256841
transform 1 0 364 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1712256841
transform 1 0 356 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1712256841
transform 1 0 348 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1712256841
transform 1 0 348 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1712256841
transform 1 0 332 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1712256841
transform 1 0 332 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1712256841
transform 1 0 324 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1712256841
transform 1 0 244 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1712256841
transform 1 0 244 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1712256841
transform 1 0 2716 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1712256841
transform 1 0 2692 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1712256841
transform 1 0 2668 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1712256841
transform 1 0 2588 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1712256841
transform 1 0 2588 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1712256841
transform 1 0 2188 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1712256841
transform 1 0 3372 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1712256841
transform 1 0 3276 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1712256841
transform 1 0 3052 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1712256841
transform 1 0 2972 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1712256841
transform 1 0 3356 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1712256841
transform 1 0 3316 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1712256841
transform 1 0 2940 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1712256841
transform 1 0 2892 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1712256841
transform 1 0 3436 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1712256841
transform 1 0 3388 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1712256841
transform 1 0 3436 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1712256841
transform 1 0 3436 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1712256841
transform 1 0 3396 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1712256841
transform 1 0 3396 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1712256841
transform 1 0 3412 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1712256841
transform 1 0 3372 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1712256841
transform 1 0 3324 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1712256841
transform 1 0 3324 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1712256841
transform 1 0 2964 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1712256841
transform 1 0 2876 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1712256841
transform 1 0 2780 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1712256841
transform 1 0 2724 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1712256841
transform 1 0 3340 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1712256841
transform 1 0 3276 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1712256841
transform 1 0 2772 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1712256841
transform 1 0 2684 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1712256841
transform 1 0 3188 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1712256841
transform 1 0 2788 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1712256841
transform 1 0 2724 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1712256841
transform 1 0 2724 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1712256841
transform 1 0 2628 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1712256841
transform 1 0 3220 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1712256841
transform 1 0 3108 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1712256841
transform 1 0 2732 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1712256841
transform 1 0 2708 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1712256841
transform 1 0 2692 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1712256841
transform 1 0 2580 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1712256841
transform 1 0 2940 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1712256841
transform 1 0 2836 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1712256841
transform 1 0 2828 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1712256841
transform 1 0 2796 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1712256841
transform 1 0 2700 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1712256841
transform 1 0 3260 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1712256841
transform 1 0 3060 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1712256841
transform 1 0 3372 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1712256841
transform 1 0 3308 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1712256841
transform 1 0 3284 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1712256841
transform 1 0 3228 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1712256841
transform 1 0 2844 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1712256841
transform 1 0 2820 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1712256841
transform 1 0 2140 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1712256841
transform 1 0 2052 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1712256841
transform 1 0 1828 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1712256841
transform 1 0 1756 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1712256841
transform 1 0 1700 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1712256841
transform 1 0 1644 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1712256841
transform 1 0 804 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1712256841
transform 1 0 652 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1712256841
transform 1 0 252 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1712256841
transform 1 0 132 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1712256841
transform 1 0 420 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1712256841
transform 1 0 380 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1712256841
transform 1 0 724 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1712256841
transform 1 0 604 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1712256841
transform 1 0 796 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1712256841
transform 1 0 708 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1712256841
transform 1 0 1092 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1712256841
transform 1 0 940 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1712256841
transform 1 0 1340 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1712256841
transform 1 0 1252 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1712256841
transform 1 0 2092 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1712256841
transform 1 0 1636 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1712256841
transform 1 0 3412 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1712256841
transform 1 0 3364 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1712256841
transform 1 0 3196 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1712256841
transform 1 0 3100 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1712256841
transform 1 0 2956 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1712256841
transform 1 0 3228 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1712256841
transform 1 0 3180 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1712256841
transform 1 0 2756 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1712256841
transform 1 0 2684 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1712256841
transform 1 0 2684 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1712256841
transform 1 0 2572 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1712256841
transform 1 0 3412 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1712256841
transform 1 0 3372 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1712256841
transform 1 0 3308 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1712256841
transform 1 0 3340 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1712256841
transform 1 0 3292 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1712256841
transform 1 0 2900 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1712256841
transform 1 0 1708 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1712256841
transform 1 0 1708 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1712256841
transform 1 0 1612 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1712256841
transform 1 0 1692 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1712256841
transform 1 0 1580 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1712256841
transform 1 0 1572 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1712256841
transform 1 0 1500 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1712256841
transform 1 0 1532 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1712256841
transform 1 0 1444 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1712256841
transform 1 0 1492 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1712256841
transform 1 0 1468 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1712256841
transform 1 0 1572 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1712256841
transform 1 0 1484 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1712256841
transform 1 0 1548 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1712256841
transform 1 0 1492 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1712256841
transform 1 0 2116 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1712256841
transform 1 0 1508 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1712256841
transform 1 0 1492 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1712256841
transform 1 0 860 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1712256841
transform 1 0 836 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1712256841
transform 1 0 268 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1712256841
transform 1 0 868 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1712256841
transform 1 0 844 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1712256841
transform 1 0 1044 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1712256841
transform 1 0 852 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1712256841
transform 1 0 852 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1712256841
transform 1 0 668 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1712256841
transform 1 0 1724 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1712256841
transform 1 0 1428 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1712256841
transform 1 0 1428 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1712256841
transform 1 0 828 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1712256841
transform 1 0 828 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1712256841
transform 1 0 660 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1712256841
transform 1 0 1020 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1712256841
transform 1 0 868 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1712256841
transform 1 0 1540 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1712256841
transform 1 0 1508 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1712256841
transform 1 0 1476 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1712256841
transform 1 0 1300 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1712256841
transform 1 0 1004 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1712256841
transform 1 0 1324 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1712256841
transform 1 0 1196 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1712256841
transform 1 0 1044 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1712256841
transform 1 0 668 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1712256841
transform 1 0 524 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1712256841
transform 1 0 356 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1712256841
transform 1 0 740 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1712256841
transform 1 0 684 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1712256841
transform 1 0 588 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1712256841
transform 1 0 1172 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1712256841
transform 1 0 1012 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1712256841
transform 1 0 972 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1712256841
transform 1 0 900 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1712256841
transform 1 0 1284 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1712256841
transform 1 0 1108 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1712256841
transform 1 0 220 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1712256841
transform 1 0 180 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1712256841
transform 1 0 236 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1712256841
transform 1 0 188 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1712256841
transform 1 0 300 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1712256841
transform 1 0 180 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1712256841
transform 1 0 268 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1712256841
transform 1 0 180 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1712256841
transform 1 0 324 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1712256841
transform 1 0 236 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1712256841
transform 1 0 212 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1712256841
transform 1 0 524 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1712256841
transform 1 0 308 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1712256841
transform 1 0 268 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1712256841
transform 1 0 212 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1712256841
transform 1 0 548 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1712256841
transform 1 0 180 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1712256841
transform 1 0 252 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2584
timestamp 1712256841
transform 1 0 220 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1712256841
transform 1 0 2212 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1712256841
transform 1 0 2180 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1712256841
transform 1 0 2220 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1712256841
transform 1 0 1956 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1712256841
transform 1 0 1956 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1712256841
transform 1 0 1820 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1712256841
transform 1 0 1780 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1712256841
transform 1 0 2268 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1712256841
transform 1 0 2164 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1712256841
transform 1 0 2332 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1712256841
transform 1 0 2116 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1712256841
transform 1 0 2404 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1712256841
transform 1 0 2324 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1712256841
transform 1 0 2300 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2599
timestamp 1712256841
transform 1 0 2404 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1712256841
transform 1 0 2340 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1712256841
transform 1 0 2196 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1712256841
transform 1 0 2164 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1712256841
transform 1 0 2084 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1712256841
transform 1 0 2100 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1712256841
transform 1 0 1908 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1712256841
transform 1 0 1860 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1712256841
transform 1 0 1500 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1712256841
transform 1 0 1116 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1712256841
transform 1 0 1108 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1712256841
transform 1 0 1020 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1712256841
transform 1 0 1140 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1712256841
transform 1 0 1052 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1712256841
transform 1 0 1028 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1712256841
transform 1 0 892 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1712256841
transform 1 0 428 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1712256841
transform 1 0 332 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1712256841
transform 1 0 1604 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1712256841
transform 1 0 1540 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1712256841
transform 1 0 2236 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1712256841
transform 1 0 1564 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1712256841
transform 1 0 2492 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1712256841
transform 1 0 2388 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1712256841
transform 1 0 2388 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1712256841
transform 1 0 2220 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1712256841
transform 1 0 2284 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1712256841
transform 1 0 2236 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1712256841
transform 1 0 2180 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1712256841
transform 1 0 1740 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1712256841
transform 1 0 1708 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1712256841
transform 1 0 1604 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1712256841
transform 1 0 1620 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1712256841
transform 1 0 1420 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1712256841
transform 1 0 1420 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1712256841
transform 1 0 1380 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1712256841
transform 1 0 1812 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1712256841
transform 1 0 1708 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1712256841
transform 1 0 1708 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1712256841
transform 1 0 1516 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1712256841
transform 1 0 1660 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1712256841
transform 1 0 1548 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1712256841
transform 1 0 1516 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1712256841
transform 1 0 644 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1712256841
transform 1 0 580 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1712256841
transform 1 0 548 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1712256841
transform 1 0 612 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1712256841
transform 1 0 500 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1712256841
transform 1 0 460 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1712256841
transform 1 0 436 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1712256841
transform 1 0 436 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1712256841
transform 1 0 420 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1712256841
transform 1 0 668 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1712256841
transform 1 0 444 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1712256841
transform 1 0 796 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1712256841
transform 1 0 684 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1712256841
transform 1 0 916 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1712256841
transform 1 0 796 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1712256841
transform 1 0 820 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1712256841
transform 1 0 780 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1712256841
transform 1 0 2964 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1712256841
transform 1 0 2964 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1712256841
transform 1 0 2844 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1712256841
transform 1 0 2580 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1712256841
transform 1 0 2516 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1712256841
transform 1 0 2516 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1712256841
transform 1 0 2476 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1712256841
transform 1 0 1708 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1712256841
transform 1 0 1708 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1712256841
transform 1 0 1652 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1712256841
transform 1 0 1652 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1712256841
transform 1 0 1516 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1712256841
transform 1 0 2596 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1712256841
transform 1 0 2540 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1712256841
transform 1 0 1708 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1712256841
transform 1 0 1708 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1712256841
transform 1 0 1684 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1712256841
transform 1 0 484 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1712256841
transform 1 0 444 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1712256841
transform 1 0 404 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1712256841
transform 1 0 444 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1712256841
transform 1 0 420 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1712256841
transform 1 0 420 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1712256841
transform 1 0 388 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1712256841
transform 1 0 980 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1712256841
transform 1 0 516 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1712256841
transform 1 0 484 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1712256841
transform 1 0 436 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1712256841
transform 1 0 1124 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1712256841
transform 1 0 1012 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1712256841
transform 1 0 972 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1712256841
transform 1 0 500 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1712256841
transform 1 0 412 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1712256841
transform 1 0 1780 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1712256841
transform 1 0 1636 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1712256841
transform 1 0 1748 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1712256841
transform 1 0 1668 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1712256841
transform 1 0 1748 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1712256841
transform 1 0 1716 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1712256841
transform 1 0 1748 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1712256841
transform 1 0 1588 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1712256841
transform 1 0 1572 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1712256841
transform 1 0 1468 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1712256841
transform 1 0 1468 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1712256841
transform 1 0 1372 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1712256841
transform 1 0 1356 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1712256841
transform 1 0 1348 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1712256841
transform 1 0 1348 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1712256841
transform 1 0 1260 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1712256841
transform 1 0 1252 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1712256841
transform 1 0 932 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1712256841
transform 1 0 596 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1712256841
transform 1 0 1548 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1712256841
transform 1 0 1348 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1712256841
transform 1 0 1332 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1712256841
transform 1 0 1580 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1712256841
transform 1 0 1388 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1712256841
transform 1 0 1300 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1712256841
transform 1 0 1300 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2718
timestamp 1712256841
transform 1 0 1044 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1712256841
transform 1 0 1044 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1712256841
transform 1 0 996 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1712256841
transform 1 0 748 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1712256841
transform 1 0 748 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1712256841
transform 1 0 644 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1712256841
transform 1 0 156 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1712256841
transform 1 0 2140 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1712256841
transform 1 0 1820 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1712256841
transform 1 0 2500 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1712256841
transform 1 0 2324 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1712256841
transform 1 0 2124 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1712256841
transform 1 0 2380 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1712256841
transform 1 0 2340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1712256841
transform 1 0 2132 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1712256841
transform 1 0 2588 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1712256841
transform 1 0 2244 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1712256841
transform 1 0 2172 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1712256841
transform 1 0 2548 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1712256841
transform 1 0 2140 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1712256841
transform 1 0 1836 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1712256841
transform 1 0 1828 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1712256841
transform 1 0 1724 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1712256841
transform 1 0 1924 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1712256841
transform 1 0 1732 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2743
timestamp 1712256841
transform 1 0 1652 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1712256841
transform 1 0 1316 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1712256841
transform 1 0 2548 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1712256841
transform 1 0 1828 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1712256841
transform 1 0 1804 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1712256841
transform 1 0 1372 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1712256841
transform 1 0 2156 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1712256841
transform 1 0 1884 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1712256841
transform 1 0 1876 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1712256841
transform 1 0 1844 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1712256841
transform 1 0 1844 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1712256841
transform 1 0 1796 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1712256841
transform 1 0 1796 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1712256841
transform 1 0 1772 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2757
timestamp 1712256841
transform 1 0 1756 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1712256841
transform 1 0 1748 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1712256841
transform 1 0 1692 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1712256841
transform 1 0 1692 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1712256841
transform 1 0 1556 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1712256841
transform 1 0 1980 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2763
timestamp 1712256841
transform 1 0 1900 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1712256841
transform 1 0 2148 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1712256841
transform 1 0 2084 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1712256841
transform 1 0 1972 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2767
timestamp 1712256841
transform 1 0 1980 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1712256841
transform 1 0 1868 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1712256841
transform 1 0 1772 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1712256841
transform 1 0 2636 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1712256841
transform 1 0 2524 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1712256841
transform 1 0 2620 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1712256841
transform 1 0 2508 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1712256841
transform 1 0 2548 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1712256841
transform 1 0 2500 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1712256841
transform 1 0 2356 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1712256841
transform 1 0 2660 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1712256841
transform 1 0 2508 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1712256841
transform 1 0 2420 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1712256841
transform 1 0 1596 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1712256841
transform 1 0 1508 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1712256841
transform 1 0 1484 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1712256841
transform 1 0 1460 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1712256841
transform 1 0 1460 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1712256841
transform 1 0 948 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1712256841
transform 1 0 884 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1712256841
transform 1 0 588 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1712256841
transform 1 0 924 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1712256841
transform 1 0 884 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1712256841
transform 1 0 868 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1712256841
transform 1 0 588 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1712256841
transform 1 0 1556 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1712256841
transform 1 0 924 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1712256841
transform 1 0 1556 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1712256841
transform 1 0 1028 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1712256841
transform 1 0 1100 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1712256841
transform 1 0 972 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1712256841
transform 1 0 932 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1712256841
transform 1 0 1212 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1712256841
transform 1 0 1052 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1712256841
transform 1 0 1052 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1712256841
transform 1 0 1020 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1712256841
transform 1 0 2548 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1712256841
transform 1 0 2524 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1712256841
transform 1 0 1548 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1712256841
transform 1 0 532 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2807
timestamp 1712256841
transform 1 0 484 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1712256841
transform 1 0 580 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1712256841
transform 1 0 524 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1712256841
transform 1 0 668 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1712256841
transform 1 0 564 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1712256841
transform 1 0 500 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1712256841
transform 1 0 628 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1712256841
transform 1 0 556 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1712256841
transform 1 0 500 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2816
timestamp 1712256841
transform 1 0 468 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1712256841
transform 1 0 652 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1712256841
transform 1 0 540 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1712256841
transform 1 0 1004 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1712256841
transform 1 0 868 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1712256841
transform 1 0 884 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1712256841
transform 1 0 724 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1712256841
transform 1 0 732 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1712256841
transform 1 0 628 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1712256841
transform 1 0 1076 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1712256841
transform 1 0 1052 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2827
timestamp 1712256841
transform 1 0 1996 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2828
timestamp 1712256841
transform 1 0 1988 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1712256841
transform 1 0 1820 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1712256841
transform 1 0 1572 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1712256841
transform 1 0 1572 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1712256841
transform 1 0 1404 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1712256841
transform 1 0 1316 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1712256841
transform 1 0 1308 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1712256841
transform 1 0 1252 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2836
timestamp 1712256841
transform 1 0 1244 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1712256841
transform 1 0 612 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1712256841
transform 1 0 508 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1712256841
transform 1 0 596 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2840
timestamp 1712256841
transform 1 0 508 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1712256841
transform 1 0 692 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1712256841
transform 1 0 612 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1712256841
transform 1 0 1572 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1712256841
transform 1 0 1572 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1712256841
transform 1 0 2124 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2846
timestamp 1712256841
transform 1 0 1596 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1712256841
transform 1 0 1732 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1712256841
transform 1 0 1588 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1712256841
transform 1 0 2396 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1712256841
transform 1 0 1708 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1712256841
transform 1 0 1956 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1712256841
transform 1 0 1748 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1712256841
transform 1 0 2028 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1712256841
transform 1 0 1924 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1712256841
transform 1 0 1972 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1712256841
transform 1 0 1820 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1712256841
transform 1 0 2276 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1712256841
transform 1 0 2244 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1712256841
transform 1 0 2212 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1712256841
transform 1 0 2124 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1712256841
transform 1 0 1980 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1712256841
transform 1 0 1948 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1712256841
transform 1 0 1564 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1712256841
transform 1 0 1444 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1712256841
transform 1 0 2436 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1712256841
transform 1 0 2420 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1712256841
transform 1 0 2388 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1712256841
transform 1 0 2012 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1712256841
transform 1 0 2476 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1712256841
transform 1 0 2412 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2871
timestamp 1712256841
transform 1 0 2412 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1712256841
transform 1 0 2356 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2873
timestamp 1712256841
transform 1 0 2140 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1712256841
transform 1 0 2404 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1712256841
transform 1 0 2356 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2876
timestamp 1712256841
transform 1 0 2132 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1712256841
transform 1 0 2452 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1712256841
transform 1 0 2268 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1712256841
transform 1 0 2084 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1712256841
transform 1 0 2356 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1712256841
transform 1 0 2108 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1712256841
transform 1 0 2180 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1712256841
transform 1 0 2132 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1712256841
transform 1 0 2100 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1712256841
transform 1 0 1996 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1712256841
transform 1 0 2260 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1712256841
transform 1 0 2220 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1712256841
transform 1 0 2476 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1712256841
transform 1 0 2452 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1712256841
transform 1 0 2452 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1712256841
transform 1 0 2332 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1712256841
transform 1 0 1532 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1712256841
transform 1 0 1260 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1712256841
transform 1 0 1628 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1712256841
transform 1 0 1548 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1712256841
transform 1 0 1748 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1712256841
transform 1 0 1668 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1712256841
transform 1 0 1668 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1712256841
transform 1 0 1628 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1712256841
transform 1 0 1636 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1712256841
transform 1 0 1540 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1712256841
transform 1 0 1332 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1712256841
transform 1 0 1228 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1712256841
transform 1 0 1068 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1712256841
transform 1 0 1268 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1712256841
transform 1 0 1156 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1712256841
transform 1 0 1124 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1712256841
transform 1 0 1476 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1712256841
transform 1 0 1388 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1712256841
transform 1 0 1388 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1712256841
transform 1 0 1196 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1712256841
transform 1 0 1196 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1712256841
transform 1 0 1028 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1712256841
transform 1 0 604 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1712256841
transform 1 0 564 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1712256841
transform 1 0 156 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1712256841
transform 1 0 1964 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1712256841
transform 1 0 1940 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1712256841
transform 1 0 1932 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1712256841
transform 1 0 1388 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1712256841
transform 1 0 1404 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1712256841
transform 1 0 772 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1712256841
transform 1 0 708 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1712256841
transform 1 0 668 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1712256841
transform 1 0 908 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1712256841
transform 1 0 812 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1712256841
transform 1 0 1284 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1712256841
transform 1 0 1284 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1712256841
transform 1 0 1244 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1712256841
transform 1 0 1244 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1712256841
transform 1 0 972 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1712256841
transform 1 0 972 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1712256841
transform 1 0 924 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1712256841
transform 1 0 868 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1712256841
transform 1 0 812 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1712256841
transform 1 0 812 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1712256841
transform 1 0 332 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1712256841
transform 1 0 332 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1712256841
transform 1 0 268 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1712256841
transform 1 0 1092 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1712256841
transform 1 0 1028 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1712256841
transform 1 0 916 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1712256841
transform 1 0 916 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1712256841
transform 1 0 860 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1712256841
transform 1 0 924 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1712256841
transform 1 0 756 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1712256841
transform 1 0 772 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1712256841
transform 1 0 700 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1712256841
transform 1 0 988 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1712256841
transform 1 0 844 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1712256841
transform 1 0 740 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1712256841
transform 1 0 644 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1712256841
transform 1 0 644 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1712256841
transform 1 0 604 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1712256841
transform 1 0 740 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2956
timestamp 1712256841
transform 1 0 700 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1712256841
transform 1 0 668 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1712256841
transform 1 0 604 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1712256841
transform 1 0 1156 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1712256841
transform 1 0 1060 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2961
timestamp 1712256841
transform 1 0 996 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1712256841
transform 1 0 916 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2963
timestamp 1712256841
transform 1 0 1356 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1712256841
transform 1 0 1268 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1712256841
transform 1 0 1268 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1712256841
transform 1 0 1060 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1712256841
transform 1 0 1044 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1712256841
transform 1 0 980 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1712256841
transform 1 0 756 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1712256841
transform 1 0 708 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1712256841
transform 1 0 644 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1712256841
transform 1 0 580 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2973
timestamp 1712256841
transform 1 0 836 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1712256841
transform 1 0 780 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1712256841
transform 1 0 772 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1712256841
transform 1 0 700 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1712256841
transform 1 0 524 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1712256841
transform 1 0 964 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1712256841
transform 1 0 884 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1712256841
transform 1 0 628 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1712256841
transform 1 0 2524 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1712256841
transform 1 0 2492 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1712256841
transform 1 0 2412 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1712256841
transform 1 0 2380 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1712256841
transform 1 0 2380 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1712256841
transform 1 0 1468 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1712256841
transform 1 0 1164 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1712256841
transform 1 0 1156 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1712256841
transform 1 0 1148 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1712256841
transform 1 0 1148 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1712256841
transform 1 0 1052 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1712256841
transform 1 0 1004 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1712256841
transform 1 0 652 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1712256841
transform 1 0 1084 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2995
timestamp 1712256841
transform 1 0 940 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2996
timestamp 1712256841
transform 1 0 700 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2997
timestamp 1712256841
transform 1 0 636 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1712256841
transform 1 0 852 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1712256841
transform 1 0 804 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1712256841
transform 1 0 764 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1712256841
transform 1 0 580 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1712256841
transform 1 0 852 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1712256841
transform 1 0 700 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1712256841
transform 1 0 692 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1712256841
transform 1 0 612 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1712256841
transform 1 0 564 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1712256841
transform 1 0 2084 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1712256841
transform 1 0 1940 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3009
timestamp 1712256841
transform 1 0 2452 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1712256841
transform 1 0 1932 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1712256841
transform 1 0 1956 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1712256841
transform 1 0 1924 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3013
timestamp 1712256841
transform 1 0 1956 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1712256841
transform 1 0 1884 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1712256841
transform 1 0 1900 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1712256841
transform 1 0 1452 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1712256841
transform 1 0 2252 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1712256841
transform 1 0 2244 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3019
timestamp 1712256841
transform 1 0 1868 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1712256841
transform 1 0 1868 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1712256841
transform 1 0 1828 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1712256841
transform 1 0 1780 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1712256841
transform 1 0 1764 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3024
timestamp 1712256841
transform 1 0 1764 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1712256841
transform 1 0 1764 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1712256841
transform 1 0 1724 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1712256841
transform 1 0 1724 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1712256841
transform 1 0 1620 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1712256841
transform 1 0 1428 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1712256841
transform 1 0 1420 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3031
timestamp 1712256841
transform 1 0 1484 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1712256841
transform 1 0 1468 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1712256841
transform 1 0 1388 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1712256841
transform 1 0 1380 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1712256841
transform 1 0 1276 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1712256841
transform 1 0 1220 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1712256841
transform 1 0 1500 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1712256841
transform 1 0 1412 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1712256841
transform 1 0 1212 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3040
timestamp 1712256841
transform 1 0 1196 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1712256841
transform 1 0 1188 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1712256841
transform 1 0 1124 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1712256841
transform 1 0 1092 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1712256841
transform 1 0 1084 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1712256841
transform 1 0 2228 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1712256841
transform 1 0 1988 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1712256841
transform 1 0 2516 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1712256841
transform 1 0 2460 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3049
timestamp 1712256841
transform 1 0 2460 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1712256841
transform 1 0 2372 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3051
timestamp 1712256841
transform 1 0 2188 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1712256841
transform 1 0 2188 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1712256841
transform 1 0 2084 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1712256841
transform 1 0 2084 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1712256841
transform 1 0 2060 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1712256841
transform 1 0 2060 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1712256841
transform 1 0 1612 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1712256841
transform 1 0 1612 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1712256841
transform 1 0 1572 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1712256841
transform 1 0 2244 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1712256841
transform 1 0 2188 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1712256841
transform 1 0 2180 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1712256841
transform 1 0 1932 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1712256841
transform 1 0 1908 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1712256841
transform 1 0 1908 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1712256841
transform 1 0 1908 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1712256841
transform 1 0 1828 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1712256841
transform 1 0 2076 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1712256841
transform 1 0 1940 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1712256841
transform 1 0 1932 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1712256841
transform 1 0 1900 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1712256841
transform 1 0 1852 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1712256841
transform 1 0 1956 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1712256841
transform 1 0 1844 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1712256841
transform 1 0 1732 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1712256841
transform 1 0 1620 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1712256841
transform 1 0 1588 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1712256841
transform 1 0 2612 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1712256841
transform 1 0 2588 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1712256841
transform 1 0 2580 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1712256841
transform 1 0 2460 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1712256841
transform 1 0 2428 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1712256841
transform 1 0 2404 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1712256841
transform 1 0 2452 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1712256841
transform 1 0 2444 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1712256841
transform 1 0 2372 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1712256841
transform 1 0 2356 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1712256841
transform 1 0 2316 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1712256841
transform 1 0 2284 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1712256841
transform 1 0 2676 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1712256841
transform 1 0 2628 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1712256841
transform 1 0 2524 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1712256841
transform 1 0 2508 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1712256841
transform 1 0 2508 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1712256841
transform 1 0 2436 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1712256841
transform 1 0 2412 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1712256841
transform 1 0 3068 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1712256841
transform 1 0 3012 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1712256841
transform 1 0 2932 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1712256841
transform 1 0 2916 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1712256841
transform 1 0 2548 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1712256841
transform 1 0 2548 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1712256841
transform 1 0 2540 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1712256841
transform 1 0 2276 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1712256841
transform 1 0 2244 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1712256841
transform 1 0 2236 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1712256841
transform 1 0 2236 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1712256841
transform 1 0 2236 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1712256841
transform 1 0 2180 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1712256841
transform 1 0 2092 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1712256841
transform 1 0 2044 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1712256841
transform 1 0 2020 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1712256841
transform 1 0 2060 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1712256841
transform 1 0 1972 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1712256841
transform 1 0 1924 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1712256841
transform 1 0 1860 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1712256841
transform 1 0 1780 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1712256841
transform 1 0 1724 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1712256841
transform 1 0 2228 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1712256841
transform 1 0 2220 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1712256841
transform 1 0 2212 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1712256841
transform 1 0 2092 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1712256841
transform 1 0 2076 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1712256841
transform 1 0 2076 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1712256841
transform 1 0 2060 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1712256841
transform 1 0 2028 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1712256841
transform 1 0 1716 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1712256841
transform 1 0 1660 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1712256841
transform 1 0 1700 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1712256841
transform 1 0 1660 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1712256841
transform 1 0 1636 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1712256841
transform 1 0 1612 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1712256841
transform 1 0 3236 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1712256841
transform 1 0 1916 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1712256841
transform 1 0 1908 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1712256841
transform 1 0 1604 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1712256841
transform 1 0 1596 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1712256841
transform 1 0 1388 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1712256841
transform 1 0 1596 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3140
timestamp 1712256841
transform 1 0 1596 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1712256841
transform 1 0 1572 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1712256841
transform 1 0 1572 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1712256841
transform 1 0 1836 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1712256841
transform 1 0 1604 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1712256841
transform 1 0 1548 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1712256841
transform 1 0 372 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1712256841
transform 1 0 1580 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1712256841
transform 1 0 1428 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1712256841
transform 1 0 1468 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1712256841
transform 1 0 1428 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1712256841
transform 1 0 1468 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1712256841
transform 1 0 1420 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1712256841
transform 1 0 1380 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1712256841
transform 1 0 772 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1712256841
transform 1 0 540 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1712256841
transform 1 0 420 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1712256841
transform 1 0 484 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1712256841
transform 1 0 412 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1712256841
transform 1 0 428 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1712256841
transform 1 0 356 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1712256841
transform 1 0 1444 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1712256841
transform 1 0 1340 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1712256841
transform 1 0 1284 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1712256841
transform 1 0 2044 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1712256841
transform 1 0 1996 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3166
timestamp 1712256841
transform 1 0 1996 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1712256841
transform 1 0 1532 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1712256841
transform 1 0 372 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1712256841
transform 1 0 348 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1712256841
transform 1 0 436 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1712256841
transform 1 0 340 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1712256841
transform 1 0 404 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3173
timestamp 1712256841
transform 1 0 404 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1712256841
transform 1 0 324 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1712256841
transform 1 0 316 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1712256841
transform 1 0 428 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1712256841
transform 1 0 348 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1712256841
transform 1 0 468 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1712256841
transform 1 0 404 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3180
timestamp 1712256841
transform 1 0 356 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1712256841
transform 1 0 436 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1712256841
transform 1 0 332 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1712256841
transform 1 0 524 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1712256841
transform 1 0 340 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1712256841
transform 1 0 420 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3186
timestamp 1712256841
transform 1 0 340 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1712256841
transform 1 0 2684 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1712256841
transform 1 0 1892 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1712256841
transform 1 0 2892 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1712256841
transform 1 0 2660 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1712256841
transform 1 0 2684 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1712256841
transform 1 0 2620 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1712256841
transform 1 0 2588 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3194
timestamp 1712256841
transform 1 0 2228 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1712256841
transform 1 0 2628 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1712256841
transform 1 0 2412 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3197
timestamp 1712256841
transform 1 0 2268 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1712256841
transform 1 0 2644 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1712256841
transform 1 0 2476 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1712256841
transform 1 0 2452 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1712256841
transform 1 0 2148 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1712256841
transform 1 0 1916 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1712256841
transform 1 0 2428 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1712256841
transform 1 0 2308 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1712256841
transform 1 0 2132 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3206
timestamp 1712256841
transform 1 0 2236 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1712256841
transform 1 0 2196 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1712256841
transform 1 0 1940 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1712256841
transform 1 0 1820 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1712256841
transform 1 0 1852 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1712256841
transform 1 0 1788 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1712256841
transform 1 0 1732 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1712256841
transform 1 0 1732 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1712256841
transform 1 0 2028 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1712256841
transform 1 0 1572 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1712256841
transform 1 0 1588 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1712256841
transform 1 0 1292 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1712256841
transform 1 0 1276 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3219
timestamp 1712256841
transform 1 0 1108 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3220
timestamp 1712256841
transform 1 0 1124 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3221
timestamp 1712256841
transform 1 0 940 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1712256841
transform 1 0 2484 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3223
timestamp 1712256841
transform 1 0 2060 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1712256841
transform 1 0 2508 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1712256841
transform 1 0 2212 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1712256841
transform 1 0 2132 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1712256841
transform 1 0 1804 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3228
timestamp 1712256841
transform 1 0 1700 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1712256841
transform 1 0 1372 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1712256841
transform 1 0 204 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1712256841
transform 1 0 1356 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1712256841
transform 1 0 684 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1712256841
transform 1 0 1628 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3234
timestamp 1712256841
transform 1 0 1372 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3235
timestamp 1712256841
transform 1 0 1988 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1712256841
transform 1 0 1660 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1712256841
transform 1 0 2164 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3238
timestamp 1712256841
transform 1 0 1644 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1712256841
transform 1 0 1660 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3240
timestamp 1712256841
transform 1 0 1620 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3241
timestamp 1712256841
transform 1 0 1724 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1712256841
transform 1 0 1604 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1712256841
transform 1 0 1644 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3244
timestamp 1712256841
transform 1 0 1524 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1712256841
transform 1 0 1204 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1712256841
transform 1 0 1148 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3247
timestamp 1712256841
transform 1 0 1100 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3248
timestamp 1712256841
transform 1 0 2132 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1712256841
transform 1 0 2116 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1712256841
transform 1 0 2012 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1712256841
transform 1 0 2220 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1712256841
transform 1 0 2196 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1712256841
transform 1 0 2244 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1712256841
transform 1 0 2204 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1712256841
transform 1 0 2228 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1712256841
transform 1 0 2148 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1712256841
transform 1 0 2028 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1712256841
transform 1 0 1980 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1712256841
transform 1 0 2244 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1712256841
transform 1 0 1980 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1712256841
transform 1 0 2108 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1712256841
transform 1 0 2052 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1712256841
transform 1 0 2036 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1712256841
transform 1 0 1964 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3265
timestamp 1712256841
transform 1 0 2148 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1712256841
transform 1 0 1996 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1712256841
transform 1 0 2020 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1712256841
transform 1 0 1820 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1712256841
transform 1 0 2476 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1712256841
transform 1 0 2196 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1712256841
transform 1 0 2196 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1712256841
transform 1 0 2068 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1712256841
transform 1 0 2332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1712256841
transform 1 0 2284 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1712256841
transform 1 0 2172 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1712256841
transform 1 0 2116 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1712256841
transform 1 0 2020 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1712256841
transform 1 0 2036 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1712256841
transform 1 0 1892 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1712256841
transform 1 0 668 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1712256841
transform 1 0 316 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1712256841
transform 1 0 260 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1712256841
transform 1 0 108 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1712256841
transform 1 0 276 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1712256841
transform 1 0 220 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1712256841
transform 1 0 228 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1712256841
transform 1 0 164 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1712256841
transform 1 0 164 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1712256841
transform 1 0 116 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3290
timestamp 1712256841
transform 1 0 812 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1712256841
transform 1 0 708 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3292
timestamp 1712256841
transform 1 0 724 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1712256841
transform 1 0 524 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1712256841
transform 1 0 540 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1712256841
transform 1 0 196 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1712256841
transform 1 0 260 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1712256841
transform 1 0 116 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1712256841
transform 1 0 1140 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1712256841
transform 1 0 132 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1712256841
transform 1 0 132 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1712256841
transform 1 0 84 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3302
timestamp 1712256841
transform 1 0 604 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1712256841
transform 1 0 476 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1712256841
transform 1 0 268 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3305
timestamp 1712256841
transform 1 0 148 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3306
timestamp 1712256841
transform 1 0 116 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1712256841
transform 1 0 148 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1712256841
transform 1 0 100 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3309
timestamp 1712256841
transform 1 0 108 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1712256841
transform 1 0 84 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1712256841
transform 1 0 1796 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1712256841
transform 1 0 1684 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3313
timestamp 1712256841
transform 1 0 1652 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3314
timestamp 1712256841
transform 1 0 1436 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3315
timestamp 1712256841
transform 1 0 3156 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3316
timestamp 1712256841
transform 1 0 1724 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1712256841
transform 1 0 1700 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3318
timestamp 1712256841
transform 1 0 1452 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1712256841
transform 1 0 1388 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3320
timestamp 1712256841
transform 1 0 1372 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3321
timestamp 1712256841
transform 1 0 1276 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3322
timestamp 1712256841
transform 1 0 1276 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3323
timestamp 1712256841
transform 1 0 820 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3324
timestamp 1712256841
transform 1 0 1420 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1712256841
transform 1 0 364 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1712256841
transform 1 0 380 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3327
timestamp 1712256841
transform 1 0 348 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1712256841
transform 1 0 1036 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1712256841
transform 1 0 492 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3330
timestamp 1712256841
transform 1 0 492 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3331
timestamp 1712256841
transform 1 0 316 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3332
timestamp 1712256841
transform 1 0 404 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3333
timestamp 1712256841
transform 1 0 348 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3334
timestamp 1712256841
transform 1 0 348 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1712256841
transform 1 0 292 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3336
timestamp 1712256841
transform 1 0 428 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3337
timestamp 1712256841
transform 1 0 308 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3338
timestamp 1712256841
transform 1 0 1660 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3339
timestamp 1712256841
transform 1 0 1500 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1712256841
transform 1 0 1428 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3341
timestamp 1712256841
transform 1 0 1428 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1712256841
transform 1 0 796 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3343
timestamp 1712256841
transform 1 0 548 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1712256841
transform 1 0 1964 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3345
timestamp 1712256841
transform 1 0 1732 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3346
timestamp 1712256841
transform 1 0 1732 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1712256841
transform 1 0 564 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1712256841
transform 1 0 276 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1712256841
transform 1 0 228 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1712256841
transform 1 0 364 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3351
timestamp 1712256841
transform 1 0 332 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3352
timestamp 1712256841
transform 1 0 356 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1712256841
transform 1 0 300 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3354
timestamp 1712256841
transform 1 0 380 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3355
timestamp 1712256841
transform 1 0 348 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1712256841
transform 1 0 284 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1712256841
transform 1 0 2148 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1712256841
transform 1 0 2100 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1712256841
transform 1 0 1676 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3360
timestamp 1712256841
transform 1 0 1668 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1712256841
transform 1 0 748 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1712256841
transform 1 0 2076 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3363
timestamp 1712256841
transform 1 0 2036 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1712256841
transform 1 0 2036 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1712256841
transform 1 0 860 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3366
timestamp 1712256841
transform 1 0 844 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1712256841
transform 1 0 828 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3368
timestamp 1712256841
transform 1 0 372 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3369
timestamp 1712256841
transform 1 0 252 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1712256841
transform 1 0 212 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3371
timestamp 1712256841
transform 1 0 2116 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1712256841
transform 1 0 2116 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1712256841
transform 1 0 2036 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1712256841
transform 1 0 572 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_3375
timestamp 1712256841
transform 1 0 852 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1712256841
transform 1 0 756 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3377
timestamp 1712256841
transform 1 0 756 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3378
timestamp 1712256841
transform 1 0 588 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3379
timestamp 1712256841
transform 1 0 436 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3380
timestamp 1712256841
transform 1 0 260 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3381
timestamp 1712256841
transform 1 0 228 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3382
timestamp 1712256841
transform 1 0 1020 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3383
timestamp 1712256841
transform 1 0 1012 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3384
timestamp 1712256841
transform 1 0 932 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3385
timestamp 1712256841
transform 1 0 932 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3386
timestamp 1712256841
transform 1 0 828 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3387
timestamp 1712256841
transform 1 0 572 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1712256841
transform 1 0 780 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3389
timestamp 1712256841
transform 1 0 676 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1712256841
transform 1 0 652 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3391
timestamp 1712256841
transform 1 0 556 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1712256841
transform 1 0 556 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1712256841
transform 1 0 516 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3394
timestamp 1712256841
transform 1 0 508 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3395
timestamp 1712256841
transform 1 0 772 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3396
timestamp 1712256841
transform 1 0 748 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3397
timestamp 1712256841
transform 1 0 748 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3398
timestamp 1712256841
transform 1 0 668 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3399
timestamp 1712256841
transform 1 0 636 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3400
timestamp 1712256841
transform 1 0 564 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3401
timestamp 1712256841
transform 1 0 1476 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3402
timestamp 1712256841
transform 1 0 1436 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1712256841
transform 1 0 1988 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3404
timestamp 1712256841
transform 1 0 1620 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3405
timestamp 1712256841
transform 1 0 1548 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3406
timestamp 1712256841
transform 1 0 1548 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3407
timestamp 1712256841
transform 1 0 1460 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3408
timestamp 1712256841
transform 1 0 1484 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3409
timestamp 1712256841
transform 1 0 1380 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3410
timestamp 1712256841
transform 1 0 1340 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3411
timestamp 1712256841
transform 1 0 892 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3412
timestamp 1712256841
transform 1 0 884 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3413
timestamp 1712256841
transform 1 0 836 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1712256841
transform 1 0 644 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3415
timestamp 1712256841
transform 1 0 324 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3416
timestamp 1712256841
transform 1 0 324 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1712256841
transform 1 0 140 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3418
timestamp 1712256841
transform 1 0 140 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3419
timestamp 1712256841
transform 1 0 116 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_3420
timestamp 1712256841
transform 1 0 1476 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3421
timestamp 1712256841
transform 1 0 1452 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1712256841
transform 1 0 1628 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1712256841
transform 1 0 1532 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3424
timestamp 1712256841
transform 1 0 1428 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3425
timestamp 1712256841
transform 1 0 1444 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3426
timestamp 1712256841
transform 1 0 1364 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3427
timestamp 1712256841
transform 1 0 2332 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3428
timestamp 1712256841
transform 1 0 2140 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3429
timestamp 1712256841
transform 1 0 2132 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1712256841
transform 1 0 1780 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3431
timestamp 1712256841
transform 1 0 1804 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3432
timestamp 1712256841
transform 1 0 1764 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3433
timestamp 1712256841
transform 1 0 1836 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1712256841
transform 1 0 1788 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3435
timestamp 1712256841
transform 1 0 1972 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1712256841
transform 1 0 1828 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3437
timestamp 1712256841
transform 1 0 1860 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3438
timestamp 1712256841
transform 1 0 1396 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1712256841
transform 1 0 1468 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1712256841
transform 1 0 1412 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3441
timestamp 1712256841
transform 1 0 1308 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1712256841
transform 1 0 1348 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3443
timestamp 1712256841
transform 1 0 1220 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1712256841
transform 1 0 1828 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3445
timestamp 1712256841
transform 1 0 1788 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3446
timestamp 1712256841
transform 1 0 1780 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1712256841
transform 1 0 1780 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3448
timestamp 1712256841
transform 1 0 1732 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1712256841
transform 1 0 1540 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3450
timestamp 1712256841
transform 1 0 1540 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3451
timestamp 1712256841
transform 1 0 1300 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1712256841
transform 1 0 1300 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3453
timestamp 1712256841
transform 1 0 1004 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1712256841
transform 1 0 2412 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1712256841
transform 1 0 1988 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1712256841
transform 1 0 2436 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3457
timestamp 1712256841
transform 1 0 2340 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3458
timestamp 1712256841
transform 1 0 2484 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1712256841
transform 1 0 2452 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1712256841
transform 1 0 2436 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1712256841
transform 1 0 2428 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3462
timestamp 1712256841
transform 1 0 2428 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1712256841
transform 1 0 2396 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1712256841
transform 1 0 2372 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3465
timestamp 1712256841
transform 1 0 2364 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1712256841
transform 1 0 2356 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1712256841
transform 1 0 2036 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1712256841
transform 1 0 2564 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3469
timestamp 1712256841
transform 1 0 2540 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1712256841
transform 1 0 1852 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3471
timestamp 1712256841
transform 1 0 1788 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3472
timestamp 1712256841
transform 1 0 2276 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1712256841
transform 1 0 1772 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3474
timestamp 1712256841
transform 1 0 1820 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1712256841
transform 1 0 1788 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3476
timestamp 1712256841
transform 1 0 1908 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3477
timestamp 1712256841
transform 1 0 1844 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1712256841
transform 1 0 1844 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3479
timestamp 1712256841
transform 1 0 1804 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3480
timestamp 1712256841
transform 1 0 2020 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3481
timestamp 1712256841
transform 1 0 1892 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3482
timestamp 1712256841
transform 1 0 1844 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3483
timestamp 1712256841
transform 1 0 1844 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1712256841
transform 1 0 2852 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3485
timestamp 1712256841
transform 1 0 2564 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1712256841
transform 1 0 2524 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3487
timestamp 1712256841
transform 1 0 2500 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3488
timestamp 1712256841
transform 1 0 2020 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3489
timestamp 1712256841
transform 1 0 2020 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1712256841
transform 1 0 1972 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3491
timestamp 1712256841
transform 1 0 3084 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3492
timestamp 1712256841
transform 1 0 3036 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3493
timestamp 1712256841
transform 1 0 3012 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3494
timestamp 1712256841
transform 1 0 3012 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3495
timestamp 1712256841
transform 1 0 3012 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3496
timestamp 1712256841
transform 1 0 2604 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3497
timestamp 1712256841
transform 1 0 2580 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3498
timestamp 1712256841
transform 1 0 2572 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1712256841
transform 1 0 2772 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1712256841
transform 1 0 2044 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3501
timestamp 1712256841
transform 1 0 1860 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3502
timestamp 1712256841
transform 1 0 2300 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3503
timestamp 1712256841
transform 1 0 2236 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3504
timestamp 1712256841
transform 1 0 2484 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3505
timestamp 1712256841
transform 1 0 2428 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3506
timestamp 1712256841
transform 1 0 2308 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3507
timestamp 1712256841
transform 1 0 3068 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3508
timestamp 1712256841
transform 1 0 2796 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1712256841
transform 1 0 2636 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3510
timestamp 1712256841
transform 1 0 2636 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3511
timestamp 1712256841
transform 1 0 2604 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3512
timestamp 1712256841
transform 1 0 2508 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1712256841
transform 1 0 2380 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1712256841
transform 1 0 2308 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3515
timestamp 1712256841
transform 1 0 2364 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3516
timestamp 1712256841
transform 1 0 2260 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1712256841
transform 1 0 2228 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3518
timestamp 1712256841
transform 1 0 2404 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3519
timestamp 1712256841
transform 1 0 2284 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3520
timestamp 1712256841
transform 1 0 2180 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3521
timestamp 1712256841
transform 1 0 2836 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3522
timestamp 1712256841
transform 1 0 2764 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3523
timestamp 1712256841
transform 1 0 2700 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3524
timestamp 1712256841
transform 1 0 3140 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3525
timestamp 1712256841
transform 1 0 3004 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1712256841
transform 1 0 1796 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3527
timestamp 1712256841
transform 1 0 1692 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3528
timestamp 1712256841
transform 1 0 1700 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1712256841
transform 1 0 204 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3530
timestamp 1712256841
transform 1 0 140 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1712256841
transform 1 0 108 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3532
timestamp 1712256841
transform 1 0 68 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3533
timestamp 1712256841
transform 1 0 68 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3534
timestamp 1712256841
transform 1 0 156 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3535
timestamp 1712256841
transform 1 0 140 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3536
timestamp 1712256841
transform 1 0 140 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3537
timestamp 1712256841
transform 1 0 100 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3538
timestamp 1712256841
transform 1 0 684 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3539
timestamp 1712256841
transform 1 0 92 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3540
timestamp 1712256841
transform 1 0 140 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3541
timestamp 1712256841
transform 1 0 84 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1712256841
transform 1 0 2196 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3543
timestamp 1712256841
transform 1 0 2156 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3544
timestamp 1712256841
transform 1 0 1716 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1712256841
transform 1 0 1716 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1712256841
transform 1 0 1292 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3547
timestamp 1712256841
transform 1 0 1292 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3548
timestamp 1712256841
transform 1 0 692 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_3549
timestamp 1712256841
transform 1 0 692 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3550
timestamp 1712256841
transform 1 0 524 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3551
timestamp 1712256841
transform 1 0 396 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3552
timestamp 1712256841
transform 1 0 380 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1712256841
transform 1 0 380 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3554
timestamp 1712256841
transform 1 0 324 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3555
timestamp 1712256841
transform 1 0 100 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3556
timestamp 1712256841
transform 1 0 164 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1712256841
transform 1 0 92 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3558
timestamp 1712256841
transform 1 0 1084 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3559
timestamp 1712256841
transform 1 0 1012 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3560
timestamp 1712256841
transform 1 0 748 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1712256841
transform 1 0 164 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1712256841
transform 1 0 84 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3563
timestamp 1712256841
transform 1 0 156 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3564
timestamp 1712256841
transform 1 0 84 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3565
timestamp 1712256841
transform 1 0 172 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3566
timestamp 1712256841
transform 1 0 116 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1712256841
transform 1 0 100 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1712256841
transform 1 0 164 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3569
timestamp 1712256841
transform 1 0 84 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1712256841
transform 1 0 196 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1712256841
transform 1 0 100 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3572
timestamp 1712256841
transform 1 0 516 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3573
timestamp 1712256841
transform 1 0 180 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3574
timestamp 1712256841
transform 1 0 212 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3575
timestamp 1712256841
transform 1 0 108 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3576
timestamp 1712256841
transform 1 0 1220 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3577
timestamp 1712256841
transform 1 0 1124 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1712256841
transform 1 0 1380 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3579
timestamp 1712256841
transform 1 0 1380 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3580
timestamp 1712256841
transform 1 0 1340 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3581
timestamp 1712256841
transform 1 0 1196 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3582
timestamp 1712256841
transform 1 0 1356 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3583
timestamp 1712256841
transform 1 0 1332 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3584
timestamp 1712256841
transform 1 0 1260 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3585
timestamp 1712256841
transform 1 0 1212 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3586
timestamp 1712256841
transform 1 0 1428 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3587
timestamp 1712256841
transform 1 0 1332 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3588
timestamp 1712256841
transform 1 0 1188 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3589
timestamp 1712256841
transform 1 0 1108 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1712256841
transform 1 0 1620 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3591
timestamp 1712256841
transform 1 0 1508 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3592
timestamp 1712256841
transform 1 0 1308 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3593
timestamp 1712256841
transform 1 0 1124 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1712256841
transform 1 0 1956 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_3595
timestamp 1712256841
transform 1 0 1772 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_3596
timestamp 1712256841
transform 1 0 2108 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3597
timestamp 1712256841
transform 1 0 1860 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3598
timestamp 1712256841
transform 1 0 1900 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3599
timestamp 1712256841
transform 1 0 1868 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1712256841
transform 1 0 1852 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1712256841
transform 1 0 1532 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3602
timestamp 1712256841
transform 1 0 1532 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3603
timestamp 1712256841
transform 1 0 1356 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3604
timestamp 1712256841
transform 1 0 2476 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3605
timestamp 1712256841
transform 1 0 2428 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3606
timestamp 1712256841
transform 1 0 2364 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3607
timestamp 1712256841
transform 1 0 2364 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1712256841
transform 1 0 2332 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1712256841
transform 1 0 2044 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1712256841
transform 1 0 2044 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3611
timestamp 1712256841
transform 1 0 2028 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1712256841
transform 1 0 2020 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1712256841
transform 1 0 1980 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1712256841
transform 1 0 1980 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3615
timestamp 1712256841
transform 1 0 1948 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1712256841
transform 1 0 1948 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3617
timestamp 1712256841
transform 1 0 1916 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1712256841
transform 1 0 1892 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1712256841
transform 1 0 1892 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1712256841
transform 1 0 1892 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1712256841
transform 1 0 2100 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3622
timestamp 1712256841
transform 1 0 2020 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1712256841
transform 1 0 1932 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1712256841
transform 1 0 1732 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3625
timestamp 1712256841
transform 1 0 2932 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1712256841
transform 1 0 2612 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3627
timestamp 1712256841
transform 1 0 2540 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3628
timestamp 1712256841
transform 1 0 2540 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3629
timestamp 1712256841
transform 1 0 2500 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3630
timestamp 1712256841
transform 1 0 2468 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3631
timestamp 1712256841
transform 1 0 2468 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1712256841
transform 1 0 2332 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1712256841
transform 1 0 2332 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1712256841
transform 1 0 2188 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1712256841
transform 1 0 2132 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1712256841
transform 1 0 2124 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3637
timestamp 1712256841
transform 1 0 2124 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3638
timestamp 1712256841
transform 1 0 2100 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3639
timestamp 1712256841
transform 1 0 2092 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3640
timestamp 1712256841
transform 1 0 2068 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1712256841
transform 1 0 2068 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3642
timestamp 1712256841
transform 1 0 2060 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1712256841
transform 1 0 1996 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1712256841
transform 1 0 1996 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1712256841
transform 1 0 1988 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3646
timestamp 1712256841
transform 1 0 2196 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3647
timestamp 1712256841
transform 1 0 2164 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3648
timestamp 1712256841
transform 1 0 2164 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1712256841
transform 1 0 2084 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3650
timestamp 1712256841
transform 1 0 1700 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1712256841
transform 1 0 1596 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3652
timestamp 1712256841
transform 1 0 2228 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1712256841
transform 1 0 1724 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1712256841
transform 1 0 1996 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1712256841
transform 1 0 1676 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1712256841
transform 1 0 1580 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1712256841
transform 1 0 1628 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3658
timestamp 1712256841
transform 1 0 1156 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3659
timestamp 1712256841
transform 1 0 1156 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3660
timestamp 1712256841
transform 1 0 1076 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1712256841
transform 1 0 1076 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1712256841
transform 1 0 716 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3663
timestamp 1712256841
transform 1 0 716 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1712256841
transform 1 0 652 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_3665
timestamp 1712256841
transform 1 0 2044 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1712256841
transform 1 0 1932 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3667
timestamp 1712256841
transform 1 0 1852 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1712256841
transform 1 0 1788 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3669
timestamp 1712256841
transform 1 0 1916 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3670
timestamp 1712256841
transform 1 0 1820 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3671
timestamp 1712256841
transform 1 0 1572 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3672
timestamp 1712256841
transform 1 0 1356 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3673
timestamp 1712256841
transform 1 0 1612 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3674
timestamp 1712256841
transform 1 0 1540 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1712256841
transform 1 0 1492 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1712256841
transform 1 0 1460 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3677
timestamp 1712256841
transform 1 0 1516 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3678
timestamp 1712256841
transform 1 0 1460 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3679
timestamp 1712256841
transform 1 0 1300 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3680
timestamp 1712256841
transform 1 0 892 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3681
timestamp 1712256841
transform 1 0 892 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3682
timestamp 1712256841
transform 1 0 868 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1712256841
transform 1 0 868 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3684
timestamp 1712256841
transform 1 0 860 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3685
timestamp 1712256841
transform 1 0 852 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1712256841
transform 1 0 836 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3687
timestamp 1712256841
transform 1 0 812 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1712256841
transform 1 0 532 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3689
timestamp 1712256841
transform 1 0 500 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3690
timestamp 1712256841
transform 1 0 1340 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3691
timestamp 1712256841
transform 1 0 1284 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1712256841
transform 1 0 3156 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1712256841
transform 1 0 2260 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3694
timestamp 1712256841
transform 1 0 2260 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3695
timestamp 1712256841
transform 1 0 1596 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3696
timestamp 1712256841
transform 1 0 1580 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1712256841
transform 1 0 1412 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1712256841
transform 1 0 1356 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3699
timestamp 1712256841
transform 1 0 1660 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3700
timestamp 1712256841
transform 1 0 1292 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3701
timestamp 1712256841
transform 1 0 1252 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3702
timestamp 1712256841
transform 1 0 1236 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3703
timestamp 1712256841
transform 1 0 1228 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3704
timestamp 1712256841
transform 1 0 1164 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3705
timestamp 1712256841
transform 1 0 1268 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3706
timestamp 1712256841
transform 1 0 1236 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1712256841
transform 1 0 1220 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3708
timestamp 1712256841
transform 1 0 1148 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1712256841
transform 1 0 828 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1712256841
transform 1 0 1428 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3711
timestamp 1712256841
transform 1 0 1372 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3712
timestamp 1712256841
transform 1 0 1340 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3713
timestamp 1712256841
transform 1 0 1340 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1712256841
transform 1 0 1204 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1712256841
transform 1 0 1220 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3716
timestamp 1712256841
transform 1 0 1188 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3717
timestamp 1712256841
transform 1 0 1164 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3718
timestamp 1712256841
transform 1 0 1156 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3719
timestamp 1712256841
transform 1 0 1068 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3720
timestamp 1712256841
transform 1 0 1068 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3721
timestamp 1712256841
transform 1 0 748 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3722
timestamp 1712256841
transform 1 0 748 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3723
timestamp 1712256841
transform 1 0 492 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1712256841
transform 1 0 1276 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1712256841
transform 1 0 1116 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3726
timestamp 1712256841
transform 1 0 1372 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1712256841
transform 1 0 1252 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3728
timestamp 1712256841
transform 1 0 1084 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3729
timestamp 1712256841
transform 1 0 1044 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1712256841
transform 1 0 940 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3731
timestamp 1712256841
transform 1 0 924 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1712256841
transform 1 0 908 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1712256841
transform 1 0 636 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1712256841
transform 1 0 636 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3735
timestamp 1712256841
transform 1 0 340 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3736
timestamp 1712256841
transform 1 0 292 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3737
timestamp 1712256841
transform 1 0 284 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1712256841
transform 1 0 1188 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3739
timestamp 1712256841
transform 1 0 1060 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3740
timestamp 1712256841
transform 1 0 1036 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1712256841
transform 1 0 948 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3742
timestamp 1712256841
transform 1 0 916 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3743
timestamp 1712256841
transform 1 0 900 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1712256841
transform 1 0 812 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3745
timestamp 1712256841
transform 1 0 1124 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3746
timestamp 1712256841
transform 1 0 820 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1712256841
transform 1 0 1340 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3748
timestamp 1712256841
transform 1 0 1084 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_3749
timestamp 1712256841
transform 1 0 1156 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3750
timestamp 1712256841
transform 1 0 1092 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3751
timestamp 1712256841
transform 1 0 1084 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3752
timestamp 1712256841
transform 1 0 980 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3753
timestamp 1712256841
transform 1 0 660 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1712256841
transform 1 0 380 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3755
timestamp 1712256841
transform 1 0 316 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3756
timestamp 1712256841
transform 1 0 316 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1712256841
transform 1 0 236 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3758
timestamp 1712256841
transform 1 0 1188 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3759
timestamp 1712256841
transform 1 0 1100 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3760
timestamp 1712256841
transform 1 0 1372 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3761
timestamp 1712256841
transform 1 0 1340 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3762
timestamp 1712256841
transform 1 0 3132 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3763
timestamp 1712256841
transform 1 0 3044 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3764
timestamp 1712256841
transform 1 0 2988 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3765
timestamp 1712256841
transform 1 0 1012 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3766
timestamp 1712256841
transform 1 0 764 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3767
timestamp 1712256841
transform 1 0 1356 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3768
timestamp 1712256841
transform 1 0 988 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3769
timestamp 1712256841
transform 1 0 1044 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3770
timestamp 1712256841
transform 1 0 996 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3771
timestamp 1712256841
transform 1 0 1012 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3772
timestamp 1712256841
transform 1 0 940 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3773
timestamp 1712256841
transform 1 0 1380 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3774
timestamp 1712256841
transform 1 0 1348 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3775
timestamp 1712256841
transform 1 0 1340 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3776
timestamp 1712256841
transform 1 0 1308 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3777
timestamp 1712256841
transform 1 0 1308 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3778
timestamp 1712256841
transform 1 0 1140 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3779
timestamp 1712256841
transform 1 0 1060 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1712256841
transform 1 0 892 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3781
timestamp 1712256841
transform 1 0 1356 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3782
timestamp 1712256841
transform 1 0 1356 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3783
timestamp 1712256841
transform 1 0 1292 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1712256841
transform 1 0 1188 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3785
timestamp 1712256841
transform 1 0 1212 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3786
timestamp 1712256841
transform 1 0 1148 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3787
timestamp 1712256841
transform 1 0 2884 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3788
timestamp 1712256841
transform 1 0 2724 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3789
timestamp 1712256841
transform 1 0 2228 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3790
timestamp 1712256841
transform 1 0 1468 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3791
timestamp 1712256841
transform 1 0 1380 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3792
timestamp 1712256841
transform 1 0 1380 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3793
timestamp 1712256841
transform 1 0 1380 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1712256841
transform 1 0 1372 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3795
timestamp 1712256841
transform 1 0 1348 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3796
timestamp 1712256841
transform 1 0 1332 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1712256841
transform 1 0 1316 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1712256841
transform 1 0 1316 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3799
timestamp 1712256841
transform 1 0 1316 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1712256841
transform 1 0 1268 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1712256841
transform 1 0 1268 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3802
timestamp 1712256841
transform 1 0 2820 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3803
timestamp 1712256841
transform 1 0 1716 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3804
timestamp 1712256841
transform 1 0 1716 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3805
timestamp 1712256841
transform 1 0 1348 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3806
timestamp 1712256841
transform 1 0 1348 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3807
timestamp 1712256841
transform 1 0 1332 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3808
timestamp 1712256841
transform 1 0 1260 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3809
timestamp 1712256841
transform 1 0 1260 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3810
timestamp 1712256841
transform 1 0 1356 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3811
timestamp 1712256841
transform 1 0 1316 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3812
timestamp 1712256841
transform 1 0 1476 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1712256841
transform 1 0 1316 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1712256841
transform 1 0 1412 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1712256841
transform 1 0 1332 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3816
timestamp 1712256841
transform 1 0 1300 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3817
timestamp 1712256841
transform 1 0 1132 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3818
timestamp 1712256841
transform 1 0 1132 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3819
timestamp 1712256841
transform 1 0 1044 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3820
timestamp 1712256841
transform 1 0 1036 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3821
timestamp 1712256841
transform 1 0 1004 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1712256841
transform 1 0 956 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1712256841
transform 1 0 1572 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3824
timestamp 1712256841
transform 1 0 1484 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1712256841
transform 1 0 564 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1712256841
transform 1 0 524 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1712256841
transform 1 0 764 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1712256841
transform 1 0 540 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1712256841
transform 1 0 956 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1712256841
transform 1 0 812 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3831
timestamp 1712256841
transform 1 0 804 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1712256841
transform 1 0 740 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3833
timestamp 1712256841
transform 1 0 1140 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1712256841
transform 1 0 1100 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3835
timestamp 1712256841
transform 1 0 924 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3836
timestamp 1712256841
transform 1 0 836 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1712256841
transform 1 0 820 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1712256841
transform 1 0 812 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1712256841
transform 1 0 780 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1712256841
transform 1 0 316 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3841
timestamp 1712256841
transform 1 0 316 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3842
timestamp 1712256841
transform 1 0 284 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1712256841
transform 1 0 908 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3844
timestamp 1712256841
transform 1 0 804 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3845
timestamp 1712256841
transform 1 0 1228 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3846
timestamp 1712256841
transform 1 0 1084 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1712256841
transform 1 0 1140 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1712256841
transform 1 0 1100 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3849
timestamp 1712256841
transform 1 0 1596 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1712256841
transform 1 0 1572 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1712256841
transform 1 0 1516 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3852
timestamp 1712256841
transform 1 0 1516 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3853
timestamp 1712256841
transform 1 0 1340 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3854
timestamp 1712256841
transform 1 0 1316 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3855
timestamp 1712256841
transform 1 0 1276 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1712256841
transform 1 0 1276 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3857
timestamp 1712256841
transform 1 0 1204 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3858
timestamp 1712256841
transform 1 0 868 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3859
timestamp 1712256841
transform 1 0 1212 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3860
timestamp 1712256841
transform 1 0 1188 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3861
timestamp 1712256841
transform 1 0 2772 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3862
timestamp 1712256841
transform 1 0 2772 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3863
timestamp 1712256841
transform 1 0 2756 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3864
timestamp 1712256841
transform 1 0 2748 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3865
timestamp 1712256841
transform 1 0 2580 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3866
timestamp 1712256841
transform 1 0 1636 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3867
timestamp 1712256841
transform 1 0 1628 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3868
timestamp 1712256841
transform 1 0 1612 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3869
timestamp 1712256841
transform 1 0 1292 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3870
timestamp 1712256841
transform 1 0 1172 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3871
timestamp 1712256841
transform 1 0 1172 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3872
timestamp 1712256841
transform 1 0 1044 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3873
timestamp 1712256841
transform 1 0 596 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3874
timestamp 1712256841
transform 1 0 516 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3875
timestamp 1712256841
transform 1 0 2932 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3876
timestamp 1712256841
transform 1 0 2492 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3877
timestamp 1712256841
transform 1 0 2492 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3878
timestamp 1712256841
transform 1 0 1172 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3879
timestamp 1712256841
transform 1 0 1076 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3880
timestamp 1712256841
transform 1 0 1076 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3881
timestamp 1712256841
transform 1 0 1068 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3882
timestamp 1712256841
transform 1 0 1044 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3883
timestamp 1712256841
transform 1 0 1028 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3884
timestamp 1712256841
transform 1 0 884 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1712256841
transform 1 0 772 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3886
timestamp 1712256841
transform 1 0 1124 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3887
timestamp 1712256841
transform 1 0 844 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1712256841
transform 1 0 1556 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1712256841
transform 1 0 1548 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1712256841
transform 1 0 1308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3891
timestamp 1712256841
transform 1 0 1300 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3892
timestamp 1712256841
transform 1 0 1236 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3893
timestamp 1712256841
transform 1 0 1236 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3894
timestamp 1712256841
transform 1 0 1100 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3895
timestamp 1712256841
transform 1 0 948 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3896
timestamp 1712256841
transform 1 0 1212 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3897
timestamp 1712256841
transform 1 0 1108 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3898
timestamp 1712256841
transform 1 0 572 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1712256841
transform 1 0 444 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3900
timestamp 1712256841
transform 1 0 1276 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3901
timestamp 1712256841
transform 1 0 628 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1712256841
transform 1 0 628 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3903
timestamp 1712256841
transform 1 0 628 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3904
timestamp 1712256841
transform 1 0 572 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3905
timestamp 1712256841
transform 1 0 500 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3906
timestamp 1712256841
transform 1 0 476 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3907
timestamp 1712256841
transform 1 0 436 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3908
timestamp 1712256841
transform 1 0 348 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1712256841
transform 1 0 332 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3910
timestamp 1712256841
transform 1 0 324 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3911
timestamp 1712256841
transform 1 0 300 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3912
timestamp 1712256841
transform 1 0 716 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3913
timestamp 1712256841
transform 1 0 548 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3914
timestamp 1712256841
transform 1 0 676 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3915
timestamp 1712256841
transform 1 0 540 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3916
timestamp 1712256841
transform 1 0 532 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3917
timestamp 1712256841
transform 1 0 460 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1712256841
transform 1 0 340 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1712256841
transform 1 0 796 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3920
timestamp 1712256841
transform 1 0 628 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3921
timestamp 1712256841
transform 1 0 676 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3922
timestamp 1712256841
transform 1 0 644 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3923
timestamp 1712256841
transform 1 0 308 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1712256841
transform 1 0 308 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3925
timestamp 1712256841
transform 1 0 204 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3926
timestamp 1712256841
transform 1 0 1884 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1712256841
transform 1 0 1268 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1712256841
transform 1 0 1268 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1712256841
transform 1 0 1212 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3930
timestamp 1712256841
transform 1 0 1204 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3931
timestamp 1712256841
transform 1 0 780 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1712256841
transform 1 0 2836 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1712256841
transform 1 0 2772 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3934
timestamp 1712256841
transform 1 0 2772 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3935
timestamp 1712256841
transform 1 0 1852 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3936
timestamp 1712256841
transform 1 0 1852 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3937
timestamp 1712256841
transform 1 0 1780 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1712256841
transform 1 0 1468 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1712256841
transform 1 0 964 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1712256841
transform 1 0 932 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3941
timestamp 1712256841
transform 1 0 2844 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1712256841
transform 1 0 2460 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1712256841
transform 1 0 2460 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1712256841
transform 1 0 2316 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1712256841
transform 1 0 2316 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1712256841
transform 1 0 1444 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1712256841
transform 1 0 1436 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3948
timestamp 1712256841
transform 1 0 1276 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3949
timestamp 1712256841
transform 1 0 1028 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1712256841
transform 1 0 1028 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1712256841
transform 1 0 996 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1712256841
transform 1 0 996 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3953
timestamp 1712256841
transform 1 0 908 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1712256841
transform 1 0 908 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3955
timestamp 1712256841
transform 1 0 820 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3956
timestamp 1712256841
transform 1 0 820 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3957
timestamp 1712256841
transform 1 0 708 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1712256841
transform 1 0 684 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3959
timestamp 1712256841
transform 1 0 1972 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3960
timestamp 1712256841
transform 1 0 1364 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1712256841
transform 1 0 660 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3962
timestamp 1712256841
transform 1 0 660 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1712256841
transform 1 0 660 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1712256841
transform 1 0 628 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3965
timestamp 1712256841
transform 1 0 596 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3966
timestamp 1712256841
transform 1 0 1052 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3967
timestamp 1712256841
transform 1 0 940 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3968
timestamp 1712256841
transform 1 0 868 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3969
timestamp 1712256841
transform 1 0 868 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3970
timestamp 1712256841
transform 1 0 868 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3971
timestamp 1712256841
transform 1 0 764 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3972
timestamp 1712256841
transform 1 0 732 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3973
timestamp 1712256841
transform 1 0 2764 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3974
timestamp 1712256841
transform 1 0 1364 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3975
timestamp 1712256841
transform 1 0 1364 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_3976
timestamp 1712256841
transform 1 0 1300 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3977
timestamp 1712256841
transform 1 0 1268 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3978
timestamp 1712256841
transform 1 0 1268 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3979
timestamp 1712256841
transform 1 0 1268 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3980
timestamp 1712256841
transform 1 0 1236 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3981
timestamp 1712256841
transform 1 0 1220 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3982
timestamp 1712256841
transform 1 0 1212 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3983
timestamp 1712256841
transform 1 0 1204 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3984
timestamp 1712256841
transform 1 0 1196 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3985
timestamp 1712256841
transform 1 0 1116 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3986
timestamp 1712256841
transform 1 0 1108 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3987
timestamp 1712256841
transform 1 0 1028 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3988
timestamp 1712256841
transform 1 0 1028 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3989
timestamp 1712256841
transform 1 0 364 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3990
timestamp 1712256841
transform 1 0 292 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3991
timestamp 1712256841
transform 1 0 268 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1712256841
transform 1 0 236 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3993
timestamp 1712256841
transform 1 0 564 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1712256841
transform 1 0 308 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3995
timestamp 1712256841
transform 1 0 364 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3996
timestamp 1712256841
transform 1 0 332 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3997
timestamp 1712256841
transform 1 0 740 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3998
timestamp 1712256841
transform 1 0 340 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3999
timestamp 1712256841
transform 1 0 828 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4000
timestamp 1712256841
transform 1 0 300 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4001
timestamp 1712256841
transform 1 0 252 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4002
timestamp 1712256841
transform 1 0 220 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4003
timestamp 1712256841
transform 1 0 212 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4004
timestamp 1712256841
transform 1 0 148 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4005
timestamp 1712256841
transform 1 0 996 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4006
timestamp 1712256841
transform 1 0 596 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4007
timestamp 1712256841
transform 1 0 572 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4008
timestamp 1712256841
transform 1 0 180 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4009
timestamp 1712256841
transform 1 0 132 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4010
timestamp 1712256841
transform 1 0 108 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4011
timestamp 1712256841
transform 1 0 1932 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4012
timestamp 1712256841
transform 1 0 1876 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4013
timestamp 1712256841
transform 1 0 1876 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4014
timestamp 1712256841
transform 1 0 1492 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1712256841
transform 1 0 1492 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4016
timestamp 1712256841
transform 1 0 972 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4017
timestamp 1712256841
transform 1 0 956 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4018
timestamp 1712256841
transform 1 0 956 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1712256841
transform 1 0 148 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4020
timestamp 1712256841
transform 1 0 108 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4021
timestamp 1712256841
transform 1 0 2772 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4022
timestamp 1712256841
transform 1 0 2388 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4023
timestamp 1712256841
transform 1 0 2388 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4024
timestamp 1712256841
transform 1 0 2340 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1712256841
transform 1 0 1564 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4026
timestamp 1712256841
transform 1 0 1516 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4027
timestamp 1712256841
transform 1 0 1516 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4028
timestamp 1712256841
transform 1 0 892 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4029
timestamp 1712256841
transform 1 0 796 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4030
timestamp 1712256841
transform 1 0 796 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4031
timestamp 1712256841
transform 1 0 788 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4032
timestamp 1712256841
transform 1 0 708 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4033
timestamp 1712256841
transform 1 0 2028 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4034
timestamp 1712256841
transform 1 0 1732 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4035
timestamp 1712256841
transform 1 0 1684 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4036
timestamp 1712256841
transform 1 0 1684 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4037
timestamp 1712256841
transform 1 0 836 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4038
timestamp 1712256841
transform 1 0 1124 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1712256841
transform 1 0 1060 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4040
timestamp 1712256841
transform 1 0 1060 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1712256841
transform 1 0 964 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4042
timestamp 1712256841
transform 1 0 900 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4043
timestamp 1712256841
transform 1 0 900 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4044
timestamp 1712256841
transform 1 0 628 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4045
timestamp 1712256841
transform 1 0 428 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4046
timestamp 1712256841
transform 1 0 228 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4047
timestamp 1712256841
transform 1 0 564 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4048
timestamp 1712256841
transform 1 0 388 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4049
timestamp 1712256841
transform 1 0 1076 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4050
timestamp 1712256841
transform 1 0 812 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4051
timestamp 1712256841
transform 1 0 612 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4052
timestamp 1712256841
transform 1 0 612 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4053
timestamp 1712256841
transform 1 0 540 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4054
timestamp 1712256841
transform 1 0 532 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4055
timestamp 1712256841
transform 1 0 532 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4056
timestamp 1712256841
transform 1 0 516 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4057
timestamp 1712256841
transform 1 0 516 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4058
timestamp 1712256841
transform 1 0 372 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4059
timestamp 1712256841
transform 1 0 340 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4060
timestamp 1712256841
transform 1 0 316 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4061
timestamp 1712256841
transform 1 0 292 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4062
timestamp 1712256841
transform 1 0 292 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4063
timestamp 1712256841
transform 1 0 260 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4064
timestamp 1712256841
transform 1 0 252 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4065
timestamp 1712256841
transform 1 0 948 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4066
timestamp 1712256841
transform 1 0 348 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4067
timestamp 1712256841
transform 1 0 1092 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4068
timestamp 1712256841
transform 1 0 388 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4069
timestamp 1712256841
transform 1 0 340 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4070
timestamp 1712256841
transform 1 0 268 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4071
timestamp 1712256841
transform 1 0 196 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4072
timestamp 1712256841
transform 1 0 188 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4073
timestamp 1712256841
transform 1 0 988 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4074
timestamp 1712256841
transform 1 0 500 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1712256841
transform 1 0 516 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4076
timestamp 1712256841
transform 1 0 492 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4077
timestamp 1712256841
transform 1 0 164 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4078
timestamp 1712256841
transform 1 0 196 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4079
timestamp 1712256841
transform 1 0 116 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4080
timestamp 1712256841
transform 1 0 1188 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4081
timestamp 1712256841
transform 1 0 924 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4082
timestamp 1712256841
transform 1 0 1268 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4083
timestamp 1712256841
transform 1 0 1196 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4084
timestamp 1712256841
transform 1 0 1116 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4085
timestamp 1712256841
transform 1 0 1116 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4086
timestamp 1712256841
transform 1 0 1116 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4087
timestamp 1712256841
transform 1 0 1116 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1712256841
transform 1 0 1092 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4089
timestamp 1712256841
transform 1 0 1012 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4090
timestamp 1712256841
transform 1 0 1012 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4091
timestamp 1712256841
transform 1 0 900 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4092
timestamp 1712256841
transform 1 0 788 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4093
timestamp 1712256841
transform 1 0 1212 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4094
timestamp 1712256841
transform 1 0 1068 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1712256841
transform 1 0 1172 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4096
timestamp 1712256841
transform 1 0 1076 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4097
timestamp 1712256841
transform 1 0 1124 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4098
timestamp 1712256841
transform 1 0 940 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1712256841
transform 1 0 940 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4100
timestamp 1712256841
transform 1 0 932 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1712256841
transform 1 0 916 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4102
timestamp 1712256841
transform 1 0 884 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4103
timestamp 1712256841
transform 1 0 676 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1712256841
transform 1 0 1108 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4105
timestamp 1712256841
transform 1 0 1084 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4106
timestamp 1712256841
transform 1 0 1740 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4107
timestamp 1712256841
transform 1 0 1340 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4108
timestamp 1712256841
transform 1 0 1156 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4109
timestamp 1712256841
transform 1 0 356 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4110
timestamp 1712256841
transform 1 0 220 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4111
timestamp 1712256841
transform 1 0 564 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1712256841
transform 1 0 388 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4113
timestamp 1712256841
transform 1 0 732 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4114
timestamp 1712256841
transform 1 0 500 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1712256841
transform 1 0 460 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4116
timestamp 1712256841
transform 1 0 452 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4117
timestamp 1712256841
transform 1 0 1220 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4118
timestamp 1712256841
transform 1 0 708 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4119
timestamp 1712256841
transform 1 0 652 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1712256841
transform 1 0 476 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4121
timestamp 1712256841
transform 1 0 436 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4122
timestamp 1712256841
transform 1 0 420 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4123
timestamp 1712256841
transform 1 0 420 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4124
timestamp 1712256841
transform 1 0 420 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4125
timestamp 1712256841
transform 1 0 324 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4126
timestamp 1712256841
transform 1 0 276 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4127
timestamp 1712256841
transform 1 0 276 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4128
timestamp 1712256841
transform 1 0 228 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4129
timestamp 1712256841
transform 1 0 212 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4130
timestamp 1712256841
transform 1 0 204 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4131
timestamp 1712256841
transform 1 0 740 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4132
timestamp 1712256841
transform 1 0 644 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4133
timestamp 1712256841
transform 1 0 860 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4134
timestamp 1712256841
transform 1 0 796 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4135
timestamp 1712256841
transform 1 0 756 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4136
timestamp 1712256841
transform 1 0 708 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4137
timestamp 1712256841
transform 1 0 204 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4138
timestamp 1712256841
transform 1 0 100 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4139
timestamp 1712256841
transform 1 0 276 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4140
timestamp 1712256841
transform 1 0 252 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4141
timestamp 1712256841
transform 1 0 772 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4142
timestamp 1712256841
transform 1 0 740 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1712256841
transform 1 0 844 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1712256841
transform 1 0 324 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4145
timestamp 1712256841
transform 1 0 940 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1712256841
transform 1 0 812 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4147
timestamp 1712256841
transform 1 0 1004 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4148
timestamp 1712256841
transform 1 0 1004 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4149
timestamp 1712256841
transform 1 0 908 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4150
timestamp 1712256841
transform 1 0 852 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4151
timestamp 1712256841
transform 1 0 652 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4152
timestamp 1712256841
transform 1 0 988 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1712256841
transform 1 0 964 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4154
timestamp 1712256841
transform 1 0 2764 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4155
timestamp 1712256841
transform 1 0 2764 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4156
timestamp 1712256841
transform 1 0 2740 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4157
timestamp 1712256841
transform 1 0 2740 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1712256841
transform 1 0 1884 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4159
timestamp 1712256841
transform 1 0 1844 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4160
timestamp 1712256841
transform 1 0 1588 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4161
timestamp 1712256841
transform 1 0 1372 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4162
timestamp 1712256841
transform 1 0 1372 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4163
timestamp 1712256841
transform 1 0 1372 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4164
timestamp 1712256841
transform 1 0 1308 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4165
timestamp 1712256841
transform 1 0 1292 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4166
timestamp 1712256841
transform 1 0 156 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1712256841
transform 1 0 124 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4168
timestamp 1712256841
transform 1 0 108 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4169
timestamp 1712256841
transform 1 0 108 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4170
timestamp 1712256841
transform 1 0 132 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4171
timestamp 1712256841
transform 1 0 84 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4172
timestamp 1712256841
transform 1 0 420 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4173
timestamp 1712256841
transform 1 0 108 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4174
timestamp 1712256841
transform 1 0 516 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4175
timestamp 1712256841
transform 1 0 444 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4176
timestamp 1712256841
transform 1 0 668 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4177
timestamp 1712256841
transform 1 0 580 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4178
timestamp 1712256841
transform 1 0 724 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4179
timestamp 1712256841
transform 1 0 668 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4180
timestamp 1712256841
transform 1 0 596 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4181
timestamp 1712256841
transform 1 0 132 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4182
timestamp 1712256841
transform 1 0 108 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4183
timestamp 1712256841
transform 1 0 612 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1712256841
transform 1 0 468 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4185
timestamp 1712256841
transform 1 0 708 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4186
timestamp 1712256841
transform 1 0 644 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4187
timestamp 1712256841
transform 1 0 772 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4188
timestamp 1712256841
transform 1 0 164 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1712256841
transform 1 0 860 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4190
timestamp 1712256841
transform 1 0 756 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4191
timestamp 1712256841
transform 1 0 852 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4192
timestamp 1712256841
transform 1 0 796 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4193
timestamp 1712256841
transform 1 0 884 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4194
timestamp 1712256841
transform 1 0 860 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4195
timestamp 1712256841
transform 1 0 932 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1712256841
transform 1 0 796 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4197
timestamp 1712256841
transform 1 0 740 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4198
timestamp 1712256841
transform 1 0 988 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4199
timestamp 1712256841
transform 1 0 868 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4200
timestamp 1712256841
transform 1 0 172 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1712256841
transform 1 0 116 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1712256841
transform 1 0 68 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4203
timestamp 1712256841
transform 1 0 68 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4204
timestamp 1712256841
transform 1 0 380 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4205
timestamp 1712256841
transform 1 0 84 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4206
timestamp 1712256841
transform 1 0 516 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4207
timestamp 1712256841
transform 1 0 404 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4208
timestamp 1712256841
transform 1 0 668 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4209
timestamp 1712256841
transform 1 0 452 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1712256841
transform 1 0 1060 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1712256841
transform 1 0 1044 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4212
timestamp 1712256841
transform 1 0 988 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4213
timestamp 1712256841
transform 1 0 884 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1712256841
transform 1 0 836 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1712256841
transform 1 0 836 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4216
timestamp 1712256841
transform 1 0 580 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4217
timestamp 1712256841
transform 1 0 580 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4218
timestamp 1712256841
transform 1 0 276 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4219
timestamp 1712256841
transform 1 0 228 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4220
timestamp 1712256841
transform 1 0 692 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4221
timestamp 1712256841
transform 1 0 564 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4222
timestamp 1712256841
transform 1 0 732 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4223
timestamp 1712256841
transform 1 0 628 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4224
timestamp 1712256841
transform 1 0 108 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1712256841
transform 1 0 84 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4226
timestamp 1712256841
transform 1 0 164 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4227
timestamp 1712256841
transform 1 0 140 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4228
timestamp 1712256841
transform 1 0 724 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4229
timestamp 1712256841
transform 1 0 692 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4230
timestamp 1712256841
transform 1 0 796 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4231
timestamp 1712256841
transform 1 0 212 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1712256841
transform 1 0 844 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4233
timestamp 1712256841
transform 1 0 756 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4234
timestamp 1712256841
transform 1 0 860 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4235
timestamp 1712256841
transform 1 0 820 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4236
timestamp 1712256841
transform 1 0 868 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4237
timestamp 1712256841
transform 1 0 836 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1712256841
transform 1 0 1308 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4239
timestamp 1712256841
transform 1 0 1124 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1712256841
transform 1 0 1060 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4241
timestamp 1712256841
transform 1 0 972 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4242
timestamp 1712256841
transform 1 0 900 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4243
timestamp 1712256841
transform 1 0 860 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4244
timestamp 1712256841
transform 1 0 972 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4245
timestamp 1712256841
transform 1 0 836 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4246
timestamp 1712256841
transform 1 0 2956 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4247
timestamp 1712256841
transform 1 0 2924 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4248
timestamp 1712256841
transform 1 0 2916 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4249
timestamp 1712256841
transform 1 0 2572 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4250
timestamp 1712256841
transform 1 0 2572 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4251
timestamp 1712256841
transform 1 0 2412 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4252
timestamp 1712256841
transform 1 0 2396 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4253
timestamp 1712256841
transform 1 0 2284 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1712256841
transform 1 0 2284 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4255
timestamp 1712256841
transform 1 0 1348 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4256
timestamp 1712256841
transform 1 0 1348 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4257
timestamp 1712256841
transform 1 0 1276 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4258
timestamp 1712256841
transform 1 0 1236 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4259
timestamp 1712256841
transform 1 0 1220 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1712256841
transform 1 0 1068 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4261
timestamp 1712256841
transform 1 0 644 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4262
timestamp 1712256841
transform 1 0 372 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4263
timestamp 1712256841
transform 1 0 364 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4264
timestamp 1712256841
transform 1 0 284 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4265
timestamp 1712256841
transform 1 0 228 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4266
timestamp 1712256841
transform 1 0 132 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4267
timestamp 1712256841
transform 1 0 340 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4268
timestamp 1712256841
transform 1 0 236 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4269
timestamp 1712256841
transform 1 0 620 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4270
timestamp 1712256841
transform 1 0 316 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4271
timestamp 1712256841
transform 1 0 420 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4272
timestamp 1712256841
transform 1 0 380 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4273
timestamp 1712256841
transform 1 0 1284 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4274
timestamp 1712256841
transform 1 0 1132 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4275
timestamp 1712256841
transform 1 0 1132 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1712256841
transform 1 0 1060 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4277
timestamp 1712256841
transform 1 0 676 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4278
timestamp 1712256841
transform 1 0 668 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1712256841
transform 1 0 468 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4280
timestamp 1712256841
transform 1 0 444 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4281
timestamp 1712256841
transform 1 0 412 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4282
timestamp 1712256841
transform 1 0 284 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4283
timestamp 1712256841
transform 1 0 588 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4284
timestamp 1712256841
transform 1 0 460 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4285
timestamp 1712256841
transform 1 0 316 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4286
timestamp 1712256841
transform 1 0 964 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4287
timestamp 1712256841
transform 1 0 820 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4288
timestamp 1712256841
transform 1 0 812 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4289
timestamp 1712256841
transform 1 0 524 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4290
timestamp 1712256841
transform 1 0 524 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4291
timestamp 1712256841
transform 1 0 252 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4292
timestamp 1712256841
transform 1 0 180 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4293
timestamp 1712256841
transform 1 0 932 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4294
timestamp 1712256841
transform 1 0 676 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4295
timestamp 1712256841
transform 1 0 220 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4296
timestamp 1712256841
transform 1 0 140 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4297
timestamp 1712256841
transform 1 0 1148 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1712256841
transform 1 0 628 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4299
timestamp 1712256841
transform 1 0 1388 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4300
timestamp 1712256841
transform 1 0 1172 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1712256841
transform 1 0 1068 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4302
timestamp 1712256841
transform 1 0 1036 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4303
timestamp 1712256841
transform 1 0 1276 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4304
timestamp 1712256841
transform 1 0 940 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4305
timestamp 1712256841
transform 1 0 996 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1712256841
transform 1 0 948 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4307
timestamp 1712256841
transform 1 0 1060 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4308
timestamp 1712256841
transform 1 0 980 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4309
timestamp 1712256841
transform 1 0 1684 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4310
timestamp 1712256841
transform 1 0 1588 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4311
timestamp 1712256841
transform 1 0 1380 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4312
timestamp 1712256841
transform 1 0 1020 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4313
timestamp 1712256841
transform 1 0 2956 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4314
timestamp 1712256841
transform 1 0 2476 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4315
timestamp 1712256841
transform 1 0 2476 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4316
timestamp 1712256841
transform 1 0 1772 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4317
timestamp 1712256841
transform 1 0 1764 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4318
timestamp 1712256841
transform 1 0 1404 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4319
timestamp 1712256841
transform 1 0 1388 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4320
timestamp 1712256841
transform 1 0 1148 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4321
timestamp 1712256841
transform 1 0 1076 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4322
timestamp 1712256841
transform 1 0 2708 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1712256841
transform 1 0 2540 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4324
timestamp 1712256841
transform 1 0 1748 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4325
timestamp 1712256841
transform 1 0 1500 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4326
timestamp 1712256841
transform 1 0 1348 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4327
timestamp 1712256841
transform 1 0 1036 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4328
timestamp 1712256841
transform 1 0 396 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4329
timestamp 1712256841
transform 1 0 396 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1712256841
transform 1 0 396 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4331
timestamp 1712256841
transform 1 0 388 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4332
timestamp 1712256841
transform 1 0 356 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1712256841
transform 1 0 356 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4334
timestamp 1712256841
transform 1 0 244 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4335
timestamp 1712256841
transform 1 0 172 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4336
timestamp 1712256841
transform 1 0 172 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4337
timestamp 1712256841
transform 1 0 788 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_4338
timestamp 1712256841
transform 1 0 260 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_4339
timestamp 1712256841
transform 1 0 412 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4340
timestamp 1712256841
transform 1 0 324 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4341
timestamp 1712256841
transform 1 0 788 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1712256841
transform 1 0 396 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4343
timestamp 1712256841
transform 1 0 300 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1712256841
transform 1 0 1028 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_4345
timestamp 1712256841
transform 1 0 580 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_4346
timestamp 1712256841
transform 1 0 284 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4347
timestamp 1712256841
transform 1 0 284 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4348
timestamp 1712256841
transform 1 0 236 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_4349
timestamp 1712256841
transform 1 0 156 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4350
timestamp 1712256841
transform 1 0 1060 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4351
timestamp 1712256841
transform 1 0 1012 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4352
timestamp 1712256841
transform 1 0 804 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4353
timestamp 1712256841
transform 1 0 908 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4354
timestamp 1712256841
transform 1 0 756 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4355
timestamp 1712256841
transform 1 0 900 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4356
timestamp 1712256841
transform 1 0 860 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4357
timestamp 1712256841
transform 1 0 1204 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4358
timestamp 1712256841
transform 1 0 988 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4359
timestamp 1712256841
transform 1 0 1188 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4360
timestamp 1712256841
transform 1 0 1164 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4361
timestamp 1712256841
transform 1 0 2908 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4362
timestamp 1712256841
transform 1 0 2844 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4363
timestamp 1712256841
transform 1 0 2508 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4364
timestamp 1712256841
transform 1 0 2508 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4365
timestamp 1712256841
transform 1 0 1844 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4366
timestamp 1712256841
transform 1 0 1804 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4367
timestamp 1712256841
transform 1 0 1572 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4368
timestamp 1712256841
transform 1 0 1412 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4369
timestamp 1712256841
transform 1 0 1092 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4370
timestamp 1712256841
transform 1 0 1148 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4371
timestamp 1712256841
transform 1 0 644 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1712256841
transform 1 0 76 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4373
timestamp 1712256841
transform 1 0 76 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4374
timestamp 1712256841
transform 1 0 620 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4375
timestamp 1712256841
transform 1 0 412 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4376
timestamp 1712256841
transform 1 0 612 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4377
timestamp 1712256841
transform 1 0 500 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4378
timestamp 1712256841
transform 1 0 692 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4379
timestamp 1712256841
transform 1 0 660 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4380
timestamp 1712256841
transform 1 0 660 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_4381
timestamp 1712256841
transform 1 0 564 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_4382
timestamp 1712256841
transform 1 0 636 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4383
timestamp 1712256841
transform 1 0 588 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4384
timestamp 1712256841
transform 1 0 588 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4385
timestamp 1712256841
transform 1 0 532 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4386
timestamp 1712256841
transform 1 0 380 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4387
timestamp 1712256841
transform 1 0 1204 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4388
timestamp 1712256841
transform 1 0 732 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1712256841
transform 1 0 692 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4390
timestamp 1712256841
transform 1 0 644 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4391
timestamp 1712256841
transform 1 0 812 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4392
timestamp 1712256841
transform 1 0 692 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4393
timestamp 1712256841
transform 1 0 796 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4394
timestamp 1712256841
transform 1 0 756 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4395
timestamp 1712256841
transform 1 0 516 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4396
timestamp 1712256841
transform 1 0 404 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_4397
timestamp 1712256841
transform 1 0 420 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_4398
timestamp 1712256841
transform 1 0 340 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_4399
timestamp 1712256841
transform 1 0 1588 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4400
timestamp 1712256841
transform 1 0 1548 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1712256841
transform 1 0 1484 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4402
timestamp 1712256841
transform 1 0 1484 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4403
timestamp 1712256841
transform 1 0 1268 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4404
timestamp 1712256841
transform 1 0 1268 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4405
timestamp 1712256841
transform 1 0 1172 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4406
timestamp 1712256841
transform 1 0 2748 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4407
timestamp 1712256841
transform 1 0 2460 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4408
timestamp 1712256841
transform 1 0 2460 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1712256841
transform 1 0 1268 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4410
timestamp 1712256841
transform 1 0 1244 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4411
timestamp 1712256841
transform 1 0 1204 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4412
timestamp 1712256841
transform 1 0 1204 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4413
timestamp 1712256841
transform 1 0 1068 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4414
timestamp 1712256841
transform 1 0 1060 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4415
timestamp 1712256841
transform 1 0 1004 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4416
timestamp 1712256841
transform 1 0 1388 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1712256841
transform 1 0 892 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4418
timestamp 1712256841
transform 1 0 876 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1712256841
transform 1 0 876 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4420
timestamp 1712256841
transform 1 0 900 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4421
timestamp 1712256841
transform 1 0 868 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1712256841
transform 1 0 940 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4423
timestamp 1712256841
transform 1 0 908 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4424
timestamp 1712256841
transform 1 0 2444 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4425
timestamp 1712256841
transform 1 0 2412 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4426
timestamp 1712256841
transform 1 0 2260 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1712256841
transform 1 0 1476 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4428
timestamp 1712256841
transform 1 0 1476 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4429
timestamp 1712256841
transform 1 0 956 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4430
timestamp 1712256841
transform 1 0 956 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1712256841
transform 1 0 916 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4432
timestamp 1712256841
transform 1 0 876 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4433
timestamp 1712256841
transform 1 0 812 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4434
timestamp 1712256841
transform 1 0 948 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4435
timestamp 1712256841
transform 1 0 932 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4436
timestamp 1712256841
transform 1 0 836 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_4437
timestamp 1712256841
transform 1 0 1252 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4438
timestamp 1712256841
transform 1 0 1132 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4439
timestamp 1712256841
transform 1 0 1132 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4440
timestamp 1712256841
transform 1 0 940 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4441
timestamp 1712256841
transform 1 0 908 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4442
timestamp 1712256841
transform 1 0 1796 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4443
timestamp 1712256841
transform 1 0 1740 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4444
timestamp 1712256841
transform 1 0 1740 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4445
timestamp 1712256841
transform 1 0 1620 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1712256841
transform 1 0 1332 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1712256841
transform 1 0 1316 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4448
timestamp 1712256841
transform 1 0 1228 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4449
timestamp 1712256841
transform 1 0 1444 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4450
timestamp 1712256841
transform 1 0 1228 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4451
timestamp 1712256841
transform 1 0 1180 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4452
timestamp 1712256841
transform 1 0 1180 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4453
timestamp 1712256841
transform 1 0 1180 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4454
timestamp 1712256841
transform 1 0 1180 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4455
timestamp 1712256841
transform 1 0 1140 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4456
timestamp 1712256841
transform 1 0 1132 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4457
timestamp 1712256841
transform 1 0 1140 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4458
timestamp 1712256841
transform 1 0 1076 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4459
timestamp 1712256841
transform 1 0 1212 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1712256841
transform 1 0 1140 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4461
timestamp 1712256841
transform 1 0 1092 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4462
timestamp 1712256841
transform 1 0 1092 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4463
timestamp 1712256841
transform 1 0 1052 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_4464
timestamp 1712256841
transform 1 0 1108 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1712256841
transform 1 0 1044 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1712256841
transform 1 0 1764 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4467
timestamp 1712256841
transform 1 0 1668 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4468
timestamp 1712256841
transform 1 0 1668 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4469
timestamp 1712256841
transform 1 0 1532 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4470
timestamp 1712256841
transform 1 0 1532 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4471
timestamp 1712256841
transform 1 0 1412 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4472
timestamp 1712256841
transform 1 0 1196 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1712256841
transform 1 0 1196 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4474
timestamp 1712256841
transform 1 0 1132 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4475
timestamp 1712256841
transform 1 0 2004 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4476
timestamp 1712256841
transform 1 0 1844 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4477
timestamp 1712256841
transform 1 0 1724 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4478
timestamp 1712256841
transform 1 0 1652 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4479
timestamp 1712256841
transform 1 0 1516 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4480
timestamp 1712256841
transform 1 0 1452 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4481
timestamp 1712256841
transform 1 0 1564 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1712256841
transform 1 0 1524 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4483
timestamp 1712256841
transform 1 0 1468 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4484
timestamp 1712256841
transform 1 0 1444 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4485
timestamp 1712256841
transform 1 0 1468 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1712256841
transform 1 0 1316 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4487
timestamp 1712256841
transform 1 0 1372 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4488
timestamp 1712256841
transform 1 0 1332 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4489
timestamp 1712256841
transform 1 0 1444 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4490
timestamp 1712256841
transform 1 0 1332 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4491
timestamp 1712256841
transform 1 0 1332 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4492
timestamp 1712256841
transform 1 0 1252 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4493
timestamp 1712256841
transform 1 0 1532 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4494
timestamp 1712256841
transform 1 0 1460 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_4495
timestamp 1712256841
transform 1 0 1372 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4496
timestamp 1712256841
transform 1 0 1356 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4497
timestamp 1712256841
transform 1 0 1500 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4498
timestamp 1712256841
transform 1 0 1412 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1712256841
transform 1 0 1620 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4500
timestamp 1712256841
transform 1 0 1532 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1712256841
transform 1 0 1908 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4502
timestamp 1712256841
transform 1 0 1884 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4503
timestamp 1712256841
transform 1 0 1820 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4504
timestamp 1712256841
transform 1 0 1700 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4505
timestamp 1712256841
transform 1 0 1708 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4506
timestamp 1712256841
transform 1 0 1652 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4507
timestamp 1712256841
transform 1 0 1612 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4508
timestamp 1712256841
transform 1 0 1772 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1712256841
transform 1 0 1716 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4510
timestamp 1712256841
transform 1 0 1900 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4511
timestamp 1712256841
transform 1 0 1852 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4512
timestamp 1712256841
transform 1 0 1780 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4513
timestamp 1712256841
transform 1 0 1700 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4514
timestamp 1712256841
transform 1 0 1372 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4515
timestamp 1712256841
transform 1 0 2060 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4516
timestamp 1712256841
transform 1 0 1876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4517
timestamp 1712256841
transform 1 0 1876 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4518
timestamp 1712256841
transform 1 0 1828 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4519
timestamp 1712256841
transform 1 0 1828 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4520
timestamp 1712256841
transform 1 0 1828 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_4521
timestamp 1712256841
transform 1 0 1708 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4522
timestamp 1712256841
transform 1 0 1700 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4523
timestamp 1712256841
transform 1 0 1660 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4524
timestamp 1712256841
transform 1 0 1652 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4525
timestamp 1712256841
transform 1 0 1588 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_4526
timestamp 1712256841
transform 1 0 1588 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4527
timestamp 1712256841
transform 1 0 1516 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4528
timestamp 1712256841
transform 1 0 1508 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4529
timestamp 1712256841
transform 1 0 2188 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4530
timestamp 1712256841
transform 1 0 2036 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_4531
timestamp 1712256841
transform 1 0 2044 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4532
timestamp 1712256841
transform 1 0 1852 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4533
timestamp 1712256841
transform 1 0 836 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1712256841
transform 1 0 836 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4535
timestamp 1712256841
transform 1 0 636 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4536
timestamp 1712256841
transform 1 0 2004 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4537
timestamp 1712256841
transform 1 0 1924 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4538
timestamp 1712256841
transform 1 0 1924 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4539
timestamp 1712256841
transform 1 0 1884 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4540
timestamp 1712256841
transform 1 0 2188 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4541
timestamp 1712256841
transform 1 0 1972 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4542
timestamp 1712256841
transform 1 0 1908 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4543
timestamp 1712256841
transform 1 0 1876 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4544
timestamp 1712256841
transform 1 0 1860 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4545
timestamp 1712256841
transform 1 0 1844 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4546
timestamp 1712256841
transform 1 0 1572 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4547
timestamp 1712256841
transform 1 0 3420 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4548
timestamp 1712256841
transform 1 0 3420 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4549
timestamp 1712256841
transform 1 0 2380 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4550
timestamp 1712256841
transform 1 0 1932 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4551
timestamp 1712256841
transform 1 0 2380 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4552
timestamp 1712256841
transform 1 0 2300 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4553
timestamp 1712256841
transform 1 0 2500 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4554
timestamp 1712256841
transform 1 0 2420 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4555
timestamp 1712256841
transform 1 0 2436 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4556
timestamp 1712256841
transform 1 0 2396 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4557
timestamp 1712256841
transform 1 0 2180 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4558
timestamp 1712256841
transform 1 0 2340 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4559
timestamp 1712256841
transform 1 0 2140 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4560
timestamp 1712256841
transform 1 0 2140 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4561
timestamp 1712256841
transform 1 0 2092 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4562
timestamp 1712256841
transform 1 0 2092 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4563
timestamp 1712256841
transform 1 0 1820 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4564
timestamp 1712256841
transform 1 0 2020 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4565
timestamp 1712256841
transform 1 0 1948 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4566
timestamp 1712256841
transform 1 0 1900 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4567
timestamp 1712256841
transform 1 0 1796 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4568
timestamp 1712256841
transform 1 0 2132 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4569
timestamp 1712256841
transform 1 0 2060 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4570
timestamp 1712256841
transform 1 0 2420 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1712256841
transform 1 0 2204 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1712256841
transform 1 0 2204 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4573
timestamp 1712256841
transform 1 0 2068 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4574
timestamp 1712256841
transform 1 0 2020 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4575
timestamp 1712256841
transform 1 0 2020 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4576
timestamp 1712256841
transform 1 0 1940 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4577
timestamp 1712256841
transform 1 0 1748 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4578
timestamp 1712256841
transform 1 0 1724 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4579
timestamp 1712256841
transform 1 0 1684 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4580
timestamp 1712256841
transform 1 0 1668 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4581
timestamp 1712256841
transform 1 0 1684 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4582
timestamp 1712256841
transform 1 0 1604 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4583
timestamp 1712256841
transform 1 0 1692 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4584
timestamp 1712256841
transform 1 0 1516 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4585
timestamp 1712256841
transform 1 0 1476 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4586
timestamp 1712256841
transform 1 0 2348 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4587
timestamp 1712256841
transform 1 0 2156 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4588
timestamp 1712256841
transform 1 0 2436 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4589
timestamp 1712256841
transform 1 0 2308 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4590
timestamp 1712256841
transform 1 0 2444 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4591
timestamp 1712256841
transform 1 0 2364 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4592
timestamp 1712256841
transform 1 0 2564 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4593
timestamp 1712256841
transform 1 0 2404 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4594
timestamp 1712256841
transform 1 0 2340 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4595
timestamp 1712256841
transform 1 0 2332 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4596
timestamp 1712256841
transform 1 0 2284 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4597
timestamp 1712256841
transform 1 0 2260 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4598
timestamp 1712256841
transform 1 0 2260 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4599
timestamp 1712256841
transform 1 0 2252 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4600
timestamp 1712256841
transform 1 0 2252 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1712256841
transform 1 0 2212 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1712256841
transform 1 0 2196 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1712256841
transform 1 0 2188 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4604
timestamp 1712256841
transform 1 0 2060 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1712256841
transform 1 0 2060 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1712256841
transform 1 0 2052 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4607
timestamp 1712256841
transform 1 0 1988 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4608
timestamp 1712256841
transform 1 0 2588 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1712256841
transform 1 0 2532 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4610
timestamp 1712256841
transform 1 0 2388 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4611
timestamp 1712256841
transform 1 0 2340 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4612
timestamp 1712256841
transform 1 0 2204 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4613
timestamp 1712256841
transform 1 0 2204 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1712256841
transform 1 0 2172 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4615
timestamp 1712256841
transform 1 0 1604 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4616
timestamp 1712256841
transform 1 0 2084 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1712256841
transform 1 0 1660 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4618
timestamp 1712256841
transform 1 0 2284 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4619
timestamp 1712256841
transform 1 0 2236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1712256841
transform 1 0 2404 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1712256841
transform 1 0 2340 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1712256841
transform 1 0 1500 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1712256841
transform 1 0 1468 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4624
timestamp 1712256841
transform 1 0 1556 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4625
timestamp 1712256841
transform 1 0 1468 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1712256841
transform 1 0 1692 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4627
timestamp 1712256841
transform 1 0 1556 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1712256841
transform 1 0 1604 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4629
timestamp 1712256841
transform 1 0 1444 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4630
timestamp 1712256841
transform 1 0 3052 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4631
timestamp 1712256841
transform 1 0 2972 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1712256841
transform 1 0 2884 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1712256841
transform 1 0 2884 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4634
timestamp 1712256841
transform 1 0 2716 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1712256841
transform 1 0 2668 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4636
timestamp 1712256841
transform 1 0 2564 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4637
timestamp 1712256841
transform 1 0 2132 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4638
timestamp 1712256841
transform 1 0 2132 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4639
timestamp 1712256841
transform 1 0 2060 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4640
timestamp 1712256841
transform 1 0 2060 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4641
timestamp 1712256841
transform 1 0 1652 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4642
timestamp 1712256841
transform 1 0 1604 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4643
timestamp 1712256841
transform 1 0 2276 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4644
timestamp 1712256841
transform 1 0 2268 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4645
timestamp 1712256841
transform 1 0 2220 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4646
timestamp 1712256841
transform 1 0 2220 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4647
timestamp 1712256841
transform 1 0 2500 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4648
timestamp 1712256841
transform 1 0 2260 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4649
timestamp 1712256841
transform 1 0 2524 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4650
timestamp 1712256841
transform 1 0 2388 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4651
timestamp 1712256841
transform 1 0 2548 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4652
timestamp 1712256841
transform 1 0 2476 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4653
timestamp 1712256841
transform 1 0 2348 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4654
timestamp 1712256841
transform 1 0 2308 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4655
timestamp 1712256841
transform 1 0 2188 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4656
timestamp 1712256841
transform 1 0 2140 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4657
timestamp 1712256841
transform 1 0 2052 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4658
timestamp 1712256841
transform 1 0 2396 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4659
timestamp 1712256841
transform 1 0 2348 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4660
timestamp 1712256841
transform 1 0 2340 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4661
timestamp 1712256841
transform 1 0 2308 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4662
timestamp 1712256841
transform 1 0 2004 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4663
timestamp 1712256841
transform 1 0 2004 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4664
timestamp 1712256841
transform 1 0 1964 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4665
timestamp 1712256841
transform 1 0 2052 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4666
timestamp 1712256841
transform 1 0 1940 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4667
timestamp 1712256841
transform 1 0 2532 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4668
timestamp 1712256841
transform 1 0 2436 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4669
timestamp 1712256841
transform 1 0 2436 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4670
timestamp 1712256841
transform 1 0 2412 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4671
timestamp 1712256841
transform 1 0 2356 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4672
timestamp 1712256841
transform 1 0 2244 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4673
timestamp 1712256841
transform 1 0 2116 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4674
timestamp 1712256841
transform 1 0 1428 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4675
timestamp 1712256841
transform 1 0 1348 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4676
timestamp 1712256841
transform 1 0 2708 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1712256841
transform 1 0 1796 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4678
timestamp 1712256841
transform 1 0 1388 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4679
timestamp 1712256841
transform 1 0 2716 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4680
timestamp 1712256841
transform 1 0 2604 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4681
timestamp 1712256841
transform 1 0 2572 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4682
timestamp 1712256841
transform 1 0 2572 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4683
timestamp 1712256841
transform 1 0 2444 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4684
timestamp 1712256841
transform 1 0 2308 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4685
timestamp 1712256841
transform 1 0 2260 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4686
timestamp 1712256841
transform 1 0 1572 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4687
timestamp 1712256841
transform 1 0 1404 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1712256841
transform 1 0 2900 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4689
timestamp 1712256841
transform 1 0 2900 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4690
timestamp 1712256841
transform 1 0 2732 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4691
timestamp 1712256841
transform 1 0 2692 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4692
timestamp 1712256841
transform 1 0 2396 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4693
timestamp 1712256841
transform 1 0 2356 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4694
timestamp 1712256841
transform 1 0 2300 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4695
timestamp 1712256841
transform 1 0 2244 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4696
timestamp 1712256841
transform 1 0 2436 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4697
timestamp 1712256841
transform 1 0 2340 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1712256841
transform 1 0 2492 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4699
timestamp 1712256841
transform 1 0 2420 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4700
timestamp 1712256841
transform 1 0 2604 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4701
timestamp 1712256841
transform 1 0 2524 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4702
timestamp 1712256841
transform 1 0 2548 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4703
timestamp 1712256841
transform 1 0 2356 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4704
timestamp 1712256841
transform 1 0 2356 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4705
timestamp 1712256841
transform 1 0 2316 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4706
timestamp 1712256841
transform 1 0 2172 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4707
timestamp 1712256841
transform 1 0 2100 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1712256841
transform 1 0 2084 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4709
timestamp 1712256841
transform 1 0 2052 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4710
timestamp 1712256841
transform 1 0 2420 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4711
timestamp 1712256841
transform 1 0 2356 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4712
timestamp 1712256841
transform 1 0 2084 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4713
timestamp 1712256841
transform 1 0 2076 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4714
timestamp 1712256841
transform 1 0 2052 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4715
timestamp 1712256841
transform 1 0 2172 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4716
timestamp 1712256841
transform 1 0 2148 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4717
timestamp 1712256841
transform 1 0 2268 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4718
timestamp 1712256841
transform 1 0 2236 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4719
timestamp 1712256841
transform 1 0 2460 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4720
timestamp 1712256841
transform 1 0 2428 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4721
timestamp 1712256841
transform 1 0 2380 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4722
timestamp 1712256841
transform 1 0 2300 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4723
timestamp 1712256841
transform 1 0 2604 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4724
timestamp 1712256841
transform 1 0 1860 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4725
timestamp 1712256841
transform 1 0 1764 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4726
timestamp 1712256841
transform 1 0 1652 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1712256841
transform 1 0 1572 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1712256841
transform 1 0 1620 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4729
timestamp 1712256841
transform 1 0 1588 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1712256841
transform 1 0 2012 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1712256841
transform 1 0 1892 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4732
timestamp 1712256841
transform 1 0 1828 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4733
timestamp 1712256841
transform 1 0 1804 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4734
timestamp 1712256841
transform 1 0 1740 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4735
timestamp 1712256841
transform 1 0 1692 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4736
timestamp 1712256841
transform 1 0 1788 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4737
timestamp 1712256841
transform 1 0 1740 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1712256841
transform 1 0 1836 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1712256841
transform 1 0 1788 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4740
timestamp 1712256841
transform 1 0 1756 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4741
timestamp 1712256841
transform 1 0 1860 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4742
timestamp 1712256841
transform 1 0 1772 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4743
timestamp 1712256841
transform 1 0 1932 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4744
timestamp 1712256841
transform 1 0 1732 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4745
timestamp 1712256841
transform 1 0 2972 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4746
timestamp 1712256841
transform 1 0 2892 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4747
timestamp 1712256841
transform 1 0 2876 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4748
timestamp 1712256841
transform 1 0 2820 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4749
timestamp 1712256841
transform 1 0 2692 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4750
timestamp 1712256841
transform 1 0 2644 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4751
timestamp 1712256841
transform 1 0 2636 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4752
timestamp 1712256841
transform 1 0 2604 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4753
timestamp 1712256841
transform 1 0 2604 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4754
timestamp 1712256841
transform 1 0 2596 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4755
timestamp 1712256841
transform 1 0 2596 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4756
timestamp 1712256841
transform 1 0 2588 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4757
timestamp 1712256841
transform 1 0 2588 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4758
timestamp 1712256841
transform 1 0 2556 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4759
timestamp 1712256841
transform 1 0 2548 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4760
timestamp 1712256841
transform 1 0 2076 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4761
timestamp 1712256841
transform 1 0 1876 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4762
timestamp 1712256841
transform 1 0 1700 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4763
timestamp 1712256841
transform 1 0 2876 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4764
timestamp 1712256841
transform 1 0 2740 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4765
timestamp 1712256841
transform 1 0 2732 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4766
timestamp 1712256841
transform 1 0 2628 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4767
timestamp 1712256841
transform 1 0 2604 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4768
timestamp 1712256841
transform 1 0 2596 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4769
timestamp 1712256841
transform 1 0 2516 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4770
timestamp 1712256841
transform 1 0 2516 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4771
timestamp 1712256841
transform 1 0 2004 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4772
timestamp 1712256841
transform 1 0 1780 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4773
timestamp 1712256841
transform 1 0 1716 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4774
timestamp 1712256841
transform 1 0 1444 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4775
timestamp 1712256841
transform 1 0 1348 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4776
timestamp 1712256841
transform 1 0 2084 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1712256841
transform 1 0 1980 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4778
timestamp 1712256841
transform 1 0 2004 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4779
timestamp 1712256841
transform 1 0 1956 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4780
timestamp 1712256841
transform 1 0 2332 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1712256841
transform 1 0 2164 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4782
timestamp 1712256841
transform 1 0 2244 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4783
timestamp 1712256841
transform 1 0 2212 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4784
timestamp 1712256841
transform 1 0 2052 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4785
timestamp 1712256841
transform 1 0 1884 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1712256841
transform 1 0 1860 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1712256841
transform 1 0 1908 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4788
timestamp 1712256841
transform 1 0 1884 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4789
timestamp 1712256841
transform 1 0 2068 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1712256841
transform 1 0 1940 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4791
timestamp 1712256841
transform 1 0 2228 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4792
timestamp 1712256841
transform 1 0 2140 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4793
timestamp 1712256841
transform 1 0 2444 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4794
timestamp 1712256841
transform 1 0 2180 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4795
timestamp 1712256841
transform 1 0 3068 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1712256841
transform 1 0 3004 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4797
timestamp 1712256841
transform 1 0 2820 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4798
timestamp 1712256841
transform 1 0 2708 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4799
timestamp 1712256841
transform 1 0 2708 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4800
timestamp 1712256841
transform 1 0 2500 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4801
timestamp 1712256841
transform 1 0 2428 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4802
timestamp 1712256841
transform 1 0 2196 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4803
timestamp 1712256841
transform 1 0 2140 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4804
timestamp 1712256841
transform 1 0 2444 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4805
timestamp 1712256841
transform 1 0 2236 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4806
timestamp 1712256841
transform 1 0 2164 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4807
timestamp 1712256841
transform 1 0 2140 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4808
timestamp 1712256841
transform 1 0 2276 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4809
timestamp 1712256841
transform 1 0 2220 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4810
timestamp 1712256841
transform 1 0 2460 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4811
timestamp 1712256841
transform 1 0 2244 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4812
timestamp 1712256841
transform 1 0 2380 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4813
timestamp 1712256841
transform 1 0 2300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4814
timestamp 1712256841
transform 1 0 2164 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1712256841
transform 1 0 2148 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4816
timestamp 1712256841
transform 1 0 2188 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1712256841
transform 1 0 2164 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4818
timestamp 1712256841
transform 1 0 2364 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4819
timestamp 1712256841
transform 1 0 2356 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4820
timestamp 1712256841
transform 1 0 2340 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4821
timestamp 1712256841
transform 1 0 2300 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4822
timestamp 1712256841
transform 1 0 2372 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1712256841
transform 1 0 2260 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4824
timestamp 1712256841
transform 1 0 2412 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1712256841
transform 1 0 2340 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4826
timestamp 1712256841
transform 1 0 2476 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4827
timestamp 1712256841
transform 1 0 2404 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4828
timestamp 1712256841
transform 1 0 2476 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4829
timestamp 1712256841
transform 1 0 2460 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1712256841
transform 1 0 2812 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1712256841
transform 1 0 2748 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4832
timestamp 1712256841
transform 1 0 2524 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4833
timestamp 1712256841
transform 1 0 2508 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4834
timestamp 1712256841
transform 1 0 2412 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4835
timestamp 1712256841
transform 1 0 2372 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4836
timestamp 1712256841
transform 1 0 2332 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1712256841
transform 1 0 2932 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4838
timestamp 1712256841
transform 1 0 2924 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4839
timestamp 1712256841
transform 1 0 2916 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4840
timestamp 1712256841
transform 1 0 2692 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4841
timestamp 1712256841
transform 1 0 2524 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4842
timestamp 1712256841
transform 1 0 2468 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4843
timestamp 1712256841
transform 1 0 2452 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4844
timestamp 1712256841
transform 1 0 2452 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4845
timestamp 1712256841
transform 1 0 2436 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4846
timestamp 1712256841
transform 1 0 2404 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4847
timestamp 1712256841
transform 1 0 2684 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4848
timestamp 1712256841
transform 1 0 2452 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4849
timestamp 1712256841
transform 1 0 2364 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4850
timestamp 1712256841
transform 1 0 2308 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4851
timestamp 1712256841
transform 1 0 2412 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4852
timestamp 1712256841
transform 1 0 2388 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4853
timestamp 1712256841
transform 1 0 2572 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4854
timestamp 1712256841
transform 1 0 2556 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4855
timestamp 1712256841
transform 1 0 2604 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1712256841
transform 1 0 2460 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4857
timestamp 1712256841
transform 1 0 2692 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4858
timestamp 1712256841
transform 1 0 2628 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4859
timestamp 1712256841
transform 1 0 2748 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4860
timestamp 1712256841
transform 1 0 2620 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4861
timestamp 1712256841
transform 1 0 2564 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4862
timestamp 1712256841
transform 1 0 2524 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4863
timestamp 1712256841
transform 1 0 2628 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1712256841
transform 1 0 2588 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4865
timestamp 1712256841
transform 1 0 2548 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4866
timestamp 1712256841
transform 1 0 2116 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4867
timestamp 1712256841
transform 1 0 2540 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4868
timestamp 1712256841
transform 1 0 2516 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4869
timestamp 1712256841
transform 1 0 2692 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4870
timestamp 1712256841
transform 1 0 2540 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4871
timestamp 1712256841
transform 1 0 2676 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4872
timestamp 1712256841
transform 1 0 2652 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4873
timestamp 1712256841
transform 1 0 2628 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4874
timestamp 1712256841
transform 1 0 2844 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4875
timestamp 1712256841
transform 1 0 2716 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4876
timestamp 1712256841
transform 1 0 2716 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4877
timestamp 1712256841
transform 1 0 2716 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4878
timestamp 1712256841
transform 1 0 2676 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4879
timestamp 1712256841
transform 1 0 2652 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4880
timestamp 1712256841
transform 1 0 2604 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4881
timestamp 1712256841
transform 1 0 2092 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4882
timestamp 1712256841
transform 1 0 2028 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4883
timestamp 1712256841
transform 1 0 3316 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4884
timestamp 1712256841
transform 1 0 3156 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4885
timestamp 1712256841
transform 1 0 3140 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4886
timestamp 1712256841
transform 1 0 2676 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4887
timestamp 1712256841
transform 1 0 2724 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4888
timestamp 1712256841
transform 1 0 2540 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4889
timestamp 1712256841
transform 1 0 2044 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4890
timestamp 1712256841
transform 1 0 2044 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4891
timestamp 1712256841
transform 1 0 1980 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4892
timestamp 1712256841
transform 1 0 1668 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4893
timestamp 1712256841
transform 1 0 1652 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4894
timestamp 1712256841
transform 1 0 3196 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4895
timestamp 1712256841
transform 1 0 3132 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4896
timestamp 1712256841
transform 1 0 3284 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4897
timestamp 1712256841
transform 1 0 3180 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4898
timestamp 1712256841
transform 1 0 2780 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4899
timestamp 1712256841
transform 1 0 2676 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4900
timestamp 1712256841
transform 1 0 2636 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4901
timestamp 1712256841
transform 1 0 2932 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4902
timestamp 1712256841
transform 1 0 2860 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4903
timestamp 1712256841
transform 1 0 2924 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4904
timestamp 1712256841
transform 1 0 2900 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4905
timestamp 1712256841
transform 1 0 2996 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4906
timestamp 1712256841
transform 1 0 2908 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4907
timestamp 1712256841
transform 1 0 3020 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4908
timestamp 1712256841
transform 1 0 2988 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4909
timestamp 1712256841
transform 1 0 3036 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4910
timestamp 1712256841
transform 1 0 2996 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4911
timestamp 1712256841
transform 1 0 2972 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1712256841
transform 1 0 2948 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4913
timestamp 1712256841
transform 1 0 3260 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4914
timestamp 1712256841
transform 1 0 3260 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4915
timestamp 1712256841
transform 1 0 3108 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4916
timestamp 1712256841
transform 1 0 3076 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4917
timestamp 1712256841
transform 1 0 2956 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4918
timestamp 1712256841
transform 1 0 3044 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4919
timestamp 1712256841
transform 1 0 2980 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4920
timestamp 1712256841
transform 1 0 2972 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4921
timestamp 1712256841
transform 1 0 2956 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1712256841
transform 1 0 2932 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4923
timestamp 1712256841
transform 1 0 2908 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4924
timestamp 1712256841
transform 1 0 3092 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4925
timestamp 1712256841
transform 1 0 3020 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4926
timestamp 1712256841
transform 1 0 3036 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4927
timestamp 1712256841
transform 1 0 2804 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4928
timestamp 1712256841
transform 1 0 3092 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4929
timestamp 1712256841
transform 1 0 2916 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4930
timestamp 1712256841
transform 1 0 3020 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4931
timestamp 1712256841
transform 1 0 2996 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4932
timestamp 1712256841
transform 1 0 2996 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4933
timestamp 1712256841
transform 1 0 2956 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4934
timestamp 1712256841
transform 1 0 2956 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4935
timestamp 1712256841
transform 1 0 2940 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4936
timestamp 1712256841
transform 1 0 2956 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4937
timestamp 1712256841
transform 1 0 2932 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1712256841
transform 1 0 2988 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4939
timestamp 1712256841
transform 1 0 2924 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4940
timestamp 1712256841
transform 1 0 3092 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4941
timestamp 1712256841
transform 1 0 2972 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4942
timestamp 1712256841
transform 1 0 2860 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4943
timestamp 1712256841
transform 1 0 3276 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1712256841
transform 1 0 3268 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4945
timestamp 1712256841
transform 1 0 3204 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1712256841
transform 1 0 3204 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4947
timestamp 1712256841
transform 1 0 3204 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4948
timestamp 1712256841
transform 1 0 2948 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4949
timestamp 1712256841
transform 1 0 2876 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4950
timestamp 1712256841
transform 1 0 2844 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4951
timestamp 1712256841
transform 1 0 3156 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4952
timestamp 1712256841
transform 1 0 3052 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4953
timestamp 1712256841
transform 1 0 3172 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4954
timestamp 1712256841
transform 1 0 3116 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4955
timestamp 1712256841
transform 1 0 3108 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4956
timestamp 1712256841
transform 1 0 3092 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4957
timestamp 1712256841
transform 1 0 2724 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4958
timestamp 1712256841
transform 1 0 2668 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1712256841
transform 1 0 2604 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4960
timestamp 1712256841
transform 1 0 2596 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4961
timestamp 1712256841
transform 1 0 2516 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4962
timestamp 1712256841
transform 1 0 2780 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4963
timestamp 1712256841
transform 1 0 2740 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4964
timestamp 1712256841
transform 1 0 3068 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4965
timestamp 1712256841
transform 1 0 3052 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4966
timestamp 1712256841
transform 1 0 3052 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4967
timestamp 1712256841
transform 1 0 2812 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4968
timestamp 1712256841
transform 1 0 2996 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4969
timestamp 1712256841
transform 1 0 2948 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4970
timestamp 1712256841
transform 1 0 3108 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4971
timestamp 1712256841
transform 1 0 3028 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4972
timestamp 1712256841
transform 1 0 2964 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4973
timestamp 1712256841
transform 1 0 3156 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4974
timestamp 1712256841
transform 1 0 3092 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1712256841
transform 1 0 3092 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4976
timestamp 1712256841
transform 1 0 3044 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4977
timestamp 1712256841
transform 1 0 2620 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4978
timestamp 1712256841
transform 1 0 2548 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_4979
timestamp 1712256841
transform 1 0 3108 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4980
timestamp 1712256841
transform 1 0 3068 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4981
timestamp 1712256841
transform 1 0 3052 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1712256841
transform 1 0 2916 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1712256841
transform 1 0 3108 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4984
timestamp 1712256841
transform 1 0 3092 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4985
timestamp 1712256841
transform 1 0 2892 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4986
timestamp 1712256841
transform 1 0 2860 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4987
timestamp 1712256841
transform 1 0 3028 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4988
timestamp 1712256841
transform 1 0 2868 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4989
timestamp 1712256841
transform 1 0 3060 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4990
timestamp 1712256841
transform 1 0 3012 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4991
timestamp 1712256841
transform 1 0 2612 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4992
timestamp 1712256841
transform 1 0 2532 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4993
timestamp 1712256841
transform 1 0 2956 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4994
timestamp 1712256841
transform 1 0 2868 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4995
timestamp 1712256841
transform 1 0 3068 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4996
timestamp 1712256841
transform 1 0 2924 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4997
timestamp 1712256841
transform 1 0 2844 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4998
timestamp 1712256841
transform 1 0 3172 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4999
timestamp 1712256841
transform 1 0 2884 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5000
timestamp 1712256841
transform 1 0 2868 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5001
timestamp 1712256841
transform 1 0 2908 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5002
timestamp 1712256841
transform 1 0 2852 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5003
timestamp 1712256841
transform 1 0 2876 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5004
timestamp 1712256841
transform 1 0 2748 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5005
timestamp 1712256841
transform 1 0 2788 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5006
timestamp 1712256841
transform 1 0 2748 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5007
timestamp 1712256841
transform 1 0 2908 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5008
timestamp 1712256841
transform 1 0 2860 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5009
timestamp 1712256841
transform 1 0 2868 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5010
timestamp 1712256841
transform 1 0 2812 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5011
timestamp 1712256841
transform 1 0 2908 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5012
timestamp 1712256841
transform 1 0 2836 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5013
timestamp 1712256841
transform 1 0 2716 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5014
timestamp 1712256841
transform 1 0 2620 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5015
timestamp 1712256841
transform 1 0 2876 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5016
timestamp 1712256841
transform 1 0 2844 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5017
timestamp 1712256841
transform 1 0 2908 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5018
timestamp 1712256841
transform 1 0 2844 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5019
timestamp 1712256841
transform 1 0 2884 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5020
timestamp 1712256841
transform 1 0 2732 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5021
timestamp 1712256841
transform 1 0 2900 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5022
timestamp 1712256841
transform 1 0 2852 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5023
timestamp 1712256841
transform 1 0 2924 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5024
timestamp 1712256841
transform 1 0 2868 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5025
timestamp 1712256841
transform 1 0 3228 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5026
timestamp 1712256841
transform 1 0 3204 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5027
timestamp 1712256841
transform 1 0 2732 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5028
timestamp 1712256841
transform 1 0 2604 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5029
timestamp 1712256841
transform 1 0 2900 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5030
timestamp 1712256841
transform 1 0 2796 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5031
timestamp 1712256841
transform 1 0 2820 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5032
timestamp 1712256841
transform 1 0 2636 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5033
timestamp 1712256841
transform 1 0 2820 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5034
timestamp 1712256841
transform 1 0 2772 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5035
timestamp 1712256841
transform 1 0 2820 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5036
timestamp 1712256841
transform 1 0 2812 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5037
timestamp 1712256841
transform 1 0 2764 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5038
timestamp 1712256841
transform 1 0 2764 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1712256841
transform 1 0 2804 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5040
timestamp 1712256841
transform 1 0 2804 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5041
timestamp 1712256841
transform 1 0 2788 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5042
timestamp 1712256841
transform 1 0 2756 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5043
timestamp 1712256841
transform 1 0 2676 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5044
timestamp 1712256841
transform 1 0 2492 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5045
timestamp 1712256841
transform 1 0 2780 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_5046
timestamp 1712256841
transform 1 0 2740 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_5047
timestamp 1712256841
transform 1 0 3180 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_5048
timestamp 1712256841
transform 1 0 3092 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_5049
timestamp 1712256841
transform 1 0 3332 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5050
timestamp 1712256841
transform 1 0 3196 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5051
timestamp 1712256841
transform 1 0 3436 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5052
timestamp 1712256841
transform 1 0 3324 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5053
timestamp 1712256841
transform 1 0 3076 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5054
timestamp 1712256841
transform 1 0 2892 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5055
timestamp 1712256841
transform 1 0 3404 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5056
timestamp 1712256841
transform 1 0 3364 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5057
timestamp 1712256841
transform 1 0 3396 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5058
timestamp 1712256841
transform 1 0 3372 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5059
timestamp 1712256841
transform 1 0 3372 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5060
timestamp 1712256841
transform 1 0 3348 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5061
timestamp 1712256841
transform 1 0 3324 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5062
timestamp 1712256841
transform 1 0 3324 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5063
timestamp 1712256841
transform 1 0 3428 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5064
timestamp 1712256841
transform 1 0 3404 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5065
timestamp 1712256841
transform 1 0 3348 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5066
timestamp 1712256841
transform 1 0 3308 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5067
timestamp 1712256841
transform 1 0 3140 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_5068
timestamp 1712256841
transform 1 0 3140 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5069
timestamp 1712256841
transform 1 0 2956 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5070
timestamp 1712256841
transform 1 0 2916 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5071
timestamp 1712256841
transform 1 0 3412 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5072
timestamp 1712256841
transform 1 0 3340 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5073
timestamp 1712256841
transform 1 0 3284 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5074
timestamp 1712256841
transform 1 0 3284 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5075
timestamp 1712256841
transform 1 0 3180 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5076
timestamp 1712256841
transform 1 0 2980 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5077
timestamp 1712256841
transform 1 0 3340 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_5078
timestamp 1712256841
transform 1 0 3300 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_5079
timestamp 1712256841
transform 1 0 3428 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5080
timestamp 1712256841
transform 1 0 3388 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5081
timestamp 1712256841
transform 1 0 3228 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5082
timestamp 1712256841
transform 1 0 3180 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5083
timestamp 1712256841
transform 1 0 3356 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5084
timestamp 1712256841
transform 1 0 3300 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5085
timestamp 1712256841
transform 1 0 3348 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5086
timestamp 1712256841
transform 1 0 3228 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5087
timestamp 1712256841
transform 1 0 3260 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5088
timestamp 1712256841
transform 1 0 3236 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5089
timestamp 1712256841
transform 1 0 3396 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5090
timestamp 1712256841
transform 1 0 3340 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5091
timestamp 1712256841
transform 1 0 3412 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5092
timestamp 1712256841
transform 1 0 3388 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5093
timestamp 1712256841
transform 1 0 3388 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5094
timestamp 1712256841
transform 1 0 3260 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5095
timestamp 1712256841
transform 1 0 3300 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5096
timestamp 1712256841
transform 1 0 3236 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5097
timestamp 1712256841
transform 1 0 3196 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5098
timestamp 1712256841
transform 1 0 3132 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1712256841
transform 1 0 3212 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5100
timestamp 1712256841
transform 1 0 3180 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5101
timestamp 1712256841
transform 1 0 3260 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5102
timestamp 1712256841
transform 1 0 3188 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5103
timestamp 1712256841
transform 1 0 3196 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5104
timestamp 1712256841
transform 1 0 3052 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5105
timestamp 1712256841
transform 1 0 2604 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5106
timestamp 1712256841
transform 1 0 2468 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5107
timestamp 1712256841
transform 1 0 2356 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5108
timestamp 1712256841
transform 1 0 2316 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5109
timestamp 1712256841
transform 1 0 1892 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5110
timestamp 1712256841
transform 1 0 1804 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5111
timestamp 1712256841
transform 1 0 1732 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5112
timestamp 1712256841
transform 1 0 1684 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5113
timestamp 1712256841
transform 1 0 1148 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5114
timestamp 1712256841
transform 1 0 1044 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5115
timestamp 1712256841
transform 1 0 1068 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5116
timestamp 1712256841
transform 1 0 940 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5117
timestamp 1712256841
transform 1 0 444 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5118
timestamp 1712256841
transform 1 0 348 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5119
timestamp 1712256841
transform 1 0 700 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5120
timestamp 1712256841
transform 1 0 548 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5121
timestamp 1712256841
transform 1 0 3180 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5122
timestamp 1712256841
transform 1 0 2948 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5123
timestamp 1712256841
transform 1 0 2916 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_5124
timestamp 1712256841
transform 1 0 2796 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_5125
timestamp 1712256841
transform 1 0 2780 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5126
timestamp 1712256841
transform 1 0 2764 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5127
timestamp 1712256841
transform 1 0 2740 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5128
timestamp 1712256841
transform 1 0 2428 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5129
timestamp 1712256841
transform 1 0 2284 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5130
timestamp 1712256841
transform 1 0 2180 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5131
timestamp 1712256841
transform 1 0 2132 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5132
timestamp 1712256841
transform 1 0 2044 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5133
timestamp 1712256841
transform 1 0 2140 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5134
timestamp 1712256841
transform 1 0 1300 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5135
timestamp 1712256841
transform 1 0 2332 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5136
timestamp 1712256841
transform 1 0 2180 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5137
timestamp 1712256841
transform 1 0 1852 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_5138
timestamp 1712256841
transform 1 0 1636 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_5139
timestamp 1712256841
transform 1 0 1364 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_5140
timestamp 1712256841
transform 1 0 1364 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5141
timestamp 1712256841
transform 1 0 1252 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5142
timestamp 1712256841
transform 1 0 1068 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5143
timestamp 1712256841
transform 1 0 1292 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5144
timestamp 1712256841
transform 1 0 1188 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5145
timestamp 1712256841
transform 1 0 948 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5146
timestamp 1712256841
transform 1 0 932 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5147
timestamp 1712256841
transform 1 0 868 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5148
timestamp 1712256841
transform 1 0 1316 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5149
timestamp 1712256841
transform 1 0 1228 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5150
timestamp 1712256841
transform 1 0 1356 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5151
timestamp 1712256841
transform 1 0 1308 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5152
timestamp 1712256841
transform 1 0 972 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5153
timestamp 1712256841
transform 1 0 804 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5154
timestamp 1712256841
transform 1 0 1996 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5155
timestamp 1712256841
transform 1 0 1764 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5156
timestamp 1712256841
transform 1 0 2004 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5157
timestamp 1712256841
transform 1 0 1972 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1712256841
transform 1 0 1964 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5159
timestamp 1712256841
transform 1 0 1924 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5160
timestamp 1712256841
transform 1 0 1844 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5161
timestamp 1712256841
transform 1 0 1556 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5162
timestamp 1712256841
transform 1 0 1508 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5163
timestamp 1712256841
transform 1 0 2108 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5164
timestamp 1712256841
transform 1 0 2044 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5165
timestamp 1712256841
transform 1 0 2444 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5166
timestamp 1712256841
transform 1 0 2364 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5167
timestamp 1712256841
transform 1 0 2060 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5168
timestamp 1712256841
transform 1 0 2036 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5169
timestamp 1712256841
transform 1 0 1956 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5170
timestamp 1712256841
transform 1 0 3164 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5171
timestamp 1712256841
transform 1 0 3068 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5172
timestamp 1712256841
transform 1 0 3020 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5173
timestamp 1712256841
transform 1 0 3020 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5174
timestamp 1712256841
transform 1 0 2524 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5175
timestamp 1712256841
transform 1 0 2460 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5176
timestamp 1712256841
transform 1 0 2388 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5177
timestamp 1712256841
transform 1 0 3052 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1712256841
transform 1 0 2860 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5179
timestamp 1712256841
transform 1 0 2860 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_5180
timestamp 1712256841
transform 1 0 972 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5181
timestamp 1712256841
transform 1 0 860 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5182
timestamp 1712256841
transform 1 0 620 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5183
timestamp 1712256841
transform 1 0 500 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5184
timestamp 1712256841
transform 1 0 468 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5185
timestamp 1712256841
transform 1 0 436 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5186
timestamp 1712256841
transform 1 0 348 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5187
timestamp 1712256841
transform 1 0 284 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5188
timestamp 1712256841
transform 1 0 2916 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5189
timestamp 1712256841
transform 1 0 2868 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5190
timestamp 1712256841
transform 1 0 2860 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1712256841
transform 1 0 2764 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5192
timestamp 1712256841
transform 1 0 2764 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5193
timestamp 1712256841
transform 1 0 2644 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5194
timestamp 1712256841
transform 1 0 3060 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5195
timestamp 1712256841
transform 1 0 2972 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5196
timestamp 1712256841
transform 1 0 2636 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5197
timestamp 1712256841
transform 1 0 2572 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5198
timestamp 1712256841
transform 1 0 2540 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5199
timestamp 1712256841
transform 1 0 2484 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5200
timestamp 1712256841
transform 1 0 2420 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5201
timestamp 1712256841
transform 1 0 2900 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5202
timestamp 1712256841
transform 1 0 2796 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5203
timestamp 1712256841
transform 1 0 2748 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5204
timestamp 1712256841
transform 1 0 2692 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5205
timestamp 1712256841
transform 1 0 2716 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5206
timestamp 1712256841
transform 1 0 2596 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5207
timestamp 1712256841
transform 1 0 2516 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5208
timestamp 1712256841
transform 1 0 2476 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5209
timestamp 1712256841
transform 1 0 2204 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5210
timestamp 1712256841
transform 1 0 2772 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5211
timestamp 1712256841
transform 1 0 2684 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5212
timestamp 1712256841
transform 1 0 2604 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5213
timestamp 1712256841
transform 1 0 2524 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5214
timestamp 1712256841
transform 1 0 2172 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5215
timestamp 1712256841
transform 1 0 2036 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5216
timestamp 1712256841
transform 1 0 2372 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5217
timestamp 1712256841
transform 1 0 2348 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5218
timestamp 1712256841
transform 1 0 2332 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5219
timestamp 1712256841
transform 1 0 2276 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5220
timestamp 1712256841
transform 1 0 2212 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5221
timestamp 1712256841
transform 1 0 2180 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5222
timestamp 1712256841
transform 1 0 2028 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5223
timestamp 1712256841
transform 1 0 2420 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5224
timestamp 1712256841
transform 1 0 2340 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5225
timestamp 1712256841
transform 1 0 2340 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5226
timestamp 1712256841
transform 1 0 2268 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5227
timestamp 1712256841
transform 1 0 2148 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5228
timestamp 1712256841
transform 1 0 2020 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5229
timestamp 1712256841
transform 1 0 2244 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5230
timestamp 1712256841
transform 1 0 2124 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5231
timestamp 1712256841
transform 1 0 2060 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5232
timestamp 1712256841
transform 1 0 1924 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5233
timestamp 1712256841
transform 1 0 2348 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5234
timestamp 1712256841
transform 1 0 2172 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5235
timestamp 1712256841
transform 1 0 2340 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5236
timestamp 1712256841
transform 1 0 2284 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5237
timestamp 1712256841
transform 1 0 2236 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5238
timestamp 1712256841
transform 1 0 2132 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5239
timestamp 1712256841
transform 1 0 1988 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5240
timestamp 1712256841
transform 1 0 2308 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_5241
timestamp 1712256841
transform 1 0 2236 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_5242
timestamp 1712256841
transform 1 0 2228 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5243
timestamp 1712256841
transform 1 0 2180 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5244
timestamp 1712256841
transform 1 0 2252 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5245
timestamp 1712256841
transform 1 0 2220 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5246
timestamp 1712256841
transform 1 0 2124 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5247
timestamp 1712256841
transform 1 0 2084 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5248
timestamp 1712256841
transform 1 0 2020 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5249
timestamp 1712256841
transform 1 0 1868 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5250
timestamp 1712256841
transform 1 0 2220 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5251
timestamp 1712256841
transform 1 0 2116 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5252
timestamp 1712256841
transform 1 0 1932 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5253
timestamp 1712256841
transform 1 0 1980 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5254
timestamp 1712256841
transform 1 0 1924 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5255
timestamp 1712256841
transform 1 0 1836 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5256
timestamp 1712256841
transform 1 0 1780 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5257
timestamp 1712256841
transform 1 0 1724 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5258
timestamp 1712256841
transform 1 0 1852 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5259
timestamp 1712256841
transform 1 0 1812 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5260
timestamp 1712256841
transform 1 0 1868 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5261
timestamp 1712256841
transform 1 0 1772 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1712256841
transform 1 0 1668 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5263
timestamp 1712256841
transform 1 0 1956 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5264
timestamp 1712256841
transform 1 0 1900 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5265
timestamp 1712256841
transform 1 0 1756 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5266
timestamp 1712256841
transform 1 0 1660 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5267
timestamp 1712256841
transform 1 0 1756 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5268
timestamp 1712256841
transform 1 0 1708 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5269
timestamp 1712256841
transform 1 0 1732 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5270
timestamp 1712256841
transform 1 0 1604 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5271
timestamp 1712256841
transform 1 0 1748 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1712256841
transform 1 0 1708 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5273
timestamp 1712256841
transform 1 0 1964 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5274
timestamp 1712256841
transform 1 0 1828 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5275
timestamp 1712256841
transform 1 0 1820 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5276
timestamp 1712256841
transform 1 0 1620 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1712256841
transform 1 0 1548 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5278
timestamp 1712256841
transform 1 0 1780 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5279
timestamp 1712256841
transform 1 0 1556 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1712256841
transform 1 0 1524 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1712256841
transform 1 0 1548 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5282
timestamp 1712256841
transform 1 0 1444 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5283
timestamp 1712256841
transform 1 0 1636 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5284
timestamp 1712256841
transform 1 0 1524 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1712256841
transform 1 0 1380 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1712256841
transform 1 0 1644 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1712256841
transform 1 0 1580 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5288
timestamp 1712256841
transform 1 0 1428 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5289
timestamp 1712256841
transform 1 0 1348 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5290
timestamp 1712256841
transform 1 0 1420 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5291
timestamp 1712256841
transform 1 0 1340 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5292
timestamp 1712256841
transform 1 0 1604 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5293
timestamp 1712256841
transform 1 0 1436 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5294
timestamp 1712256841
transform 1 0 1404 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1712256841
transform 1 0 1316 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5296
timestamp 1712256841
transform 1 0 1604 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5297
timestamp 1712256841
transform 1 0 1404 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1712256841
transform 1 0 1436 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1712256841
transform 1 0 1236 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1712256841
transform 1 0 1540 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1712256841
transform 1 0 1476 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5302
timestamp 1712256841
transform 1 0 1588 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1712256841
transform 1 0 1492 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5304
timestamp 1712256841
transform 1 0 1404 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5305
timestamp 1712256841
transform 1 0 1172 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5306
timestamp 1712256841
transform 1 0 1092 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5307
timestamp 1712256841
transform 1 0 1428 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5308
timestamp 1712256841
transform 1 0 1148 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5309
timestamp 1712256841
transform 1 0 1148 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5310
timestamp 1712256841
transform 1 0 1076 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5311
timestamp 1712256841
transform 1 0 1020 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5312
timestamp 1712256841
transform 1 0 236 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5313
timestamp 1712256841
transform 1 0 1132 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5314
timestamp 1712256841
transform 1 0 1012 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5315
timestamp 1712256841
transform 1 0 1132 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5316
timestamp 1712256841
transform 1 0 1084 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5317
timestamp 1712256841
transform 1 0 628 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5318
timestamp 1712256841
transform 1 0 276 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5319
timestamp 1712256841
transform 1 0 1140 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5320
timestamp 1712256841
transform 1 0 620 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5321
timestamp 1712256841
transform 1 0 756 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5322
timestamp 1712256841
transform 1 0 332 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5323
timestamp 1712256841
transform 1 0 1012 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5324
timestamp 1712256841
transform 1 0 748 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5325
timestamp 1712256841
transform 1 0 1100 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1712256841
transform 1 0 916 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5327
timestamp 1712256841
transform 1 0 908 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5328
timestamp 1712256841
transform 1 0 740 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1712256841
transform 1 0 1132 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5330
timestamp 1712256841
transform 1 0 884 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5331
timestamp 1712256841
transform 1 0 604 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5332
timestamp 1712256841
transform 1 0 564 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5333
timestamp 1712256841
transform 1 0 532 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5334
timestamp 1712256841
transform 1 0 604 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5335
timestamp 1712256841
transform 1 0 300 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5336
timestamp 1712256841
transform 1 0 740 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5337
timestamp 1712256841
transform 1 0 652 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5338
timestamp 1712256841
transform 1 0 988 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5339
timestamp 1712256841
transform 1 0 844 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5340
timestamp 1712256841
transform 1 0 804 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5341
timestamp 1712256841
transform 1 0 732 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5342
timestamp 1712256841
transform 1 0 660 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5343
timestamp 1712256841
transform 1 0 596 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5344
timestamp 1712256841
transform 1 0 524 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5345
timestamp 1712256841
transform 1 0 668 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5346
timestamp 1712256841
transform 1 0 596 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5347
timestamp 1712256841
transform 1 0 524 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5348
timestamp 1712256841
transform 1 0 412 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5349
timestamp 1712256841
transform 1 0 628 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5350
timestamp 1712256841
transform 1 0 556 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5351
timestamp 1712256841
transform 1 0 564 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5352
timestamp 1712256841
transform 1 0 500 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5353
timestamp 1712256841
transform 1 0 684 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5354
timestamp 1712256841
transform 1 0 612 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_5355
timestamp 1712256841
transform 1 0 908 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5356
timestamp 1712256841
transform 1 0 828 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5357
timestamp 1712256841
transform 1 0 820 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5358
timestamp 1712256841
transform 1 0 788 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5359
timestamp 1712256841
transform 1 0 788 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5360
timestamp 1712256841
transform 1 0 892 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5361
timestamp 1712256841
transform 1 0 828 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5362
timestamp 1712256841
transform 1 0 796 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5363
timestamp 1712256841
transform 1 0 780 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5364
timestamp 1712256841
transform 1 0 732 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5365
timestamp 1712256841
transform 1 0 668 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5366
timestamp 1712256841
transform 1 0 836 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5367
timestamp 1712256841
transform 1 0 732 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5368
timestamp 1712256841
transform 1 0 956 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5369
timestamp 1712256841
transform 1 0 868 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5370
timestamp 1712256841
transform 1 0 836 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5371
timestamp 1712256841
transform 1 0 804 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5372
timestamp 1712256841
transform 1 0 692 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5373
timestamp 1712256841
transform 1 0 644 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5374
timestamp 1712256841
transform 1 0 532 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5375
timestamp 1712256841
transform 1 0 716 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5376
timestamp 1712256841
transform 1 0 636 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5377
timestamp 1712256841
transform 1 0 852 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5378
timestamp 1712256841
transform 1 0 804 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5379
timestamp 1712256841
transform 1 0 1044 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5380
timestamp 1712256841
transform 1 0 996 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5381
timestamp 1712256841
transform 1 0 988 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5382
timestamp 1712256841
transform 1 0 844 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5383
timestamp 1712256841
transform 1 0 1204 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5384
timestamp 1712256841
transform 1 0 964 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1712256841
transform 1 0 860 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5386
timestamp 1712256841
transform 1 0 764 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5387
timestamp 1712256841
transform 1 0 1876 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5388
timestamp 1712256841
transform 1 0 1788 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5389
timestamp 1712256841
transform 1 0 1692 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5390
timestamp 1712256841
transform 1 0 1348 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5391
timestamp 1712256841
transform 1 0 3116 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_5392
timestamp 1712256841
transform 1 0 2964 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_5393
timestamp 1712256841
transform 1 0 2828 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_5394
timestamp 1712256841
transform 1 0 2684 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_5395
timestamp 1712256841
transform 1 0 2676 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5396
timestamp 1712256841
transform 1 0 2396 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5397
timestamp 1712256841
transform 1 0 2236 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5398
timestamp 1712256841
transform 1 0 2044 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5399
timestamp 1712256841
transform 1 0 1844 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5400
timestamp 1712256841
transform 1 0 1116 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5401
timestamp 1712256841
transform 1 0 868 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5402
timestamp 1712256841
transform 1 0 628 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5403
timestamp 1712256841
transform 1 0 628 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5404
timestamp 1712256841
transform 1 0 564 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5405
timestamp 1712256841
transform 1 0 484 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5406
timestamp 1712256841
transform 1 0 460 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5407
timestamp 1712256841
transform 1 0 3100 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5408
timestamp 1712256841
transform 1 0 2844 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5409
timestamp 1712256841
transform 1 0 2628 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5410
timestamp 1712256841
transform 1 0 2428 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5411
timestamp 1712256841
transform 1 0 2300 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5412
timestamp 1712256841
transform 1 0 2300 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5413
timestamp 1712256841
transform 1 0 2036 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5414
timestamp 1712256841
transform 1 0 2036 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5415
timestamp 1712256841
transform 1 0 1908 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5416
timestamp 1712256841
transform 1 0 1716 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5417
timestamp 1712256841
transform 1 0 1588 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5418
timestamp 1712256841
transform 1 0 1292 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5419
timestamp 1712256841
transform 1 0 1924 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5420
timestamp 1712256841
transform 1 0 1820 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5421
timestamp 1712256841
transform 1 0 2156 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5422
timestamp 1712256841
transform 1 0 1956 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5423
timestamp 1712256841
transform 1 0 3140 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5424
timestamp 1712256841
transform 1 0 3044 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5425
timestamp 1712256841
transform 1 0 2620 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5426
timestamp 1712256841
transform 1 0 2540 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5427
timestamp 1712256841
transform 1 0 2708 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5428
timestamp 1712256841
transform 1 0 2636 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5429
timestamp 1712256841
transform 1 0 2500 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5430
timestamp 1712256841
transform 1 0 2412 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5431
timestamp 1712256841
transform 1 0 2084 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5432
timestamp 1712256841
transform 1 0 2004 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1712256841
transform 1 0 2308 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5434
timestamp 1712256841
transform 1 0 2228 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5435
timestamp 1712256841
transform 1 0 2060 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5436
timestamp 1712256841
transform 1 0 1988 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5437
timestamp 1712256841
transform 1 0 1780 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5438
timestamp 1712256841
transform 1 0 1724 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5439
timestamp 1712256841
transform 1 0 1908 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5440
timestamp 1712256841
transform 1 0 1852 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5441
timestamp 1712256841
transform 1 0 1460 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5442
timestamp 1712256841
transform 1 0 1396 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5443
timestamp 1712256841
transform 1 0 1420 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5444
timestamp 1712256841
transform 1 0 1340 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5445
timestamp 1712256841
transform 1 0 1252 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5446
timestamp 1712256841
transform 1 0 1164 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5447
timestamp 1712256841
transform 1 0 1188 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5448
timestamp 1712256841
transform 1 0 1108 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5449
timestamp 1712256841
transform 1 0 212 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5450
timestamp 1712256841
transform 1 0 140 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5451
timestamp 1712256841
transform 1 0 244 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5452
timestamp 1712256841
transform 1 0 140 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5453
timestamp 1712256841
transform 1 0 308 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5454
timestamp 1712256841
transform 1 0 220 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5455
timestamp 1712256841
transform 1 0 492 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5456
timestamp 1712256841
transform 1 0 404 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5457
timestamp 1712256841
transform 1 0 660 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5458
timestamp 1712256841
transform 1 0 580 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5459
timestamp 1712256841
transform 1 0 524 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5460
timestamp 1712256841
transform 1 0 420 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5461
timestamp 1712256841
transform 1 0 892 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5462
timestamp 1712256841
transform 1 0 788 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5463
timestamp 1712256841
transform 1 0 1044 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5464
timestamp 1712256841
transform 1 0 980 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5465
timestamp 1712256841
transform 1 0 3380 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5466
timestamp 1712256841
transform 1 0 3316 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5467
timestamp 1712256841
transform 1 0 3364 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1712256841
transform 1 0 3316 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5469
timestamp 1712256841
transform 1 0 3180 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5470
timestamp 1712256841
transform 1 0 3036 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5471
timestamp 1712256841
transform 1 0 3196 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5472
timestamp 1712256841
transform 1 0 3076 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5473
timestamp 1712256841
transform 1 0 3404 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5474
timestamp 1712256841
transform 1 0 3332 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5475
timestamp 1712256841
transform 1 0 3340 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5476
timestamp 1712256841
transform 1 0 3244 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5477
timestamp 1712256841
transform 1 0 3396 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_5478
timestamp 1712256841
transform 1 0 3348 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_5479
timestamp 1712256841
transform 1 0 3348 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_5480
timestamp 1712256841
transform 1 0 3332 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1712256841
transform 1 0 3364 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5482
timestamp 1712256841
transform 1 0 3324 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1712256841
transform 1 0 3404 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5484
timestamp 1712256841
transform 1 0 3364 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1712256841
transform 1 0 3340 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1712256841
transform 1 0 3308 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5487
timestamp 1712256841
transform 1 0 3308 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5488
timestamp 1712256841
transform 1 0 3252 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1712256841
transform 1 0 3244 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1712256841
transform 1 0 3244 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5491
timestamp 1712256841
transform 1 0 3212 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5492
timestamp 1712256841
transform 1 0 3212 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5493
timestamp 1712256841
transform 1 0 3132 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5494
timestamp 1712256841
transform 1 0 3132 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1712256841
transform 1 0 3116 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5496
timestamp 1712256841
transform 1 0 3116 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5497
timestamp 1712256841
transform 1 0 3068 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5498
timestamp 1712256841
transform 1 0 2940 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1712256841
transform 1 0 2884 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5500
timestamp 1712256841
transform 1 0 2364 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1712256841
transform 1 0 2340 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_5502
timestamp 1712256841
transform 1 0 2324 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5503
timestamp 1712256841
transform 1 0 2316 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1712256841
transform 1 0 2292 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5505
timestamp 1712256841
transform 1 0 2284 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_5506
timestamp 1712256841
transform 1 0 3052 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5507
timestamp 1712256841
transform 1 0 2716 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5508
timestamp 1712256841
transform 1 0 2556 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5509
timestamp 1712256841
transform 1 0 2372 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1712256841
transform 1 0 2212 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5511
timestamp 1712256841
transform 1 0 2116 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5512
timestamp 1712256841
transform 1 0 1812 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5513
timestamp 1712256841
transform 1 0 1636 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5514
timestamp 1712256841
transform 1 0 1428 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5515
timestamp 1712256841
transform 1 0 1060 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5516
timestamp 1712256841
transform 1 0 916 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5517
timestamp 1712256841
transform 1 0 2124 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5518
timestamp 1712256841
transform 1 0 1996 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5519
timestamp 1712256841
transform 1 0 2204 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5520
timestamp 1712256841
transform 1 0 2188 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5521
timestamp 1712256841
transform 1 0 2164 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5522
timestamp 1712256841
transform 1 0 2068 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5523
timestamp 1712256841
transform 1 0 1716 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5524
timestamp 1712256841
transform 1 0 2420 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5525
timestamp 1712256841
transform 1 0 2388 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5526
timestamp 1712256841
transform 1 0 2380 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5527
timestamp 1712256841
transform 1 0 1740 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5528
timestamp 1712256841
transform 1 0 2508 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5529
timestamp 1712256841
transform 1 0 2508 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5530
timestamp 1712256841
transform 1 0 2444 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5531
timestamp 1712256841
transform 1 0 2356 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5532
timestamp 1712256841
transform 1 0 2356 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5533
timestamp 1712256841
transform 1 0 2228 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5534
timestamp 1712256841
transform 1 0 2228 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5535
timestamp 1712256841
transform 1 0 1940 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5536
timestamp 1712256841
transform 1 0 2628 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5537
timestamp 1712256841
transform 1 0 2460 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5538
timestamp 1712256841
transform 1 0 2196 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5539
timestamp 1712256841
transform 1 0 1844 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5540
timestamp 1712256841
transform 1 0 2860 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5541
timestamp 1712256841
transform 1 0 2796 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5542
timestamp 1712256841
transform 1 0 2468 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5543
timestamp 1712256841
transform 1 0 1292 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1712256841
transform 1 0 1220 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5545
timestamp 1712256841
transform 1 0 1188 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5546
timestamp 1712256841
transform 1 0 1188 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5547
timestamp 1712256841
transform 1 0 1156 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5548
timestamp 1712256841
transform 1 0 1156 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5549
timestamp 1712256841
transform 1 0 1004 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5550
timestamp 1712256841
transform 1 0 972 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5551
timestamp 1712256841
transform 1 0 1044 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5552
timestamp 1712256841
transform 1 0 956 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5553
timestamp 1712256841
transform 1 0 844 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5554
timestamp 1712256841
transform 1 0 812 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5555
timestamp 1712256841
transform 1 0 812 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5556
timestamp 1712256841
transform 1 0 3020 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5557
timestamp 1712256841
transform 1 0 2980 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5558
timestamp 1712256841
transform 1 0 2932 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5559
timestamp 1712256841
transform 1 0 2900 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5560
timestamp 1712256841
transform 1 0 2852 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5561
timestamp 1712256841
transform 1 0 940 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5562
timestamp 1712256841
transform 1 0 852 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5563
timestamp 1712256841
transform 1 0 732 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5564
timestamp 1712256841
transform 1 0 692 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5565
timestamp 1712256841
transform 1 0 956 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5566
timestamp 1712256841
transform 1 0 900 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5567
timestamp 1712256841
transform 1 0 796 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5568
timestamp 1712256841
transform 1 0 772 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5569
timestamp 1712256841
transform 1 0 700 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5570
timestamp 1712256841
transform 1 0 628 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5571
timestamp 1712256841
transform 1 0 892 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5572
timestamp 1712256841
transform 1 0 660 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5573
timestamp 1712256841
transform 1 0 596 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5574
timestamp 1712256841
transform 1 0 596 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5575
timestamp 1712256841
transform 1 0 532 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5576
timestamp 1712256841
transform 1 0 508 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5577
timestamp 1712256841
transform 1 0 708 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5578
timestamp 1712256841
transform 1 0 524 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5579
timestamp 1712256841
transform 1 0 444 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5580
timestamp 1712256841
transform 1 0 444 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5581
timestamp 1712256841
transform 1 0 404 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5582
timestamp 1712256841
transform 1 0 404 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5583
timestamp 1712256841
transform 1 0 620 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5584
timestamp 1712256841
transform 1 0 516 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_5585
timestamp 1712256841
transform 1 0 380 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_5586
timestamp 1712256841
transform 1 0 356 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5587
timestamp 1712256841
transform 1 0 692 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5588
timestamp 1712256841
transform 1 0 596 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5589
timestamp 1712256841
transform 1 0 588 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5590
timestamp 1712256841
transform 1 0 564 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5591
timestamp 1712256841
transform 1 0 324 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_5592
timestamp 1712256841
transform 1 0 324 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5593
timestamp 1712256841
transform 1 0 308 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5594
timestamp 1712256841
transform 1 0 308 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5595
timestamp 1712256841
transform 1 0 244 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5596
timestamp 1712256841
transform 1 0 244 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_5597
timestamp 1712256841
transform 1 0 772 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5598
timestamp 1712256841
transform 1 0 772 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5599
timestamp 1712256841
transform 1 0 572 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5600
timestamp 1712256841
transform 1 0 428 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5601
timestamp 1712256841
transform 1 0 396 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5602
timestamp 1712256841
transform 1 0 340 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5603
timestamp 1712256841
transform 1 0 340 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_5604
timestamp 1712256841
transform 1 0 252 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5605
timestamp 1712256841
transform 1 0 244 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_5606
timestamp 1712256841
transform 1 0 228 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5607
timestamp 1712256841
transform 1 0 644 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5608
timestamp 1712256841
transform 1 0 636 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5609
timestamp 1712256841
transform 1 0 508 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5610
timestamp 1712256841
transform 1 0 508 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5611
timestamp 1712256841
transform 1 0 380 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5612
timestamp 1712256841
transform 1 0 380 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5613
timestamp 1712256841
transform 1 0 92 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5614
timestamp 1712256841
transform 1 0 68 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5615
timestamp 1712256841
transform 1 0 908 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5616
timestamp 1712256841
transform 1 0 732 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_5617
timestamp 1712256841
transform 1 0 572 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5618
timestamp 1712256841
transform 1 0 572 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5619
timestamp 1712256841
transform 1 0 300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5620
timestamp 1712256841
transform 1 0 300 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_5621
timestamp 1712256841
transform 1 0 172 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5622
timestamp 1712256841
transform 1 0 116 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5623
timestamp 1712256841
transform 1 0 916 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5624
timestamp 1712256841
transform 1 0 876 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5625
timestamp 1712256841
transform 1 0 876 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5626
timestamp 1712256841
transform 1 0 788 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5627
timestamp 1712256841
transform 1 0 756 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5628
timestamp 1712256841
transform 1 0 740 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5629
timestamp 1712256841
transform 1 0 652 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5630
timestamp 1712256841
transform 1 0 652 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5631
timestamp 1712256841
transform 1 0 652 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5632
timestamp 1712256841
transform 1 0 596 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5633
timestamp 1712256841
transform 1 0 564 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5634
timestamp 1712256841
transform 1 0 3044 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5635
timestamp 1712256841
transform 1 0 2876 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5636
timestamp 1712256841
transform 1 0 2868 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5637
timestamp 1712256841
transform 1 0 2868 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5638
timestamp 1712256841
transform 1 0 2820 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5639
timestamp 1712256841
transform 1 0 2724 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5640
timestamp 1712256841
transform 1 0 2468 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5641
timestamp 1712256841
transform 1 0 1412 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5642
timestamp 1712256841
transform 1 0 1052 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5643
timestamp 1712256841
transform 1 0 1044 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5644
timestamp 1712256841
transform 1 0 1036 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5645
timestamp 1712256841
transform 1 0 1036 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5646
timestamp 1712256841
transform 1 0 1020 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5647
timestamp 1712256841
transform 1 0 1012 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_5648
timestamp 1712256841
transform 1 0 1012 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5649
timestamp 1712256841
transform 1 0 988 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5650
timestamp 1712256841
transform 1 0 988 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5651
timestamp 1712256841
transform 1 0 980 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1712256841
transform 1 0 1700 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5653
timestamp 1712256841
transform 1 0 1692 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5654
timestamp 1712256841
transform 1 0 1668 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5655
timestamp 1712256841
transform 1 0 1644 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5656
timestamp 1712256841
transform 1 0 1636 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5657
timestamp 1712256841
transform 1 0 1636 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_5658
timestamp 1712256841
transform 1 0 1540 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5659
timestamp 1712256841
transform 1 0 1532 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1712256841
transform 1 0 1404 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5661
timestamp 1712256841
transform 1 0 1404 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5662
timestamp 1712256841
transform 1 0 1372 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5663
timestamp 1712256841
transform 1 0 1348 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5664
timestamp 1712256841
transform 1 0 1348 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5665
timestamp 1712256841
transform 1 0 1268 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5666
timestamp 1712256841
transform 1 0 1268 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5667
timestamp 1712256841
transform 1 0 1236 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5668
timestamp 1712256841
transform 1 0 1236 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5669
timestamp 1712256841
transform 1 0 1164 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5670
timestamp 1712256841
transform 1 0 1164 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5671
timestamp 1712256841
transform 1 0 1132 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5672
timestamp 1712256841
transform 1 0 1124 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5673
timestamp 1712256841
transform 1 0 1412 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5674
timestamp 1712256841
transform 1 0 1396 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5675
timestamp 1712256841
transform 1 0 1372 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5676
timestamp 1712256841
transform 1 0 1308 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5677
timestamp 1712256841
transform 1 0 1308 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5678
timestamp 1712256841
transform 1 0 1308 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5679
timestamp 1712256841
transform 1 0 1284 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5680
timestamp 1712256841
transform 1 0 1260 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5681
timestamp 1712256841
transform 1 0 1220 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5682
timestamp 1712256841
transform 1 0 1124 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5683
timestamp 1712256841
transform 1 0 1604 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5684
timestamp 1712256841
transform 1 0 1604 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5685
timestamp 1712256841
transform 1 0 1572 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5686
timestamp 1712256841
transform 1 0 1564 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5687
timestamp 1712256841
transform 1 0 1564 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5688
timestamp 1712256841
transform 1 0 1556 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1712256841
transform 1 0 1532 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5690
timestamp 1712256841
transform 1 0 1516 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5691
timestamp 1712256841
transform 1 0 1508 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1712256841
transform 1 0 1484 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1712256841
transform 1 0 1428 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1712256841
transform 1 0 1268 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5695
timestamp 1712256841
transform 1 0 1628 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5696
timestamp 1712256841
transform 1 0 1516 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5697
timestamp 1712256841
transform 1 0 1476 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5698
timestamp 1712256841
transform 1 0 1460 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5699
timestamp 1712256841
transform 1 0 1460 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5700
timestamp 1712256841
transform 1 0 1444 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5701
timestamp 1712256841
transform 1 0 1436 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5702
timestamp 1712256841
transform 1 0 1908 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1712256841
transform 1 0 1900 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5704
timestamp 1712256841
transform 1 0 1900 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5705
timestamp 1712256841
transform 1 0 1876 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5706
timestamp 1712256841
transform 1 0 1876 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5707
timestamp 1712256841
transform 1 0 1836 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1712256841
transform 1 0 2188 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5709
timestamp 1712256841
transform 1 0 2132 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5710
timestamp 1712256841
transform 1 0 2108 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1712256841
transform 1 0 2108 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5712
timestamp 1712256841
transform 1 0 2044 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5713
timestamp 1712256841
transform 1 0 2044 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1712256841
transform 1 0 2004 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5715
timestamp 1712256841
transform 1 0 2004 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1712256841
transform 1 0 2004 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_5717
timestamp 1712256841
transform 1 0 2292 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5718
timestamp 1712256841
transform 1 0 2292 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5719
timestamp 1712256841
transform 1 0 2292 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5720
timestamp 1712256841
transform 1 0 2252 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5721
timestamp 1712256841
transform 1 0 2252 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5722
timestamp 1712256841
transform 1 0 2244 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5723
timestamp 1712256841
transform 1 0 2236 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5724
timestamp 1712256841
transform 1 0 2236 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1712256841
transform 1 0 2220 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5726
timestamp 1712256841
transform 1 0 2212 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5727
timestamp 1712256841
transform 1 0 2180 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5728
timestamp 1712256841
transform 1 0 2172 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5729
timestamp 1712256841
transform 1 0 2812 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5730
timestamp 1712256841
transform 1 0 2756 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5731
timestamp 1712256841
transform 1 0 2756 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5732
timestamp 1712256841
transform 1 0 2708 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1712256841
transform 1 0 2708 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5734
timestamp 1712256841
transform 1 0 2532 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5735
timestamp 1712256841
transform 1 0 2436 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5736
timestamp 1712256841
transform 1 0 3268 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5737
timestamp 1712256841
transform 1 0 3140 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5738
timestamp 1712256841
transform 1 0 2428 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5739
timestamp 1712256841
transform 1 0 2332 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5740
timestamp 1712256841
transform 1 0 2460 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5741
timestamp 1712256841
transform 1 0 2308 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5742
timestamp 1712256841
transform 1 0 2812 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5743
timestamp 1712256841
transform 1 0 2772 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5744
timestamp 1712256841
transform 1 0 2500 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1712256841
transform 1 0 2500 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5746
timestamp 1712256841
transform 1 0 2388 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5747
timestamp 1712256841
transform 1 0 2252 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5748
timestamp 1712256841
transform 1 0 2444 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5749
timestamp 1712256841
transform 1 0 2380 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1712256841
transform 1 0 2164 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5751
timestamp 1712256841
transform 1 0 2572 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1712256841
transform 1 0 2460 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5753
timestamp 1712256841
transform 1 0 2412 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5754
timestamp 1712256841
transform 1 0 2532 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5755
timestamp 1712256841
transform 1 0 2372 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5756
timestamp 1712256841
transform 1 0 2628 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5757
timestamp 1712256841
transform 1 0 2412 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5758
timestamp 1712256841
transform 1 0 2284 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5759
timestamp 1712256841
transform 1 0 2212 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5760
timestamp 1712256841
transform 1 0 2428 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5761
timestamp 1712256841
transform 1 0 2204 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5762
timestamp 1712256841
transform 1 0 1948 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5763
timestamp 1712256841
transform 1 0 1828 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5764
timestamp 1712256841
transform 1 0 1628 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5765
timestamp 1712256841
transform 1 0 2340 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5766
timestamp 1712256841
transform 1 0 2308 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5767
timestamp 1712256841
transform 1 0 2284 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5768
timestamp 1712256841
transform 1 0 2284 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5769
timestamp 1712256841
transform 1 0 1940 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5770
timestamp 1712256841
transform 1 0 1596 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5771
timestamp 1712256841
transform 1 0 2276 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5772
timestamp 1712256841
transform 1 0 2276 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5773
timestamp 1712256841
transform 1 0 2236 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5774
timestamp 1712256841
transform 1 0 1724 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5775
timestamp 1712256841
transform 1 0 1596 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5776
timestamp 1712256841
transform 1 0 2068 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5777
timestamp 1712256841
transform 1 0 1724 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5778
timestamp 1712256841
transform 1 0 1524 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5779
timestamp 1712256841
transform 1 0 1820 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5780
timestamp 1712256841
transform 1 0 1788 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5781
timestamp 1712256841
transform 1 0 1788 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5782
timestamp 1712256841
transform 1 0 1660 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5783
timestamp 1712256841
transform 1 0 1468 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5784
timestamp 1712256841
transform 1 0 1204 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5785
timestamp 1712256841
transform 1 0 1876 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5786
timestamp 1712256841
transform 1 0 1764 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5787
timestamp 1712256841
transform 1 0 1620 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5788
timestamp 1712256841
transform 1 0 1500 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5789
timestamp 1712256841
transform 1 0 1500 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5790
timestamp 1712256841
transform 1 0 1100 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5791
timestamp 1712256841
transform 1 0 1740 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5792
timestamp 1712256841
transform 1 0 1700 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5793
timestamp 1712256841
transform 1 0 1684 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5794
timestamp 1712256841
transform 1 0 1628 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5795
timestamp 1712256841
transform 1 0 1492 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5796
timestamp 1712256841
transform 1 0 1220 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5797
timestamp 1712256841
transform 1 0 1684 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5798
timestamp 1712256841
transform 1 0 1612 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5799
timestamp 1712256841
transform 1 0 1556 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5800
timestamp 1712256841
transform 1 0 1500 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5801
timestamp 1712256841
transform 1 0 1484 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5802
timestamp 1712256841
transform 1 0 1116 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5803
timestamp 1712256841
transform 1 0 1460 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5804
timestamp 1712256841
transform 1 0 1292 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5805
timestamp 1712256841
transform 1 0 772 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5806
timestamp 1712256841
transform 1 0 1356 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5807
timestamp 1712256841
transform 1 0 1260 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5808
timestamp 1712256841
transform 1 0 692 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5809
timestamp 1712256841
transform 1 0 1324 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_5810
timestamp 1712256841
transform 1 0 1236 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_5811
timestamp 1712256841
transform 1 0 652 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_5812
timestamp 1712256841
transform 1 0 1252 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5813
timestamp 1712256841
transform 1 0 1212 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5814
timestamp 1712256841
transform 1 0 1212 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5815
timestamp 1712256841
transform 1 0 948 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5816
timestamp 1712256841
transform 1 0 724 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5817
timestamp 1712256841
transform 1 0 1252 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5818
timestamp 1712256841
transform 1 0 1140 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5819
timestamp 1712256841
transform 1 0 924 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5820
timestamp 1712256841
transform 1 0 820 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5821
timestamp 1712256841
transform 1 0 1020 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5822
timestamp 1712256841
transform 1 0 948 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5823
timestamp 1712256841
transform 1 0 788 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5824
timestamp 1712256841
transform 1 0 1156 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5825
timestamp 1712256841
transform 1 0 924 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5826
timestamp 1712256841
transform 1 0 924 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5827
timestamp 1712256841
transform 1 0 812 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1712256841
transform 1 0 652 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5829
timestamp 1712256841
transform 1 0 1020 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5830
timestamp 1712256841
transform 1 0 900 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5831
timestamp 1712256841
transform 1 0 788 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5832
timestamp 1712256841
transform 1 0 756 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5833
timestamp 1712256841
transform 1 0 796 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5834
timestamp 1712256841
transform 1 0 724 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5835
timestamp 1712256841
transform 1 0 692 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5836
timestamp 1712256841
transform 1 0 684 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5837
timestamp 1712256841
transform 1 0 676 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5838
timestamp 1712256841
transform 1 0 612 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5839
timestamp 1712256841
transform 1 0 724 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5840
timestamp 1712256841
transform 1 0 700 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5841
timestamp 1712256841
transform 1 0 636 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5842
timestamp 1712256841
transform 1 0 540 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5843
timestamp 1712256841
transform 1 0 796 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5844
timestamp 1712256841
transform 1 0 716 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5845
timestamp 1712256841
transform 1 0 596 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5846
timestamp 1712256841
transform 1 0 588 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5847
timestamp 1712256841
transform 1 0 564 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5848
timestamp 1712256841
transform 1 0 556 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5849
timestamp 1712256841
transform 1 0 548 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5850
timestamp 1712256841
transform 1 0 836 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5851
timestamp 1712256841
transform 1 0 708 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5852
timestamp 1712256841
transform 1 0 668 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5853
timestamp 1712256841
transform 1 0 660 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5854
timestamp 1712256841
transform 1 0 620 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5855
timestamp 1712256841
transform 1 0 612 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5856
timestamp 1712256841
transform 1 0 1012 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5857
timestamp 1712256841
transform 1 0 996 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5858
timestamp 1712256841
transform 1 0 932 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5859
timestamp 1712256841
transform 1 0 3388 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5860
timestamp 1712256841
transform 1 0 3364 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1712256841
transform 1 0 3292 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1712256841
transform 1 0 3268 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1712256841
transform 1 0 3156 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5864
timestamp 1712256841
transform 1 0 3116 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5865
timestamp 1712256841
transform 1 0 2924 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5866
timestamp 1712256841
transform 1 0 2820 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5867
timestamp 1712256841
transform 1 0 2716 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5868
timestamp 1712256841
transform 1 0 2596 0 1 2955
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1712256841
transform 1 0 3096 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1712256841
transform 1 0 2080 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1712256841
transform 1 0 1512 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1712256841
transform 1 0 1784 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1712256841
transform 1 0 2520 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1712256841
transform 1 0 560 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1712256841
transform 1 0 2408 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1712256841
transform 1 0 752 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1712256841
transform 1 0 1968 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1712256841
transform 1 0 1896 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1712256841
transform 1 0 112 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1712256841
transform 1 0 328 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1712256841
transform 1 0 2552 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1712256841
transform 1 0 2504 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1712256841
transform 1 0 2576 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1712256841
transform 1 0 1320 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1712256841
transform 1 0 1040 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1712256841
transform 1 0 1120 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1712256841
transform 1 0 1088 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1712256841
transform 1 0 992 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1712256841
transform 1 0 1344 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1712256841
transform 1 0 1240 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1712256841
transform 1 0 784 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1712256841
transform 1 0 784 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1712256841
transform 1 0 704 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1712256841
transform 1 0 512 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1712256841
transform 1 0 760 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1712256841
transform 1 0 480 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1712256841
transform 1 0 1064 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1712256841
transform 1 0 416 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1712256841
transform 1 0 512 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1712256841
transform 1 0 304 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1712256841
transform 1 0 528 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1712256841
transform 1 0 312 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1712256841
transform 1 0 1184 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1712256841
transform 1 0 296 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1712256841
transform 1 0 320 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1712256841
transform 1 0 144 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1712256841
transform 1 0 280 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1712256841
transform 1 0 104 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1712256841
transform 1 0 200 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1712256841
transform 1 0 1240 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1712256841
transform 1 0 392 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1712256841
transform 1 0 336 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1712256841
transform 1 0 200 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1712256841
transform 1 0 312 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1712256841
transform 1 0 920 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1712256841
transform 1 0 160 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1712256841
transform 1 0 176 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1712256841
transform 1 0 1072 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1712256841
transform 1 0 392 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1712256841
transform 1 0 208 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1712256841
transform 1 0 152 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1712256841
transform 1 0 184 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1712256841
transform 1 0 848 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1712256841
transform 1 0 1096 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1712256841
transform 1 0 448 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1712256841
transform 1 0 424 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1712256841
transform 1 0 128 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1712256841
transform 1 0 296 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1712256841
transform 1 0 160 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1712256841
transform 1 0 736 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1712256841
transform 1 0 1240 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1712256841
transform 1 0 400 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1712256841
transform 1 0 88 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1712256841
transform 1 0 200 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1712256841
transform 1 0 600 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1712256841
transform 1 0 1136 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1712256841
transform 1 0 320 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1712256841
transform 1 0 440 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1712256841
transform 1 0 96 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1712256841
transform 1 0 296 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1712256841
transform 1 0 624 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1712256841
transform 1 0 136 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1712256841
transform 1 0 136 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1712256841
transform 1 0 1216 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1712256841
transform 1 0 256 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1712256841
transform 1 0 368 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1712256841
transform 1 0 176 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1712256841
transform 1 0 256 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1712256841
transform 1 0 560 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1712256841
transform 1 0 112 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1712256841
transform 1 0 592 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1712256841
transform 1 0 520 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1712256841
transform 1 0 400 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1712256841
transform 1 0 464 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1712256841
transform 1 0 512 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1712256841
transform 1 0 568 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_88
timestamp 1712256841
transform 1 0 1096 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_89
timestamp 1712256841
transform 1 0 896 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1712256841
transform 1 0 912 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_91
timestamp 1712256841
transform 1 0 872 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_92
timestamp 1712256841
transform 1 0 880 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1712256841
transform 1 0 824 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_94
timestamp 1712256841
transform 1 0 792 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_95
timestamp 1712256841
transform 1 0 1216 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1712256841
transform 1 0 1112 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_97
timestamp 1712256841
transform 1 0 1032 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_98
timestamp 1712256841
transform 1 0 1184 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1712256841
transform 1 0 1072 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_100
timestamp 1712256841
transform 1 0 1160 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_101
timestamp 1712256841
transform 1 0 1072 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1712256841
transform 1 0 1032 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_103
timestamp 1712256841
transform 1 0 1440 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1712256841
transform 1 0 1512 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1712256841
transform 1 0 1424 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_106
timestamp 1712256841
transform 1 0 1216 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_107
timestamp 1712256841
transform 1 0 1056 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_108
timestamp 1712256841
transform 1 0 1824 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_109
timestamp 1712256841
transform 1 0 1760 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_110
timestamp 1712256841
transform 1 0 1784 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_111
timestamp 1712256841
transform 1 0 1680 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_112
timestamp 1712256841
transform 1 0 1712 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1712256841
transform 1 0 1656 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_114
timestamp 1712256841
transform 1 0 1584 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_115
timestamp 1712256841
transform 1 0 1240 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_116
timestamp 1712256841
transform 1 0 2080 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_117
timestamp 1712256841
transform 1 0 2088 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1712256841
transform 1 0 2200 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_119
timestamp 1712256841
transform 1 0 2136 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_120
timestamp 1712256841
transform 1 0 1968 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1712256841
transform 1 0 1928 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_122
timestamp 1712256841
transform 1 0 2384 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1712256841
transform 1 0 2376 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1712256841
transform 1 0 2272 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1712256841
transform 1 0 2408 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_126
timestamp 1712256841
transform 1 0 2168 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_127
timestamp 1712256841
transform 1 0 2120 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_128
timestamp 1712256841
transform 1 0 2072 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_129
timestamp 1712256841
transform 1 0 1296 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_130
timestamp 1712256841
transform 1 0 2448 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_131
timestamp 1712256841
transform 1 0 2568 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_132
timestamp 1712256841
transform 1 0 2288 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_133
timestamp 1712256841
transform 1 0 2496 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_134
timestamp 1712256841
transform 1 0 2168 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_135
timestamp 1712256841
transform 1 0 2128 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_136
timestamp 1712256841
transform 1 0 2456 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_137
timestamp 1712256841
transform 1 0 2512 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_138
timestamp 1712256841
transform 1 0 2328 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_139
timestamp 1712256841
transform 1 0 2136 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_140
timestamp 1712256841
transform 1 0 2280 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_141
timestamp 1712256841
transform 1 0 2032 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_142
timestamp 1712256841
transform 1 0 2120 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_143
timestamp 1712256841
transform 1 0 2512 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_144
timestamp 1712256841
transform 1 0 2488 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_145
timestamp 1712256841
transform 1 0 2520 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_146
timestamp 1712256841
transform 1 0 2200 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_147
timestamp 1712256841
transform 1 0 2272 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_148
timestamp 1712256841
transform 1 0 2008 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_149
timestamp 1712256841
transform 1 0 2072 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_150
timestamp 1712256841
transform 1 0 1768 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_151
timestamp 1712256841
transform 1 0 1736 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_152
timestamp 1712256841
transform 1 0 1808 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_153
timestamp 1712256841
transform 1 0 1760 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_154
timestamp 1712256841
transform 1 0 1840 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_155
timestamp 1712256841
transform 1 0 1800 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_156
timestamp 1712256841
transform 1 0 1816 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_157
timestamp 1712256841
transform 1 0 1352 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_158
timestamp 1712256841
transform 1 0 2280 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_159
timestamp 1712256841
transform 1 0 1952 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_160
timestamp 1712256841
transform 1 0 1928 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_161
timestamp 1712256841
transform 1 0 1880 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_162
timestamp 1712256841
transform 1 0 1928 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_163
timestamp 1712256841
transform 1 0 1880 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_164
timestamp 1712256841
transform 1 0 1832 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_165
timestamp 1712256841
transform 1 0 2024 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_166
timestamp 1712256841
transform 1 0 2248 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_167
timestamp 1712256841
transform 1 0 2200 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_168
timestamp 1712256841
transform 1 0 2144 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_169
timestamp 1712256841
transform 1 0 2240 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_170
timestamp 1712256841
transform 1 0 2120 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_171
timestamp 1712256841
transform 1 0 2152 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_172
timestamp 1712256841
transform 1 0 2312 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_173
timestamp 1712256841
transform 1 0 2448 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_174
timestamp 1712256841
transform 1 0 2352 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_175
timestamp 1712256841
transform 1 0 2416 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_176
timestamp 1712256841
transform 1 0 2368 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_177
timestamp 1712256841
transform 1 0 2408 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_178
timestamp 1712256841
transform 1 0 2360 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_179
timestamp 1712256841
transform 1 0 2272 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_180
timestamp 1712256841
transform 1 0 2624 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_181
timestamp 1712256841
transform 1 0 2576 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_182
timestamp 1712256841
transform 1 0 2520 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_183
timestamp 1712256841
transform 1 0 2648 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_184
timestamp 1712256841
transform 1 0 2080 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_185
timestamp 1712256841
transform 1 0 2024 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_186
timestamp 1712256841
transform 1 0 2520 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_187
timestamp 1712256841
transform 1 0 2616 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_188
timestamp 1712256841
transform 1 0 2560 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_189
timestamp 1712256841
transform 1 0 2816 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_190
timestamp 1712256841
transform 1 0 2600 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_191
timestamp 1712256841
transform 1 0 2536 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_192
timestamp 1712256841
transform 1 0 2712 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_193
timestamp 1712256841
transform 1 0 2504 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_194
timestamp 1712256841
transform 1 0 2520 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_195
timestamp 1712256841
transform 1 0 2816 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_196
timestamp 1712256841
transform 1 0 2496 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_197
timestamp 1712256841
transform 1 0 3152 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_198
timestamp 1712256841
transform 1 0 2720 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_199
timestamp 1712256841
transform 1 0 2872 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_200
timestamp 1712256841
transform 1 0 3056 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_201
timestamp 1712256841
transform 1 0 3224 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_202
timestamp 1712256841
transform 1 0 3352 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_203
timestamp 1712256841
transform 1 0 3328 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_204
timestamp 1712256841
transform 1 0 3272 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_205
timestamp 1712256841
transform 1 0 2976 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_206
timestamp 1712256841
transform 1 0 3048 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_207
timestamp 1712256841
transform 1 0 2952 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_208
timestamp 1712256841
transform 1 0 3072 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_209
timestamp 1712256841
transform 1 0 3040 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_210
timestamp 1712256841
transform 1 0 2456 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_211
timestamp 1712256841
transform 1 0 2504 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_212
timestamp 1712256841
transform 1 0 2888 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_213
timestamp 1712256841
transform 1 0 992 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_214
timestamp 1712256841
transform 1 0 1416 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_215
timestamp 1712256841
transform 1 0 1576 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_216
timestamp 1712256841
transform 1 0 1912 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_217
timestamp 1712256841
transform 1 0 3160 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_218
timestamp 1712256841
transform 1 0 2320 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_219
timestamp 1712256841
transform 1 0 1320 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_220
timestamp 1712256841
transform 1 0 3256 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_221
timestamp 1712256841
transform 1 0 3264 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_222
timestamp 1712256841
transform 1 0 3232 0 -1 2370
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1712256841
transform 1 0 2680 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1712256841
transform 1 0 1448 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1712256841
transform 1 0 1496 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1712256841
transform 1 0 832 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1712256841
transform 1 0 224 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1712256841
transform 1 0 1536 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1712256841
transform 1 0 448 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1712256841
transform 1 0 504 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1712256841
transform 1 0 880 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1712256841
transform 1 0 1568 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1712256841
transform 1 0 736 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1712256841
transform 1 0 1936 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1712256841
transform 1 0 1664 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1712256841
transform 1 0 1592 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1712256841
transform 1 0 1408 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1712256841
transform 1 0 344 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1712256841
transform 1 0 1352 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1712256841
transform 1 0 1960 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1712256841
transform 1 0 1384 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1712256841
transform 1 0 1768 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1712256841
transform 1 0 136 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1712256841
transform 1 0 1760 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1712256841
transform 1 0 1080 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1712256841
transform 1 0 824 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1712256841
transform 1 0 456 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1712256841
transform 1 0 624 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1712256841
transform 1 0 336 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1712256841
transform 1 0 488 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1712256841
transform 1 0 288 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1712256841
transform 1 0 600 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1712256841
transform 1 0 232 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1712256841
transform 1 0 368 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1712256841
transform 1 0 504 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1712256841
transform 1 0 960 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1712256841
transform 1 0 248 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1712256841
transform 1 0 320 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1712256841
transform 1 0 640 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1712256841
transform 1 0 720 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1712256841
transform 1 0 272 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1712256841
transform 1 0 744 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1712256841
transform 1 0 816 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1712256841
transform 1 0 296 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1712256841
transform 1 0 576 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1712256841
transform 1 0 640 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1712256841
transform 1 0 320 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1712256841
transform 1 0 680 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1712256841
transform 1 0 840 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1712256841
transform 1 0 288 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_48
timestamp 1712256841
transform 1 0 568 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_49
timestamp 1712256841
transform 1 0 672 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_50
timestamp 1712256841
transform 1 0 224 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_51
timestamp 1712256841
transform 1 0 696 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_52
timestamp 1712256841
transform 1 0 824 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_53
timestamp 1712256841
transform 1 0 496 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_54
timestamp 1712256841
transform 1 0 664 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1712256841
transform 1 0 904 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_56
timestamp 1712256841
transform 1 0 280 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_57
timestamp 1712256841
transform 1 0 304 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_58
timestamp 1712256841
transform 1 0 752 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_59
timestamp 1712256841
transform 1 0 216 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_60
timestamp 1712256841
transform 1 0 1088 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_61
timestamp 1712256841
transform 1 0 408 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_62
timestamp 1712256841
transform 1 0 696 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_63
timestamp 1712256841
transform 1 0 352 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_64
timestamp 1712256841
transform 1 0 912 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_65
timestamp 1712256841
transform 1 0 944 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_66
timestamp 1712256841
transform 1 0 976 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_67
timestamp 1712256841
transform 1 0 1040 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_68
timestamp 1712256841
transform 1 0 1032 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_69
timestamp 1712256841
transform 1 0 1080 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_70
timestamp 1712256841
transform 1 0 1176 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_71
timestamp 1712256841
transform 1 0 1232 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_72
timestamp 1712256841
transform 1 0 1520 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_73
timestamp 1712256841
transform 1 0 1488 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_74
timestamp 1712256841
transform 1 0 1384 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_75
timestamp 1712256841
transform 1 0 1296 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_76
timestamp 1712256841
transform 1 0 1384 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_77
timestamp 1712256841
transform 1 0 1648 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_78
timestamp 1712256841
transform 1 0 1752 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_79
timestamp 1712256841
transform 1 0 1760 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_80
timestamp 1712256841
transform 1 0 1704 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_81
timestamp 1712256841
transform 1 0 1616 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_82
timestamp 1712256841
transform 1 0 1744 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_83
timestamp 1712256841
transform 1 0 2184 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_84
timestamp 1712256841
transform 1 0 1872 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_85
timestamp 1712256841
transform 1 0 1872 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_86
timestamp 1712256841
transform 1 0 2248 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_87
timestamp 1712256841
transform 1 0 1960 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_88
timestamp 1712256841
transform 1 0 1888 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_89
timestamp 1712256841
transform 1 0 2432 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_90
timestamp 1712256841
transform 1 0 2016 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_91
timestamp 1712256841
transform 1 0 1912 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_92
timestamp 1712256841
transform 1 0 2368 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_93
timestamp 1712256841
transform 1 0 2400 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_94
timestamp 1712256841
transform 1 0 2080 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_95
timestamp 1712256841
transform 1 0 2336 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_96
timestamp 1712256841
transform 1 0 1408 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_97
timestamp 1712256841
transform 1 0 1512 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_98
timestamp 1712256841
transform 1 0 2232 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_99
timestamp 1712256841
transform 1 0 2072 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_100
timestamp 1712256841
transform 1 0 2232 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_101
timestamp 1712256841
transform 1 0 2184 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_102
timestamp 1712256841
transform 1 0 1968 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_103
timestamp 1712256841
transform 1 0 2120 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_104
timestamp 1712256841
transform 1 0 1760 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_105
timestamp 1712256841
transform 1 0 1712 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_106
timestamp 1712256841
transform 1 0 1904 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_107
timestamp 1712256841
transform 1 0 1880 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_108
timestamp 1712256841
transform 1 0 1920 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_109
timestamp 1712256841
transform 1 0 2152 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_110
timestamp 1712256841
transform 1 0 2288 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_111
timestamp 1712256841
transform 1 0 1976 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_112
timestamp 1712256841
transform 1 0 2096 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_113
timestamp 1712256841
transform 1 0 2192 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_114
timestamp 1712256841
transform 1 0 2208 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_115
timestamp 1712256841
transform 1 0 2224 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_116
timestamp 1712256841
transform 1 0 2408 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_117
timestamp 1712256841
transform 1 0 2264 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_118
timestamp 1712256841
transform 1 0 2352 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_119
timestamp 1712256841
transform 1 0 2440 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_120
timestamp 1712256841
transform 1 0 2400 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_121
timestamp 1712256841
transform 1 0 2448 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_122
timestamp 1712256841
transform 1 0 2648 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_123
timestamp 1712256841
transform 1 0 2456 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_124
timestamp 1712256841
transform 1 0 2528 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_125
timestamp 1712256841
transform 1 0 2664 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_126
timestamp 1712256841
transform 1 0 2528 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_127
timestamp 1712256841
transform 1 0 2664 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_128
timestamp 1712256841
transform 1 0 1968 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_129
timestamp 1712256841
transform 1 0 1960 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_130
timestamp 1712256841
transform 1 0 1352 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_131
timestamp 1712256841
transform 1 0 2600 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_132
timestamp 1712256841
transform 1 0 2960 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_133
timestamp 1712256841
transform 1 0 2960 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_134
timestamp 1712256841
transform 1 0 2752 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_135
timestamp 1712256841
transform 1 0 1768 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_136
timestamp 1712256841
transform 1 0 2800 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_137
timestamp 1712256841
transform 1 0 2592 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_138
timestamp 1712256841
transform 1 0 2904 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_139
timestamp 1712256841
transform 1 0 3056 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_140
timestamp 1712256841
transform 1 0 3072 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_141
timestamp 1712256841
transform 1 0 2584 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_142
timestamp 1712256841
transform 1 0 1832 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_143
timestamp 1712256841
transform 1 0 2744 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_144
timestamp 1712256841
transform 1 0 2688 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_145
timestamp 1712256841
transform 1 0 2952 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_146
timestamp 1712256841
transform 1 0 2888 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_147
timestamp 1712256841
transform 1 0 2808 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_148
timestamp 1712256841
transform 1 0 2704 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_149
timestamp 1712256841
transform 1 0 2824 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_150
timestamp 1712256841
transform 1 0 2656 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_151
timestamp 1712256841
transform 1 0 2560 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_152
timestamp 1712256841
transform 1 0 2848 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_153
timestamp 1712256841
transform 1 0 2760 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_154
timestamp 1712256841
transform 1 0 2624 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_155
timestamp 1712256841
transform 1 0 2880 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_156
timestamp 1712256841
transform 1 0 3176 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_157
timestamp 1712256841
transform 1 0 3384 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_158
timestamp 1712256841
transform 1 0 3392 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_159
timestamp 1712256841
transform 1 0 3248 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_160
timestamp 1712256841
transform 1 0 3184 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_161
timestamp 1712256841
transform 1 0 3384 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_162
timestamp 1712256841
transform 1 0 3384 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_163
timestamp 1712256841
transform 1 0 3320 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_164
timestamp 1712256841
transform 1 0 2880 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_165
timestamp 1712256841
transform 1 0 960 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_166
timestamp 1712256841
transform 1 0 1632 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_167
timestamp 1712256841
transform 1 0 1840 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_168
timestamp 1712256841
transform 1 0 1960 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_169
timestamp 1712256841
transform 1 0 3024 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_170
timestamp 1712256841
transform 1 0 3136 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_171
timestamp 1712256841
transform 1 0 3072 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_172
timestamp 1712256841
transform 1 0 3184 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_173
timestamp 1712256841
transform 1 0 2376 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_174
timestamp 1712256841
transform 1 0 1912 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_175
timestamp 1712256841
transform 1 0 704 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_176
timestamp 1712256841
transform 1 0 928 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_177
timestamp 1712256841
transform 1 0 912 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_178
timestamp 1712256841
transform 1 0 1936 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_179
timestamp 1712256841
transform 1 0 1224 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_180
timestamp 1712256841
transform 1 0 1480 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_181
timestamp 1712256841
transform 1 0 2200 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_182
timestamp 1712256841
transform 1 0 3120 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_183
timestamp 1712256841
transform 1 0 3352 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_184
timestamp 1712256841
transform 1 0 3384 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_185
timestamp 1712256841
transform 1 0 3024 0 1 2570
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1712256841
transform 1 0 2840 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1712256841
transform 1 0 3200 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1712256841
transform 1 0 848 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1712256841
transform 1 0 848 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1712256841
transform 1 0 2120 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1712256841
transform 1 0 1480 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1712256841
transform 1 0 584 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1712256841
transform 1 0 656 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1712256841
transform 1 0 1640 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1712256841
transform 1 0 1824 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1712256841
transform 1 0 872 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1712256841
transform 1 0 1704 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1712256841
transform 1 0 776 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1712256841
transform 1 0 696 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1712256841
transform 1 0 1880 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1712256841
transform 1 0 2456 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1712256841
transform 1 0 2072 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1712256841
transform 1 0 1552 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1712256841
transform 1 0 1856 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1712256841
transform 1 0 1568 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1712256841
transform 1 0 1656 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1712256841
transform 1 0 648 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1712256841
transform 1 0 152 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1712256841
transform 1 0 352 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1712256841
transform 1 0 1456 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1712256841
transform 1 0 1832 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1712256841
transform 1 0 88 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1712256841
transform 1 0 1856 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1712256841
transform 1 0 1512 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1712256841
transform 1 0 1536 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1712256841
transform 1 0 1360 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1712256841
transform 1 0 1320 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1712256841
transform 1 0 1344 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1712256841
transform 1 0 3144 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1712256841
transform 1 0 1312 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1712256841
transform 1 0 1128 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1712256841
transform 1 0 1624 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1712256841
transform 1 0 1352 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1712256841
transform 1 0 1144 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1712256841
transform 1 0 1144 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1712256841
transform 1 0 1256 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1712256841
transform 1 0 816 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1712256841
transform 1 0 904 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1712256841
transform 1 0 664 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1712256841
transform 1 0 992 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1712256841
transform 1 0 1200 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1712256841
transform 1 0 608 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1712256841
transform 1 0 872 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1712256841
transform 1 0 1296 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1712256841
transform 1 0 504 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1712256841
transform 1 0 128 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1712256841
transform 1 0 904 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1712256841
transform 1 0 1296 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1712256841
transform 1 0 944 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1712256841
transform 1 0 160 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1712256841
transform 1 0 880 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1712256841
transform 1 0 1064 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1712256841
transform 1 0 920 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1712256841
transform 1 0 880 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1712256841
transform 1 0 1072 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1712256841
transform 1 0 1296 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1712256841
transform 1 0 1016 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1712256841
transform 1 0 848 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1712256841
transform 1 0 992 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1712256841
transform 1 0 1120 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1712256841
transform 1 0 1296 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1712256841
transform 1 0 872 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1712256841
transform 1 0 2776 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1712256841
transform 1 0 744 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1712256841
transform 1 0 952 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1712256841
transform 1 0 656 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1712256841
transform 1 0 984 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1712256841
transform 1 0 544 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1712256841
transform 1 0 1056 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1712256841
transform 1 0 1208 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1712256841
transform 1 0 496 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1712256841
transform 1 0 1360 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1712256841
transform 1 0 1312 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1712256841
transform 1 0 1496 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1712256841
transform 1 0 1272 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1712256841
transform 1 0 280 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1712256841
transform 1 0 1752 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1712256841
transform 1 0 1352 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1712256841
transform 1 0 808 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1712256841
transform 1 0 2000 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1712256841
transform 1 0 1856 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1712256841
transform 1 0 1256 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1712256841
transform 1 0 560 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1712256841
transform 1 0 1736 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1712256841
transform 1 0 1344 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1712256841
transform 1 0 1720 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1712256841
transform 1 0 608 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1712256841
transform 1 0 1608 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1712256841
transform 1 0 1392 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1712256841
transform 1 0 1696 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1712256841
transform 1 0 1384 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1712256841
transform 1 0 1248 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1712256841
transform 1 0 560 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1712256841
transform 1 0 2776 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1712256841
transform 1 0 1896 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1712256841
transform 1 0 1832 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1712256841
transform 1 0 1192 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1712256841
transform 1 0 736 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1712256841
transform 1 0 1968 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1712256841
transform 1 0 1480 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1712256841
transform 1 0 856 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1712256841
transform 1 0 1920 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1712256841
transform 1 0 1712 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1712256841
transform 1 0 1648 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1712256841
transform 1 0 1400 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1712256841
transform 1 0 2456 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1712256841
transform 1 0 1864 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1712256841
transform 1 0 1544 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1712256841
transform 1 0 2464 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1712256841
transform 1 0 2224 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1712256841
transform 1 0 1784 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1712256841
transform 1 0 2720 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1712256841
transform 1 0 2408 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1712256841
transform 1 0 2064 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1712256841
transform 1 0 2624 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1712256841
transform 1 0 2344 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1712256841
transform 1 0 2472 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1712256841
transform 1 0 2568 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1712256841
transform 1 0 2720 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1712256841
transform 1 0 2752 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1712256841
transform 1 0 2504 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_126
timestamp 1712256841
transform 1 0 1504 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_127
timestamp 1712256841
transform 1 0 2992 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_128
timestamp 1712256841
transform 1 0 2664 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_129
timestamp 1712256841
transform 1 0 2776 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_130
timestamp 1712256841
transform 1 0 2800 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_131
timestamp 1712256841
transform 1 0 2920 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_132
timestamp 1712256841
transform 1 0 3112 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_133
timestamp 1712256841
transform 1 0 3032 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_134
timestamp 1712256841
transform 1 0 2672 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_135
timestamp 1712256841
transform 1 0 2768 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_136
timestamp 1712256841
transform 1 0 2752 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_137
timestamp 1712256841
transform 1 0 3136 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_138
timestamp 1712256841
transform 1 0 2952 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_139
timestamp 1712256841
transform 1 0 2848 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_140
timestamp 1712256841
transform 1 0 2752 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_141
timestamp 1712256841
transform 1 0 3288 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_142
timestamp 1712256841
transform 1 0 3264 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_143
timestamp 1712256841
transform 1 0 2752 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_144
timestamp 1712256841
transform 1 0 2672 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_145
timestamp 1712256841
transform 1 0 3176 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_146
timestamp 1712256841
transform 1 0 3240 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_147
timestamp 1712256841
transform 1 0 3288 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_148
timestamp 1712256841
transform 1 0 2040 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_149
timestamp 1712256841
transform 1 0 2720 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_150
timestamp 1712256841
transform 1 0 2744 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_151
timestamp 1712256841
transform 1 0 2728 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_152
timestamp 1712256841
transform 1 0 2824 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_153
timestamp 1712256841
transform 1 0 2712 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_154
timestamp 1712256841
transform 1 0 3128 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_155
timestamp 1712256841
transform 1 0 3320 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_156
timestamp 1712256841
transform 1 0 3056 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_157
timestamp 1712256841
transform 1 0 3280 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_158
timestamp 1712256841
transform 1 0 3272 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_159
timestamp 1712256841
transform 1 0 3352 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_160
timestamp 1712256841
transform 1 0 3344 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_161
timestamp 1712256841
transform 1 0 3248 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_162
timestamp 1712256841
transform 1 0 2792 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_163
timestamp 1712256841
transform 1 0 2512 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_164
timestamp 1712256841
transform 1 0 2448 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_165
timestamp 1712256841
transform 1 0 752 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_166
timestamp 1712256841
transform 1 0 784 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_167
timestamp 1712256841
transform 1 0 840 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_168
timestamp 1712256841
transform 1 0 1640 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_169
timestamp 1712256841
transform 1 0 1816 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_170
timestamp 1712256841
transform 1 0 1888 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_171
timestamp 1712256841
transform 1 0 1096 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_172
timestamp 1712256841
transform 1 0 848 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_173
timestamp 1712256841
transform 1 0 536 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_174
timestamp 1712256841
transform 1 0 616 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_175
timestamp 1712256841
transform 1 0 464 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_176
timestamp 1712256841
transform 1 0 416 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_177
timestamp 1712256841
transform 1 0 440 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_178
timestamp 1712256841
transform 1 0 304 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_179
timestamp 1712256841
transform 1 0 192 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_180
timestamp 1712256841
transform 1 0 136 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_181
timestamp 1712256841
transform 1 0 160 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_182
timestamp 1712256841
transform 1 0 1064 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_183
timestamp 1712256841
transform 1 0 1168 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_184
timestamp 1712256841
transform 1 0 1232 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_185
timestamp 1712256841
transform 1 0 1432 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_186
timestamp 1712256841
transform 1 0 1456 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_187
timestamp 1712256841
transform 1 0 1520 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_188
timestamp 1712256841
transform 1 0 1720 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_189
timestamp 1712256841
transform 1 0 1880 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_190
timestamp 1712256841
transform 1 0 1824 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_191
timestamp 1712256841
transform 1 0 2024 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_192
timestamp 1712256841
transform 1 0 2048 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_193
timestamp 1712256841
transform 1 0 2216 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_194
timestamp 1712256841
transform 1 0 1952 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_195
timestamp 1712256841
transform 1 0 2376 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_196
timestamp 1712256841
transform 1 0 2608 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_197
timestamp 1712256841
transform 1 0 2648 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_198
timestamp 1712256841
transform 1 0 2576 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_199
timestamp 1712256841
transform 1 0 2808 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_200
timestamp 1712256841
transform 1 0 2992 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_201
timestamp 1712256841
transform 1 0 2704 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_202
timestamp 1712256841
transform 1 0 3168 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_203
timestamp 1712256841
transform 1 0 2432 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_204
timestamp 1712256841
transform 1 0 920 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_205
timestamp 1712256841
transform 1 0 888 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_206
timestamp 1712256841
transform 1 0 1736 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_207
timestamp 1712256841
transform 1 0 2168 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_208
timestamp 1712256841
transform 1 0 1264 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_209
timestamp 1712256841
transform 1 0 2208 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_210
timestamp 1712256841
transform 1 0 3328 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_211
timestamp 1712256841
transform 1 0 3288 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_212
timestamp 1712256841
transform 1 0 3384 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_213
timestamp 1712256841
transform 1 0 3272 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_214
timestamp 1712256841
transform 1 0 3264 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_215
timestamp 1712256841
transform 1 0 3400 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_216
timestamp 1712256841
transform 1 0 3344 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_217
timestamp 1712256841
transform 1 0 3256 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_218
timestamp 1712256841
transform 1 0 3328 0 1 770
box -8 -3 32 105
use NOR3X1  NOR3X1_0
timestamp 1712256841
transform 1 0 3176 0 -1 1970
box -7 -3 68 105
use OAI21X1  OAI21X1_0
timestamp 1712256841
transform 1 0 3128 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1712256841
transform 1 0 1576 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1712256841
transform 1 0 2176 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1712256841
transform 1 0 1080 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1712256841
transform 1 0 1672 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1712256841
transform 1 0 1832 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1712256841
transform 1 0 1504 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1712256841
transform 1 0 1528 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1712256841
transform 1 0 1696 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1712256841
transform 1 0 1416 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1712256841
transform 1 0 880 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1712256841
transform 1 0 1408 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1712256841
transform 1 0 2584 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1712256841
transform 1 0 2656 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1712256841
transform 1 0 1240 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1712256841
transform 1 0 2000 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1712256841
transform 1 0 1632 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1712256841
transform 1 0 2144 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1712256841
transform 1 0 256 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1712256841
transform 1 0 640 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1712256841
transform 1 0 96 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1712256841
transform 1 0 1664 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1712256841
transform 1 0 296 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1712256841
transform 1 0 1424 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1712256841
transform 1 0 1336 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1712256841
transform 1 0 1944 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1712256841
transform 1 0 1688 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1712256841
transform 1 0 88 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1712256841
transform 1 0 656 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1712256841
transform 1 0 1208 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1712256841
transform 1 0 1872 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1712256841
transform 1 0 2080 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1712256841
transform 1 0 1312 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1712256841
transform 1 0 1536 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1712256841
transform 1 0 1432 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1712256841
transform 1 0 1584 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1712256841
transform 1 0 1280 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1712256841
transform 1 0 1256 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1712256841
transform 1 0 1200 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1712256841
transform 1 0 1064 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1712256841
transform 1 0 1240 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1712256841
transform 1 0 1200 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1712256841
transform 1 0 1344 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1712256841
transform 1 0 1152 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1712256841
transform 1 0 1008 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1712256841
transform 1 0 824 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1712256841
transform 1 0 768 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1712256841
transform 1 0 1080 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1712256841
transform 1 0 1128 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1712256841
transform 1 0 1312 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1712256841
transform 1 0 1160 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1712256841
transform 1 0 1072 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1712256841
transform 1 0 896 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1712256841
transform 1 0 696 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1712256841
transform 1 0 992 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1712256841
transform 1 0 1184 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1712256841
transform 1 0 1320 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1712256841
transform 1 0 952 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1712256841
transform 1 0 1384 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1712256841
transform 1 0 1448 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1712256841
transform 1 0 464 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1712256841
transform 1 0 528 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1712256841
transform 1 0 1192 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1712256841
transform 1 0 872 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1712256841
transform 1 0 1096 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1712256841
transform 1 0 888 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1712256841
transform 1 0 1192 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1712256841
transform 1 0 392 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1712256841
transform 1 0 360 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1712256841
transform 1 0 776 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1712256841
transform 1 0 680 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1712256841
transform 1 0 648 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1712256841
transform 1 0 712 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1712256841
transform 1 0 336 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1712256841
transform 1 0 232 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1712256841
transform 1 0 968 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1712256841
transform 1 0 712 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1712256841
transform 1 0 816 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1712256841
transform 1 0 608 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1712256841
transform 1 0 256 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1712256841
transform 1 0 216 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1712256841
transform 1 0 1064 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1712256841
transform 1 0 672 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1712256841
transform 1 0 1128 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1712256841
transform 1 0 216 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1712256841
transform 1 0 208 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1712256841
transform 1 0 712 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1712256841
transform 1 0 816 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1712256841
transform 1 0 784 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1712256841
transform 1 0 88 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1712256841
transform 1 0 96 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1712256841
transform 1 0 592 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1712256841
transform 1 0 752 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1712256841
transform 1 0 648 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1712256841
transform 1 0 152 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1712256841
transform 1 0 88 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1712256841
transform 1 0 632 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1712256841
transform 1 0 760 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1712256841
transform 1 0 744 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1712256841
transform 1 0 592 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1712256841
transform 1 0 224 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1712256841
transform 1 0 936 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1712256841
transform 1 0 856 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1712256841
transform 1 0 968 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1712256841
transform 1 0 1000 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1712256841
transform 1 0 224 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1712256841
transform 1 0 872 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1712256841
transform 1 0 760 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1712256841
transform 1 0 976 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1712256841
transform 1 0 1032 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1712256841
transform 1 0 1160 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1712256841
transform 1 0 1120 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1712256841
transform 1 0 616 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1712256841
transform 1 0 768 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1712256841
transform 1 0 664 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1712256841
transform 1 0 608 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1712256841
transform 1 0 1176 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1712256841
transform 1 0 1360 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1712256841
transform 1 0 864 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1712256841
transform 1 0 952 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1712256841
transform 1 0 880 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1712256841
transform 1 0 824 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1712256841
transform 1 0 1224 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1712256841
transform 1 0 1416 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1712256841
transform 1 0 1168 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1712256841
transform 1 0 1184 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1712256841
transform 1 0 1464 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1712256841
transform 1 0 1128 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1712256841
transform 1 0 1464 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1712256841
transform 1 0 1496 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1712256841
transform 1 0 1344 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1712256841
transform 1 0 1320 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1712256841
transform 1 0 1440 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1712256841
transform 1 0 1672 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1712256841
transform 1 0 1768 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1712256841
transform 1 0 1600 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1712256841
transform 1 0 1680 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1712256841
transform 1 0 1632 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1712256841
transform 1 0 1800 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1712256841
transform 1 0 2032 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1712256841
transform 1 0 2016 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1712256841
transform 1 0 1960 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1712256841
transform 1 0 1800 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1712256841
transform 1 0 1864 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1712256841
transform 1 0 2296 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1712256841
transform 1 0 1768 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1712256841
transform 1 0 1888 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1712256841
transform 1 0 1656 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1712256841
transform 1 0 2112 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1712256841
transform 1 0 2288 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1712256841
transform 1 0 1616 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1712256841
transform 1 0 2488 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1712256841
transform 1 0 1544 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1712256841
transform 1 0 2016 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1712256841
transform 1 0 1472 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1712256841
transform 1 0 1528 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1712256841
transform 1 0 2240 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1712256841
transform 1 0 2248 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1712256841
transform 1 0 1920 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1712256841
transform 1 0 2304 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1712256841
transform 1 0 1976 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1712256841
transform 1 0 2256 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1712256841
transform 1 0 1336 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_163
timestamp 1712256841
transform 1 0 2296 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_164
timestamp 1712256841
transform 1 0 2328 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_165
timestamp 1712256841
transform 1 0 1952 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_166
timestamp 1712256841
transform 1 0 2328 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_167
timestamp 1712256841
transform 1 0 2056 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_168
timestamp 1712256841
transform 1 0 2320 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_169
timestamp 1712256841
transform 1 0 1704 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_170
timestamp 1712256841
transform 1 0 1544 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_171
timestamp 1712256841
transform 1 0 1984 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_172
timestamp 1712256841
transform 1 0 1824 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_173
timestamp 1712256841
transform 1 0 1752 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_174
timestamp 1712256841
transform 1 0 2032 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_175
timestamp 1712256841
transform 1 0 1704 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_176
timestamp 1712256841
transform 1 0 2056 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_177
timestamp 1712256841
transform 1 0 1928 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_178
timestamp 1712256841
transform 1 0 2040 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_179
timestamp 1712256841
transform 1 0 2200 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_180
timestamp 1712256841
transform 1 0 2064 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_181
timestamp 1712256841
transform 1 0 2416 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_182
timestamp 1712256841
transform 1 0 2176 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_183
timestamp 1712256841
transform 1 0 2304 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_184
timestamp 1712256841
transform 1 0 2344 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_185
timestamp 1712256841
transform 1 0 2416 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_186
timestamp 1712256841
transform 1 0 2480 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_187
timestamp 1712256841
transform 1 0 2360 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_188
timestamp 1712256841
transform 1 0 2560 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_189
timestamp 1712256841
transform 1 0 2576 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_190
timestamp 1712256841
transform 1 0 2496 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_191
timestamp 1712256841
transform 1 0 2600 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_192
timestamp 1712256841
transform 1 0 2536 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_193
timestamp 1712256841
transform 1 0 2680 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_194
timestamp 1712256841
transform 1 0 2648 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_195
timestamp 1712256841
transform 1 0 2648 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_196
timestamp 1712256841
transform 1 0 2816 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_197
timestamp 1712256841
transform 1 0 2896 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_198
timestamp 1712256841
transform 1 0 2968 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_199
timestamp 1712256841
transform 1 0 2992 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_200
timestamp 1712256841
transform 1 0 3008 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_201
timestamp 1712256841
transform 1 0 3008 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_202
timestamp 1712256841
transform 1 0 2888 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_203
timestamp 1712256841
transform 1 0 2856 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_204
timestamp 1712256841
transform 1 0 2920 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_205
timestamp 1712256841
transform 1 0 2968 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_206
timestamp 1712256841
transform 1 0 3040 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_207
timestamp 1712256841
transform 1 0 3072 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_208
timestamp 1712256841
transform 1 0 3128 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_209
timestamp 1712256841
transform 1 0 3080 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_210
timestamp 1712256841
transform 1 0 3032 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_211
timestamp 1712256841
transform 1 0 3136 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_212
timestamp 1712256841
transform 1 0 3008 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_213
timestamp 1712256841
transform 1 0 2848 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_214
timestamp 1712256841
transform 1 0 2864 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_215
timestamp 1712256841
transform 1 0 2856 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_216
timestamp 1712256841
transform 1 0 3008 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_217
timestamp 1712256841
transform 1 0 3008 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_218
timestamp 1712256841
transform 1 0 2968 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_219
timestamp 1712256841
transform 1 0 2840 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_220
timestamp 1712256841
transform 1 0 2832 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_221
timestamp 1712256841
transform 1 0 3032 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_222
timestamp 1712256841
transform 1 0 2808 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_223
timestamp 1712256841
transform 1 0 2696 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_224
timestamp 1712256841
transform 1 0 2744 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_225
timestamp 1712256841
transform 1 0 2704 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_226
timestamp 1712256841
transform 1 0 2856 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_227
timestamp 1712256841
transform 1 0 2872 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_228
timestamp 1712256841
transform 1 0 2600 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_229
timestamp 1712256841
transform 1 0 2760 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_230
timestamp 1712256841
transform 1 0 2664 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_231
timestamp 1712256841
transform 1 0 2744 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_232
timestamp 1712256841
transform 1 0 2800 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_233
timestamp 1712256841
transform 1 0 3168 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_234
timestamp 1712256841
transform 1 0 3216 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_235
timestamp 1712256841
transform 1 0 3328 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_236
timestamp 1712256841
transform 1 0 3280 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_237
timestamp 1712256841
transform 1 0 2744 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_238
timestamp 1712256841
transform 1 0 2896 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_239
timestamp 1712256841
transform 1 0 3080 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_240
timestamp 1712256841
transform 1 0 3168 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_241
timestamp 1712256841
transform 1 0 3320 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_242
timestamp 1712256841
transform 1 0 3368 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_243
timestamp 1712256841
transform 1 0 3336 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_244
timestamp 1712256841
transform 1 0 2936 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_245
timestamp 1712256841
transform 1 0 3016 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_246
timestamp 1712256841
transform 1 0 3096 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_247
timestamp 1712256841
transform 1 0 3248 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_248
timestamp 1712256841
transform 1 0 3392 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_249
timestamp 1712256841
transform 1 0 3160 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_250
timestamp 1712256841
transform 1 0 3128 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_251
timestamp 1712256841
transform 1 0 3240 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_252
timestamp 1712256841
transform 1 0 3016 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_253
timestamp 1712256841
transform 1 0 2944 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_254
timestamp 1712256841
transform 1 0 2848 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_255
timestamp 1712256841
transform 1 0 2712 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_256
timestamp 1712256841
transform 1 0 2400 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_257
timestamp 1712256841
transform 1 0 2152 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_258
timestamp 1712256841
transform 1 0 1992 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_259
timestamp 1712256841
transform 1 0 2080 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_260
timestamp 1712256841
transform 1 0 3120 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_261
timestamp 1712256841
transform 1 0 2944 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_262
timestamp 1712256841
transform 1 0 2512 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_263
timestamp 1712256841
transform 1 0 2528 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_264
timestamp 1712256841
transform 1 0 2592 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_265
timestamp 1712256841
transform 1 0 2384 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_266
timestamp 1712256841
transform 1 0 2456 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_267
timestamp 1712256841
transform 1 0 2184 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_268
timestamp 1712256841
transform 1 0 1976 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_269
timestamp 1712256841
transform 1 0 2120 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_270
timestamp 1712256841
transform 1 0 2208 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_271
timestamp 1712256841
transform 1 0 2296 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_272
timestamp 1712256841
transform 1 0 2152 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_273
timestamp 1712256841
transform 1 0 2232 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_274
timestamp 1712256841
transform 1 0 2040 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_275
timestamp 1712256841
transform 1 0 2096 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_276
timestamp 1712256841
transform 1 0 1992 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_277
timestamp 1712256841
transform 1 0 1936 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_278
timestamp 1712256841
transform 1 0 1760 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_279
timestamp 1712256841
transform 1 0 1832 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_280
timestamp 1712256841
transform 1 0 1888 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_281
timestamp 1712256841
transform 1 0 1928 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_282
timestamp 1712256841
transform 1 0 1632 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_283
timestamp 1712256841
transform 1 0 1728 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_284
timestamp 1712256841
transform 1 0 1536 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_285
timestamp 1712256841
transform 1 0 1704 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_286
timestamp 1712256841
transform 1 0 1432 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_287
timestamp 1712256841
transform 1 0 1520 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_288
timestamp 1712256841
transform 1 0 1392 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_289
timestamp 1712256841
transform 1 0 1392 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_290
timestamp 1712256841
transform 1 0 1280 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_291
timestamp 1712256841
transform 1 0 1376 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_292
timestamp 1712256841
transform 1 0 1224 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_293
timestamp 1712256841
transform 1 0 1408 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_294
timestamp 1712256841
transform 1 0 1520 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_295
timestamp 1712256841
transform 1 0 1472 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_296
timestamp 1712256841
transform 1 0 1168 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_297
timestamp 1712256841
transform 1 0 1208 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_298
timestamp 1712256841
transform 1 0 192 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_299
timestamp 1712256841
transform 1 0 1104 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_300
timestamp 1712256841
transform 1 0 224 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_301
timestamp 1712256841
transform 1 0 1112 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_302
timestamp 1712256841
transform 1 0 280 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_303
timestamp 1712256841
transform 1 0 984 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_304
timestamp 1712256841
transform 1 0 1064 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_305
timestamp 1712256841
transform 1 0 1112 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_306
timestamp 1712256841
transform 1 0 272 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_307
timestamp 1712256841
transform 1 0 600 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_308
timestamp 1712256841
transform 1 0 464 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_309
timestamp 1712256841
transform 1 0 568 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_310
timestamp 1712256841
transform 1 0 344 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_311
timestamp 1712256841
transform 1 0 528 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_312
timestamp 1712256841
transform 1 0 432 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_313
timestamp 1712256841
transform 1 0 560 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_314
timestamp 1712256841
transform 1 0 640 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_315
timestamp 1712256841
transform 1 0 808 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_316
timestamp 1712256841
transform 1 0 496 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_317
timestamp 1712256841
transform 1 0 688 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_318
timestamp 1712256841
transform 1 0 864 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_319
timestamp 1712256841
transform 1 0 832 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_320
timestamp 1712256841
transform 1 0 1016 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_321
timestamp 1712256841
transform 1 0 968 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_322
timestamp 1712256841
transform 1 0 3080 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_323
timestamp 1712256841
transform 1 0 2864 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_324
timestamp 1712256841
transform 1 0 3384 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_325
timestamp 1712256841
transform 1 0 3376 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_326
timestamp 1712256841
transform 1 0 3168 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_327
timestamp 1712256841
transform 1 0 3240 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_328
timestamp 1712256841
transform 1 0 3160 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_329
timestamp 1712256841
transform 1 0 3312 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_330
timestamp 1712256841
transform 1 0 3360 0 -1 2370
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1712256841
transform 1 0 1568 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1712256841
transform 1 0 744 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1712256841
transform 1 0 2064 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1712256841
transform 1 0 1432 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1712256841
transform 1 0 1160 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1712256841
transform 1 0 968 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1712256841
transform 1 0 968 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1712256841
transform 1 0 952 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1712256841
transform 1 0 1136 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1712256841
transform 1 0 1064 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1712256841
transform 1 0 1160 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1712256841
transform 1 0 1272 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1712256841
transform 1 0 1352 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1712256841
transform 1 0 1544 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1712256841
transform 1 0 2032 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1712256841
transform 1 0 1584 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1712256841
transform 1 0 1448 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1712256841
transform 1 0 1848 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1712256841
transform 1 0 1424 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1712256841
transform 1 0 2120 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1712256841
transform 1 0 2384 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1712256841
transform 1 0 2504 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1712256841
transform 1 0 2552 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1712256841
transform 1 0 2600 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1712256841
transform 1 0 2920 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1712256841
transform 1 0 2896 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1712256841
transform 1 0 1152 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1712256841
transform 1 0 3064 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1712256841
transform 1 0 2912 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1712256841
transform 1 0 1256 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1712256841
transform 1 0 3040 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1712256841
transform 1 0 2832 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1712256841
transform 1 0 1544 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1712256841
transform 1 0 2904 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1712256841
transform 1 0 3264 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1712256841
transform 1 0 3280 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_36
timestamp 1712256841
transform 1 0 2832 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_37
timestamp 1712256841
transform 1 0 2984 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_38
timestamp 1712256841
transform 1 0 3040 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1712256841
transform 1 0 3368 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_40
timestamp 1712256841
transform 1 0 3272 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_41
timestamp 1712256841
transform 1 0 3288 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1712256841
transform 1 0 3176 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_43
timestamp 1712256841
transform 1 0 1280 0 1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_44
timestamp 1712256841
transform 1 0 2728 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_45
timestamp 1712256841
transform 1 0 2832 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_46
timestamp 1712256841
transform 1 0 2688 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_47
timestamp 1712256841
transform 1 0 2744 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_48
timestamp 1712256841
transform 1 0 3224 0 1 2570
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1712256841
transform 1 0 3368 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1712256841
transform 1 0 3280 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1712256841
transform 1 0 3224 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1712256841
transform 1 0 2864 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1712256841
transform 1 0 3200 0 1 1970
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1712256841
transform 1 0 3080 0 -1 2970
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1712256841
transform 1 0 3192 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1712256841
transform 1 0 3304 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_8
timestamp 1712256841
transform 1 0 3168 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_9
timestamp 1712256841
transform 1 0 1648 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_10
timestamp 1712256841
transform 1 0 1224 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_11
timestamp 1712256841
transform 1 0 936 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_12
timestamp 1712256841
transform 1 0 888 0 1 1970
box -8 -3 40 105
use OR2X1  OR2X1_13
timestamp 1712256841
transform 1 0 1288 0 1 1770
box -8 -3 40 105
use OR2X1  OR2X1_14
timestamp 1712256841
transform 1 0 448 0 -1 1570
box -8 -3 40 105
use OR2X1  OR2X1_15
timestamp 1712256841
transform 1 0 496 0 1 1570
box -8 -3 40 105
use OR2X1  OR2X1_16
timestamp 1712256841
transform 1 0 448 0 -1 970
box -8 -3 40 105
use OR2X1  OR2X1_17
timestamp 1712256841
transform 1 0 504 0 1 970
box -8 -3 40 105
use OR2X1  OR2X1_18
timestamp 1712256841
transform 1 0 1328 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_19
timestamp 1712256841
transform 1 0 2640 0 -1 1370
box -8 -3 40 105
use OR2X1  OR2X1_20
timestamp 1712256841
transform 1 0 3128 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_21
timestamp 1712256841
transform 1 0 3064 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_22
timestamp 1712256841
transform 1 0 3240 0 -1 970
box -8 -3 40 105
use OR2X2  OR2X2_0
timestamp 1712256841
transform 1 0 3360 0 1 770
box -7 -3 35 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1712256841
transform 1 0 3480 0 1 3317
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1712256841
transform 1 0 3480 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1712256841
transform 1 0 24 0 1 3317
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1712256841
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1712256841
transform 1 0 3456 0 1 3293
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1712256841
transform 1 0 3456 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1712256841
transform 1 0 48 0 1 3293
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1712256841
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1712256841
transform 1 0 3480 0 1 3270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1712256841
transform 1 0 3480 0 1 3070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1712256841
transform 1 0 3480 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1712256841
transform 1 0 3480 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1712256841
transform 1 0 3480 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1712256841
transform 1 0 3480 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1712256841
transform 1 0 3480 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1712256841
transform 1 0 3480 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1712256841
transform 1 0 3480 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1712256841
transform 1 0 3480 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1712256841
transform 1 0 3480 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1712256841
transform 1 0 3480 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1712256841
transform 1 0 3480 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1712256841
transform 1 0 3480 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1712256841
transform 1 0 3480 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1712256841
transform 1 0 3480 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1712256841
transform 1 0 3480 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1712256841
transform 1 0 24 0 1 3270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1712256841
transform 1 0 24 0 1 3070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1712256841
transform 1 0 24 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1712256841
transform 1 0 24 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1712256841
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1712256841
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1712256841
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1712256841
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1712256841
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1712256841
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1712256841
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1712256841
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1712256841
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1712256841
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1712256841
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1712256841
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1712256841
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1712256841
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1712256841
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1712256841
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1712256841
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1712256841
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1712256841
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1712256841
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1712256841
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1712256841
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1712256841
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1712256841
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1712256841
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1712256841
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1712256841
transform 1 0 48 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1712256841
transform 1 0 48 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1712256841
transform 1 0 48 0 1 3170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_50
timestamp 1712256841
transform 1 0 3456 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_51
timestamp 1712256841
transform 1 0 3456 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_52
timestamp 1712256841
transform 1 0 3456 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_53
timestamp 1712256841
transform 1 0 3456 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_54
timestamp 1712256841
transform 1 0 3456 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_55
timestamp 1712256841
transform 1 0 3456 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_56
timestamp 1712256841
transform 1 0 3456 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_57
timestamp 1712256841
transform 1 0 3456 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_58
timestamp 1712256841
transform 1 0 3456 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_59
timestamp 1712256841
transform 1 0 3456 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_60
timestamp 1712256841
transform 1 0 3456 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_61
timestamp 1712256841
transform 1 0 3456 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_62
timestamp 1712256841
transform 1 0 3456 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_63
timestamp 1712256841
transform 1 0 3456 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_64
timestamp 1712256841
transform 1 0 3456 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_65
timestamp 1712256841
transform 1 0 3456 0 1 3170
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1712256841
transform 1 0 3016 0 -1 770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1712256841
transform 1 0 3264 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1712256841
transform 1 0 3376 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_3
timestamp 1712256841
transform 1 0 3096 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_4
timestamp 1712256841
transform 1 0 2824 0 1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_5
timestamp 1712256841
transform 1 0 2976 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1712256841
transform 1 0 2784 0 -1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1712256841
transform 1 0 2840 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1712256841
transform 1 0 2752 0 -1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_3
timestamp 1712256841
transform 1 0 2936 0 -1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1712256841
transform 1 0 3040 0 1 3170
box -8 -3 64 105
<< labels >>
rlabel electrodecontact s 3180 3135 3180 3135 4 in_clka
rlabel metal1 2164 2615 2164 2615 4 in_clkb
rlabel electrodecontact s 3340 2015 3340 2015 4 in_restart
rlabel electrodecontact s 3292 805 3292 805 4 in_move[1]
rlabel electrodecontact s 3396 805 3396 805 4 in_move[0]
rlabel metal1 1020 2925 1020 2925 4 board_out[31]
rlabel metal1 964 2815 964 2815 4 board_out[30]
rlabel metal1 684 2815 684 2815 4 board_out[29]
rlabel metal1 788 2815 788 2815 4 board_out[28]
rlabel metal1 684 2725 684 2725 4 board_out[27]
rlabel metal1 548 2615 548 2615 4 board_out[26]
rlabel electrodecontact s 540 2925 540 2925 4 board_out[25]
rlabel metal1 572 2725 572 2725 4 board_out[24]
rlabel electrodecontact s 788 3125 788 3125 4 board_out[23]
rlabel metal1 660 3125 660 3125 4 board_out[22]
rlabel metal1 940 3015 940 3015 4 board_out[21]
rlabel electrodecontact s 924 3015 924 3015 4 board_out[20]
rlabel metal1 980 3125 980 3125 4 board_out[19]
rlabel metal1 1276 3125 1276 3125 4 board_out[18]
rlabel electrodecontact s 1268 2925 1268 2925 4 board_out[17]
rlabel metal1 1316 3015 1316 3015 4 board_out[16]
rlabel metal1 1516 2725 1516 2725 4 board_out[15]
rlabel electrodecontact s 1740 2525 1740 2525 4 board_out[14]
rlabel metal1 1796 2725 1796 2725 4 board_out[13]
rlabel metal1 1860 2925 1860 2925 4 board_out[12]
rlabel metal1 2076 3125 2076 3125 4 board_out[11]
rlabel metal1 2260 2925 2260 2925 4 board_out[10]
rlabel electrodecontact s 2340 2925 2340 2925 4 board_out[9]
rlabel metal1 2004 3015 2004 3015 4 board_out[8]
rlabel metal1 2196 2925 2196 2925 4 board_out[7]
rlabel electrodecontact s 2420 3015 2420 3015 4 board_out[6]
rlabel metal1 2372 3125 2372 3125 4 board_out[5]
rlabel metal1 2476 3015 2476 3015 4 board_out[4]
rlabel metal1 2452 3015 2452 3015 4 board_out[3]
rlabel metal1 2860 3125 2860 3125 4 board_out[2]
rlabel metal1 2452 3215 2452 3215 4 board_out[1]
rlabel metal1 2436 3015 2436 3015 4 board_out[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 29340.002 6435.000 29425.502 6435.000 
<< end >>
