magic
tech scmos
timestamp 1711307567
<< metal1 >>
rect 14 2607 2818 2627
rect 38 2583 2794 2603
rect 38 2567 2794 2573
rect 994 2543 1028 2546
rect 346 2533 380 2536
rect 394 2533 412 2536
rect 418 2533 460 2536
rect 498 2533 508 2536
rect 602 2533 620 2536
rect 754 2533 780 2536
rect 834 2533 860 2536
rect 884 2533 908 2536
rect 922 2533 964 2536
rect 970 2533 988 2536
rect 994 2533 1036 2536
rect 1050 2533 1060 2536
rect 1066 2533 1100 2536
rect 1140 2533 1148 2536
rect 1228 2533 1245 2536
rect 1306 2533 1316 2536
rect 1330 2533 1340 2536
rect 322 2523 340 2526
rect 418 2525 421 2533
rect 658 2526 661 2533
rect 538 2523 556 2526
rect 596 2523 605 2526
rect 658 2523 700 2526
rect 714 2523 717 2533
rect 1354 2526 1357 2545
rect 1538 2543 1556 2546
rect 1746 2543 1756 2546
rect 1770 2543 1780 2546
rect 1532 2533 1549 2536
rect 1554 2533 1564 2536
rect 1676 2533 1701 2536
rect 1706 2533 1724 2536
rect 1738 2533 1764 2536
rect 1770 2533 1788 2536
rect 1890 2533 1908 2536
rect 1970 2533 1980 2536
rect 1994 2533 2012 2536
rect 2026 2533 2044 2536
rect 2098 2533 2108 2536
rect 2602 2533 2612 2536
rect 762 2523 788 2526
rect 828 2523 861 2526
rect 972 2523 981 2526
rect 1146 2523 1156 2526
rect 1290 2523 1324 2526
rect 1330 2523 1357 2526
rect 1378 2523 1412 2526
rect 1452 2523 1469 2526
rect 1506 2523 1516 2526
rect 1578 2523 1596 2526
rect 1642 2523 1660 2526
rect 1684 2523 1709 2526
rect 1770 2525 1773 2533
rect 1890 2523 1916 2526
rect 1922 2523 1932 2526
rect 1954 2523 1964 2526
rect 748 2513 773 2516
rect 1330 2515 1333 2523
rect 1466 2516 1469 2523
rect 1642 2516 1645 2523
rect 1466 2513 1477 2516
rect 1532 2513 1549 2516
rect 1628 2513 1645 2516
rect 1970 2515 1973 2533
rect 1978 2523 1988 2526
rect 1994 2523 2020 2526
rect 1996 2513 2013 2516
rect 2026 2515 2029 2533
rect 2674 2526 2677 2533
rect 2034 2523 2052 2526
rect 2058 2523 2076 2526
rect 2082 2523 2092 2526
rect 2236 2523 2261 2526
rect 2332 2523 2349 2526
rect 2428 2523 2453 2526
rect 2522 2523 2540 2526
rect 2596 2523 2613 2526
rect 2642 2523 2677 2526
rect 1818 2503 1844 2506
rect 2034 2503 2037 2523
rect 1818 2483 1821 2503
rect 14 2467 2818 2473
rect 1306 2426 1309 2456
rect 1850 2433 1876 2436
rect 1914 2433 1940 2436
rect 1962 2433 1980 2436
rect 1994 2433 2044 2436
rect 236 2423 253 2426
rect 316 2423 325 2426
rect 980 2423 997 2426
rect 1162 2416 1165 2426
rect 1300 2423 1309 2426
rect 1404 2423 1421 2426
rect 1468 2423 1477 2426
rect 1890 2423 1924 2426
rect 1994 2423 2028 2426
rect 2524 2423 2541 2426
rect 194 2413 220 2416
rect 282 2413 308 2416
rect 346 2406 349 2414
rect 354 2413 396 2416
rect 468 2413 485 2416
rect 492 2413 517 2416
rect 602 2413 652 2416
rect 682 2413 708 2416
rect 746 2413 756 2416
rect 762 2413 772 2416
rect 866 2413 964 2416
rect 978 2413 1044 2416
rect 1092 2413 1141 2416
rect 1162 2413 1188 2416
rect 1258 2413 1292 2416
rect 1348 2413 1381 2416
rect 1434 2413 1452 2416
rect 1474 2413 1516 2416
rect 1586 2413 1612 2416
rect 1628 2413 1661 2416
rect 1684 2413 1709 2416
rect 2058 2413 2068 2416
rect 2156 2413 2181 2416
rect 2388 2413 2413 2416
rect 2444 2413 2453 2416
rect 2492 2413 2508 2416
rect 2684 2413 2709 2416
rect 242 2403 268 2406
rect 282 2403 300 2406
rect 314 2403 340 2406
rect 346 2403 365 2406
rect 426 2403 460 2406
rect 482 2405 485 2413
rect 570 2403 580 2406
rect 602 2405 605 2413
rect 610 2403 644 2406
rect 668 2403 693 2406
rect 730 2403 748 2406
rect 778 2403 844 2406
rect 866 2405 869 2413
rect 980 2403 1029 2406
rect 1084 2403 1093 2406
rect 1106 2403 1148 2406
rect 1154 2403 1180 2406
rect 1194 2403 1228 2406
rect 1306 2403 1324 2406
rect 1354 2403 1380 2406
rect 1404 2403 1413 2406
rect 1468 2403 1485 2406
rect 1538 2403 1548 2406
rect 1578 2403 1604 2406
rect 1642 2403 1676 2406
rect 1690 2403 1724 2406
rect 2082 2403 2124 2406
rect 2458 2403 2484 2406
rect 2530 2403 2556 2406
rect 2604 2403 2620 2406
rect 2634 2403 2660 2406
rect 2698 2403 2708 2406
rect 322 2393 332 2396
rect 1050 2393 1076 2396
rect 1698 2393 1716 2396
rect 38 2367 2794 2373
rect 746 2353 781 2356
rect 578 2343 588 2346
rect 812 2343 837 2346
rect 930 2343 964 2346
rect 1242 2343 1276 2346
rect 178 2333 252 2336
rect 258 2333 341 2336
rect 346 2326 349 2334
rect 386 2326 389 2334
rect 412 2333 461 2336
rect 522 2333 548 2336
rect 596 2333 645 2336
rect 650 2326 653 2334
rect 666 2333 708 2336
rect 746 2333 796 2336
rect 852 2333 877 2336
rect 1026 2333 1036 2336
rect 1082 2333 1124 2336
rect 1236 2333 1261 2336
rect 1364 2333 1397 2336
rect 1426 2326 1429 2345
rect 1530 2343 1564 2346
rect 1482 2333 1492 2336
rect 1546 2333 1572 2336
rect 1586 2333 1596 2336
rect 1658 2326 1661 2345
rect 1690 2333 1724 2336
rect 1754 2333 1772 2336
rect 1796 2333 1805 2336
rect 1818 2333 1828 2336
rect 1956 2333 1965 2336
rect 2034 2333 2068 2336
rect 1754 2326 1757 2333
rect 116 2323 141 2326
rect 172 2323 205 2326
rect 260 2323 277 2326
rect 322 2323 349 2326
rect 356 2323 389 2326
rect 500 2323 549 2326
rect 604 2323 621 2326
rect 626 2323 653 2326
rect 660 2323 709 2326
rect 762 2323 788 2326
rect 812 2323 845 2326
rect 1074 2323 1132 2326
rect 1154 2323 1212 2326
rect 1300 2323 1325 2326
rect 1330 2323 1340 2326
rect 1420 2323 1429 2326
rect 1450 2323 1500 2326
rect 1506 2323 1516 2326
rect 1652 2323 1661 2326
rect 1748 2323 1757 2326
rect 1858 2323 1868 2326
rect 1898 2323 1932 2326
rect 2042 2323 2076 2326
rect 2114 2325 2117 2356
rect 2194 2343 2204 2346
rect 2180 2333 2205 2336
rect 2212 2333 2277 2336
rect 2394 2333 2404 2336
rect 2546 2333 2564 2336
rect 2618 2333 2644 2336
rect 2668 2333 2701 2336
rect 2484 2323 2509 2326
rect 2612 2323 2629 2326
rect 2634 2323 2652 2326
rect 2698 2325 2701 2333
rect 2732 2323 2741 2326
rect 2634 2316 2637 2323
rect 668 2313 685 2316
rect 924 2313 941 2316
rect 1796 2313 1829 2316
rect 2004 2313 2013 2316
rect 2588 2313 2597 2316
rect 2620 2313 2637 2316
rect 2002 2303 2020 2306
rect 14 2267 2818 2273
rect 212 2223 237 2226
rect 356 2223 365 2226
rect 1418 2223 1444 2226
rect 1468 2223 1477 2226
rect 1610 2223 1629 2226
rect 1828 2223 1845 2226
rect 146 2207 149 2216
rect 226 2213 252 2216
rect 274 2213 292 2216
rect 354 2213 380 2216
rect 484 2213 533 2216
rect 626 2206 629 2214
rect 674 2213 700 2216
rect 730 2213 764 2216
rect 780 2213 805 2216
rect 836 2213 845 2216
rect 908 2213 917 2216
rect 922 2213 964 2216
rect 970 2213 980 2216
rect 1052 2213 1085 2216
rect 1314 2213 1324 2216
rect 1330 2213 1397 2216
rect 1404 2213 1421 2216
rect 1508 2213 1533 2216
rect 1580 2213 1613 2216
rect 922 2206 925 2213
rect 1394 2207 1397 2213
rect 1626 2207 1629 2223
rect 2626 2216 2629 2226
rect 1642 2213 1660 2216
rect 1666 2213 1700 2216
rect 1826 2213 1860 2216
rect 1866 2213 1876 2216
rect 2012 2213 2029 2216
rect 2268 2213 2293 2216
rect 2396 2213 2413 2216
rect 2508 2213 2533 2216
rect 2594 2213 2629 2216
rect 268 2203 277 2206
rect 356 2203 373 2206
rect 378 2203 388 2206
rect 404 2203 413 2206
rect 434 2203 452 2206
rect 522 2203 532 2206
rect 564 2203 605 2206
rect 626 2203 644 2206
rect 650 2203 692 2206
rect 786 2203 820 2206
rect 834 2203 892 2206
rect 906 2203 925 2206
rect 986 2203 1044 2206
rect 1050 2203 1100 2206
rect 1148 2203 1204 2206
rect 1236 2203 1245 2206
rect 1250 2203 1309 2206
rect 1738 2203 1748 2206
rect 1834 2203 1852 2206
rect 1882 2203 1908 2206
rect 1946 2203 1980 2206
rect 1994 2203 2052 2206
rect 2116 2203 2157 2206
rect 2164 2203 2181 2206
rect 836 2193 861 2196
rect 908 2193 949 2196
rect 1130 2193 1140 2196
rect 1724 2193 1741 2196
rect 1986 2193 1996 2196
rect 2090 2193 2108 2196
rect 2122 2193 2156 2196
rect 2170 2193 2180 2196
rect 38 2167 2794 2173
rect 186 2136 189 2146
rect 300 2143 333 2146
rect 666 2143 684 2146
rect 330 2136 333 2143
rect 122 2133 132 2136
rect 186 2133 196 2136
rect 210 2133 220 2136
rect 330 2133 341 2136
rect 692 2133 709 2136
rect 714 2133 741 2136
rect 754 2133 773 2136
rect 802 2133 836 2136
rect 210 2126 213 2133
rect 754 2126 757 2133
rect 914 2126 917 2145
rect 1132 2143 1157 2146
rect 1330 2143 1372 2146
rect 1394 2143 1404 2146
rect 1394 2136 1397 2143
rect 924 2133 933 2136
rect 938 2133 956 2136
rect 1052 2133 1109 2136
rect 1130 2133 1164 2136
rect 1178 2133 1212 2136
rect 1380 2133 1397 2136
rect 1412 2133 1445 2136
rect 1290 2126 1293 2133
rect 1482 2126 1485 2156
rect 1930 2143 1956 2146
rect 2580 2143 2597 2146
rect 2594 2136 2597 2143
rect 1546 2133 1556 2136
rect 1578 2133 1628 2136
rect 1666 2133 1692 2136
rect 1780 2133 1812 2136
rect 1924 2133 1949 2136
rect 1970 2133 1989 2136
rect 2066 2133 2084 2136
rect 2116 2133 2133 2136
rect 2196 2133 2228 2136
rect 2252 2133 2269 2136
rect 2466 2133 2476 2136
rect 2498 2133 2564 2136
rect 2594 2133 2612 2136
rect 2618 2133 2628 2136
rect 2642 2133 2668 2136
rect 204 2123 213 2126
rect 228 2123 261 2126
rect 300 2123 309 2126
rect 314 2123 340 2126
rect 372 2123 389 2126
rect 450 2123 485 2126
rect 524 2123 548 2126
rect 644 2123 653 2126
rect 740 2123 757 2126
rect 762 2123 772 2126
rect 844 2123 861 2126
rect 876 2123 917 2126
rect 932 2123 949 2126
rect 1018 2123 1028 2126
rect 1060 2123 1085 2126
rect 1132 2123 1141 2126
rect 1172 2123 1220 2126
rect 1234 2123 1293 2126
rect 1426 2123 1460 2126
rect 1482 2123 1508 2126
rect 1530 2123 1548 2126
rect 1660 2123 1677 2126
rect 1700 2123 1717 2126
rect 1748 2123 1765 2126
rect 1892 2123 1917 2126
rect 1970 2125 1973 2133
rect 1978 2123 2004 2126
rect 2018 2123 2060 2126
rect 2066 2123 2092 2126
rect 2130 2123 2156 2126
rect 2162 2123 2180 2126
rect 2226 2123 2236 2126
rect 2300 2123 2309 2126
rect 2404 2123 2437 2126
rect 2450 2123 2460 2126
rect 2492 2123 2501 2126
rect 2514 2123 2556 2126
rect 2580 2123 2597 2126
rect 2642 2123 2676 2126
rect 236 2113 269 2116
rect 564 2113 597 2116
rect 602 2106 605 2115
rect 570 2103 605 2106
rect 650 2103 653 2123
rect 852 2113 869 2116
rect 884 2113 893 2116
rect 980 2113 1021 2116
rect 1468 2113 1477 2116
rect 1516 2113 1533 2116
rect 2020 2113 2045 2116
rect 2196 2113 2221 2116
rect 2252 2113 2277 2116
rect 2692 2113 2701 2116
rect 14 2067 2818 2073
rect 1170 2033 1220 2036
rect 1970 2033 1989 2036
rect 2018 2033 2052 2036
rect 1970 2026 1973 2033
rect 116 2013 141 2016
rect 268 2013 301 2016
rect 418 2013 428 2016
rect 434 2013 460 2016
rect 466 2006 469 2025
rect 620 2023 653 2026
rect 1178 2023 1204 2026
rect 1228 2023 1237 2026
rect 1828 2023 1853 2026
rect 1956 2023 1973 2026
rect 2010 2023 2036 2026
rect 2172 2023 2213 2026
rect 2260 2023 2269 2026
rect 1178 2016 1181 2023
rect 492 2013 501 2016
rect 506 2013 532 2016
rect 556 2013 581 2016
rect 594 2013 604 2016
rect 618 2013 669 2016
rect 740 2013 749 2016
rect 802 2013 812 2016
rect 866 2013 876 2016
rect 962 2013 988 2016
rect 1010 2013 1052 2016
rect 1164 2013 1181 2016
rect 1234 2013 1260 2016
rect 498 2006 501 2013
rect 250 2003 260 2006
rect 324 2003 333 2006
rect 338 2003 372 2006
rect 434 2003 452 2006
rect 466 2003 484 2006
rect 498 2003 540 2006
rect 554 2003 596 2006
rect 618 2005 621 2013
rect 1338 2006 1341 2014
rect 1434 2013 1444 2016
rect 1500 2013 1509 2016
rect 1524 2013 1557 2016
rect 1642 2013 1668 2016
rect 1674 2013 1692 2016
rect 1714 2013 1765 2016
rect 1772 2013 1789 2016
rect 1802 2013 1812 2016
rect 1922 2013 1940 2016
rect 2066 2013 2092 2016
rect 2116 2013 2125 2016
rect 2130 2013 2156 2016
rect 2170 2013 2221 2016
rect 2228 2013 2237 2016
rect 2242 2013 2252 2016
rect 2316 2013 2357 2016
rect 2396 2013 2421 2016
rect 2628 2013 2660 2016
rect 2666 2013 2676 2016
rect 658 2003 668 2006
rect 706 2003 732 2006
rect 746 2003 772 2006
rect 842 2003 868 2006
rect 906 2003 948 2006
rect 1002 2003 1044 2006
rect 1076 2003 1149 2006
rect 1258 2003 1268 2006
rect 1338 2003 1356 2006
rect 1370 2003 1404 2006
rect 1538 2003 1564 2006
rect 1626 2003 1660 2006
rect 1674 2003 1684 2006
rect 1706 2003 1740 2006
rect 1762 2005 1765 2013
rect 556 1993 581 1996
rect 746 1993 749 2003
rect 1082 1993 1124 1996
rect 1306 1993 1324 1996
rect 1338 1993 1348 1996
rect 1498 1993 1508 1996
rect 1786 1993 1789 2013
rect 1884 2003 1901 2006
rect 1956 2003 1965 2006
rect 2138 2003 2148 2006
rect 2170 2005 2173 2013
rect 2234 2006 2237 2013
rect 2210 2003 2220 2006
rect 2234 2003 2244 2006
rect 2282 2003 2308 2006
rect 2708 2003 2733 2006
rect 2730 1996 2733 2003
rect 2682 1993 2700 1996
rect 2714 1995 2733 1996
rect 2714 1993 2732 1995
rect 38 1967 2794 1973
rect 242 1943 261 1946
rect 258 1936 261 1943
rect 1202 1943 1229 1946
rect 1450 1943 1460 1946
rect 1540 1943 1557 1946
rect 2082 1943 2100 1946
rect 2114 1943 2124 1946
rect 2178 1943 2196 1946
rect 236 1933 253 1936
rect 258 1933 276 1936
rect 306 1933 324 1936
rect 338 1933 348 1936
rect 402 1926 405 1934
rect 570 1933 580 1936
rect 626 1933 652 1936
rect 698 1933 708 1936
rect 826 1933 844 1936
rect 882 1933 924 1936
rect 1026 1933 1060 1936
rect 1202 1926 1205 1943
rect 1210 1933 1236 1936
rect 1266 1933 1332 1936
rect 1348 1933 1412 1936
rect 1436 1933 1445 1936
rect 1468 1933 1517 1936
rect 1602 1933 1612 1936
rect 1626 1934 1660 1936
rect 1626 1933 1661 1934
rect 1682 1933 1708 1936
rect 1730 1933 1748 1936
rect 1780 1933 1797 1936
rect 1810 1933 1836 1936
rect 1898 1933 1908 1936
rect 1970 1933 1980 1936
rect 2060 1933 2085 1936
rect 2114 1933 2132 1936
rect 2204 1933 2220 1936
rect 2244 1933 2269 1936
rect 2346 1933 2356 1936
rect 2666 1933 2700 1936
rect 2722 1933 2732 1936
rect 204 1923 213 1926
rect 258 1923 284 1926
rect 332 1923 341 1926
rect 356 1923 405 1926
rect 426 1923 444 1926
rect 546 1923 588 1926
rect 730 1923 757 1926
rect 868 1923 893 1926
rect 898 1923 932 1926
rect 1050 1923 1068 1926
rect 1106 1923 1132 1926
rect 1138 1923 1205 1926
rect 1226 1923 1244 1926
rect 1370 1923 1420 1926
rect 1514 1925 1517 1933
rect 1546 1923 1580 1926
rect 1620 1923 1653 1926
rect 754 1916 757 1923
rect 890 1916 893 1923
rect 236 1913 269 1916
rect 620 1913 629 1916
rect 732 1913 749 1916
rect 754 1913 764 1916
rect 890 1913 909 1916
rect 948 1913 989 1916
rect 994 1906 997 1915
rect 762 1903 780 1906
rect 954 1903 997 1906
rect 1050 1903 1053 1923
rect 1658 1916 1661 1933
rect 1668 1923 1709 1926
rect 1716 1923 1725 1926
rect 1746 1923 1756 1926
rect 1868 1923 1909 1926
rect 1916 1923 1925 1926
rect 1962 1923 1988 1926
rect 1994 1923 2028 1926
rect 2068 1923 2077 1926
rect 2114 1925 2117 1933
rect 2218 1923 2228 1926
rect 2250 1923 2292 1926
rect 2330 1923 2364 1926
rect 2476 1923 2501 1926
rect 2602 1923 2620 1926
rect 2666 1925 2669 1933
rect 2730 1923 2740 1926
rect 1260 1913 1317 1916
rect 1628 1913 1661 1916
rect 1724 1913 1733 1916
rect 2580 1913 2589 1916
rect 1730 1893 1733 1913
rect 2370 1903 2388 1906
rect 14 1867 2818 1873
rect 268 1823 285 1826
rect 356 1823 365 1826
rect 524 1823 541 1826
rect 618 1823 645 1826
rect 740 1823 749 1826
rect 282 1816 285 1823
rect 770 1816 773 1846
rect 1778 1833 1797 1836
rect 2282 1833 2300 1836
rect 2322 1833 2357 1836
rect 2570 1833 2588 1836
rect 2634 1833 2652 1836
rect 1778 1826 1781 1833
rect 796 1823 821 1826
rect 860 1823 869 1826
rect 1228 1823 1269 1826
rect 1596 1823 1605 1826
rect 1732 1823 1741 1826
rect 1772 1823 1781 1826
rect 2188 1823 2197 1826
rect 2322 1823 2325 1833
rect 2636 1823 2645 1826
rect 2722 1816 2725 1825
rect 218 1813 252 1816
rect 282 1813 293 1816
rect 204 1803 213 1806
rect 226 1803 244 1806
rect 274 1803 300 1806
rect 306 1796 309 1814
rect 314 1813 348 1816
rect 394 1813 404 1816
rect 428 1813 437 1816
rect 490 1813 516 1816
rect 522 1813 580 1816
rect 586 1813 629 1816
rect 722 1813 732 1816
rect 770 1813 788 1816
rect 852 1813 901 1816
rect 964 1813 1005 1816
rect 1026 1813 1060 1816
rect 1090 1813 1109 1816
rect 1122 1813 1140 1816
rect 1162 1813 1212 1816
rect 1250 1813 1276 1816
rect 1314 1813 1364 1816
rect 1412 1813 1429 1816
rect 1500 1813 1509 1816
rect 1530 1813 1548 1816
rect 1570 1813 1580 1816
rect 1666 1813 1692 1816
rect 1724 1813 1756 1816
rect 1818 1813 1828 1816
rect 1884 1813 1900 1816
rect 1924 1813 1957 1816
rect 1964 1813 1980 1816
rect 2034 1813 2052 1816
rect 2082 1813 2116 1816
rect 2138 1813 2172 1816
rect 2460 1813 2477 1816
rect 2618 1813 2628 1816
rect 2666 1813 2692 1816
rect 2706 1813 2716 1816
rect 2722 1813 2740 1816
rect 442 1803 460 1806
rect 618 1803 660 1806
rect 684 1803 693 1806
rect 762 1803 780 1806
rect 826 1803 844 1806
rect 890 1803 900 1806
rect 1012 1803 1021 1806
rect 1106 1803 1109 1813
rect 1114 1803 1132 1806
rect 1170 1803 1204 1806
rect 1228 1803 1269 1806
rect 1300 1803 1309 1806
rect 1380 1803 1404 1806
rect 1426 1803 1429 1813
rect 1442 1803 1452 1806
rect 1482 1803 1492 1806
rect 1626 1803 1636 1806
rect 1660 1803 1677 1806
rect 1730 1803 1748 1806
rect 1938 1803 1956 1806
rect 2010 1803 2044 1806
rect 2082 1803 2108 1806
rect 2132 1803 2141 1806
rect 2188 1803 2204 1806
rect 2228 1803 2237 1806
rect 2698 1803 2708 1806
rect 2722 1803 2732 1806
rect 306 1793 317 1796
rect 762 1793 765 1803
rect 978 1793 1004 1796
rect 38 1767 2794 1773
rect 412 1743 421 1746
rect 490 1733 516 1736
rect 570 1733 612 1736
rect 658 1733 676 1736
rect 810 1733 828 1736
rect 866 1726 869 1734
rect 914 1726 917 1734
rect 970 1733 980 1736
rect 1050 1733 1092 1736
rect 1186 1733 1212 1736
rect 1268 1733 1301 1736
rect 1346 1733 1372 1736
rect 1298 1727 1301 1733
rect 132 1723 149 1726
rect 188 1723 197 1726
rect 260 1723 293 1726
rect 330 1723 340 1726
rect 354 1723 388 1726
rect 524 1723 541 1726
rect 546 1723 556 1726
rect 628 1723 637 1726
rect 698 1723 749 1726
rect 772 1723 797 1726
rect 836 1723 869 1726
rect 876 1723 917 1726
rect 954 1723 981 1726
rect 1044 1723 1093 1726
rect 1170 1723 1180 1726
rect 1298 1724 1316 1727
rect 1418 1726 1421 1734
rect 1396 1723 1421 1726
rect 1442 1726 1445 1734
rect 1450 1733 1476 1736
rect 1580 1733 1589 1736
rect 1594 1733 1620 1736
rect 1634 1733 1643 1736
rect 1666 1733 1676 1736
rect 1738 1733 1764 1736
rect 1786 1733 1804 1736
rect 1834 1726 1837 1734
rect 1922 1733 1956 1736
rect 2018 1726 2021 1734
rect 2042 1733 2068 1736
rect 2114 1733 2123 1736
rect 2162 1726 2165 1734
rect 2194 1726 2197 1736
rect 1442 1723 1453 1726
rect 1474 1723 1484 1726
rect 1500 1723 1556 1726
rect 1594 1723 1628 1726
rect 1653 1723 1661 1726
rect 1684 1723 1693 1726
rect 1698 1723 1716 1726
rect 1794 1723 1837 1726
rect 1938 1723 1964 1726
rect 1980 1723 2021 1726
rect 2058 1723 2076 1726
rect 2132 1723 2165 1726
rect 2172 1723 2197 1726
rect 2226 1725 2229 1736
rect 2354 1733 2380 1736
rect 2676 1733 2685 1736
rect 1698 1716 1701 1723
rect 476 1713 485 1716
rect 564 1713 597 1716
rect 780 1713 789 1716
rect 940 1713 965 1716
rect 1116 1713 1165 1716
rect 1308 1713 1317 1716
rect 1332 1713 1373 1716
rect 1690 1713 1701 1716
rect 1852 1713 1877 1716
rect 2180 1713 2205 1716
rect 2250 1713 2268 1716
rect 2274 1706 2277 1725
rect 2362 1723 2388 1726
rect 2562 1723 2588 1726
rect 2628 1723 2669 1726
rect 2684 1723 2716 1726
rect 2324 1713 2333 1716
rect 1282 1703 1324 1706
rect 2266 1703 2277 1706
rect 2306 1703 2340 1706
rect 14 1667 2818 1673
rect 660 1623 669 1626
rect 788 1623 821 1626
rect 844 1623 853 1626
rect 1076 1623 1117 1626
rect 1244 1623 1261 1626
rect 1580 1623 1597 1626
rect 1978 1623 1997 1626
rect 2028 1623 2045 1626
rect 2188 1623 2197 1626
rect 1978 1616 1981 1623
rect 234 1613 244 1616
rect 308 1613 317 1616
rect 396 1613 452 1616
rect 498 1613 516 1616
rect 522 1613 532 1616
rect 730 1613 748 1616
rect 762 1613 780 1616
rect 818 1613 836 1616
rect 890 1613 916 1616
rect 978 1613 988 1616
rect 1002 1613 1044 1616
rect 1050 1613 1060 1616
rect 1074 1613 1101 1616
rect 1132 1613 1165 1616
rect 1197 1613 1205 1616
rect 1332 1613 1373 1616
rect 1394 1613 1420 1616
rect 1426 1613 1469 1616
rect 1490 1613 1509 1616
rect 1516 1613 1533 1616
rect 1538 1613 1564 1616
rect 1714 1613 1748 1616
rect 1754 1613 1764 1616
rect 1778 1613 1820 1616
rect 1850 1613 1884 1616
rect 1898 1613 1916 1616
rect 1972 1613 1981 1616
rect 1986 1613 2012 1616
rect 2034 1613 2052 1616
rect 2074 1613 2100 1616
rect 2140 1613 2149 1616
rect 2330 1613 2356 1616
rect 2554 1613 2564 1616
rect 2618 1613 2629 1616
rect 2636 1613 2645 1616
rect 498 1606 501 1613
rect 1170 1606 1173 1613
rect 476 1603 501 1606
rect 554 1603 580 1606
rect 618 1603 636 1606
rect 730 1603 740 1606
rect 810 1603 828 1606
rect 842 1603 876 1606
rect 898 1603 908 1606
rect 1026 1603 1036 1606
rect 1082 1603 1124 1606
rect 1138 1603 1173 1606
rect 1218 1603 1228 1606
rect 1314 1603 1324 1606
rect 1380 1603 1405 1606
rect 1490 1605 1493 1613
rect 1586 1603 1612 1606
rect 1626 1603 1668 1606
rect 1794 1603 1812 1606
rect 1844 1603 1869 1606
rect 1922 1603 1964 1606
rect 1970 1603 2004 1606
rect 2034 1603 2037 1613
rect 2132 1603 2164 1606
rect 2188 1603 2205 1606
rect 2330 1603 2348 1606
rect 2372 1603 2405 1606
rect 2548 1603 2556 1606
rect 2618 1605 2621 1613
rect 2668 1603 2685 1606
rect 2722 1603 2732 1606
rect 268 1593 277 1596
rect 850 1593 868 1596
rect 994 1593 1013 1596
rect 1197 1593 1221 1596
rect 1354 1593 1372 1596
rect 1586 1593 1604 1596
rect 2106 1593 2123 1596
rect 922 1583 941 1586
rect 1586 1583 1589 1593
rect 38 1567 2794 1573
rect 298 1543 324 1546
rect 354 1543 364 1546
rect 450 1536 453 1546
rect 492 1543 509 1546
rect 610 1543 620 1546
rect 738 1543 748 1546
rect 738 1536 741 1543
rect 1410 1536 1413 1546
rect 1490 1543 1509 1546
rect 332 1533 349 1536
rect 354 1533 372 1536
rect 450 1533 469 1536
rect 354 1526 357 1533
rect 156 1523 181 1526
rect 276 1523 285 1526
rect 340 1523 357 1526
rect 380 1523 389 1526
rect 466 1525 469 1533
rect 490 1533 516 1536
rect 530 1533 564 1536
rect 628 1533 653 1536
rect 716 1533 741 1536
rect 756 1533 765 1536
rect 874 1533 900 1536
rect 932 1533 964 1536
rect 1028 1533 1061 1536
rect 1162 1533 1180 1536
rect 1204 1533 1237 1536
rect 1274 1533 1324 1536
rect 1410 1533 1428 1536
rect 1434 1533 1453 1536
rect 1476 1533 1501 1536
rect 490 1525 493 1533
rect 1058 1526 1061 1533
rect 524 1523 549 1526
rect 588 1523 597 1526
rect 668 1523 700 1526
rect 764 1523 773 1526
rect 818 1523 836 1526
rect 860 1523 869 1526
rect 874 1523 908 1526
rect 954 1523 972 1526
rect 978 1523 1004 1526
rect 1058 1523 1076 1526
rect 1092 1523 1125 1526
rect 1170 1523 1188 1526
rect 1210 1523 1244 1526
rect 1292 1523 1301 1526
rect 1346 1523 1372 1526
rect 1434 1525 1437 1533
rect 1506 1526 1509 1543
rect 1802 1543 1836 1546
rect 2570 1543 2612 1546
rect 1802 1536 1805 1543
rect 1580 1533 1589 1536
rect 1594 1533 1612 1536
rect 1644 1533 1669 1536
rect 1730 1533 1756 1536
rect 1794 1533 1805 1536
rect 1844 1533 1853 1536
rect 1858 1533 1868 1536
rect 1882 1533 1908 1536
rect 1484 1523 1493 1526
rect 1506 1523 1524 1526
rect 1602 1523 1620 1526
rect 1698 1523 1724 1526
rect 1794 1525 1797 1533
rect 1930 1526 1933 1534
rect 2034 1533 2052 1536
rect 2106 1533 2132 1536
rect 2234 1533 2244 1536
rect 2258 1533 2268 1536
rect 2290 1533 2324 1536
rect 2594 1533 2637 1536
rect 2674 1533 2716 1536
rect 1930 1523 1965 1526
rect 1978 1523 1996 1526
rect 2026 1523 2060 1526
rect 2074 1523 2092 1526
rect 2106 1523 2140 1526
rect 2154 1523 2188 1526
rect 2210 1523 2252 1526
rect 2266 1523 2276 1526
rect 2290 1523 2332 1526
rect 2508 1523 2533 1526
rect 2698 1523 2724 1526
rect 676 1513 685 1516
rect 716 1513 733 1516
rect 770 1513 788 1516
rect 1100 1513 1109 1516
rect 1122 1513 1132 1516
rect 1156 1513 1173 1516
rect 786 1503 804 1506
rect 1298 1503 1301 1523
rect 1388 1513 1405 1516
rect 1580 1513 1597 1516
rect 1700 1513 1709 1516
rect 1932 1513 1941 1516
rect 2100 1513 2117 1516
rect 2290 1513 2293 1523
rect 1402 1503 1405 1513
rect 14 1467 2818 1473
rect 452 1423 485 1426
rect 564 1423 573 1426
rect 932 1423 949 1426
rect 1172 1423 1197 1426
rect 1194 1416 1197 1423
rect 244 1413 269 1416
rect 346 1413 372 1416
rect 314 1403 332 1406
rect 370 1403 380 1406
rect 394 1403 397 1414
rect 508 1413 533 1416
rect 692 1413 701 1416
rect 812 1413 829 1416
rect 418 1403 428 1406
rect 458 1403 484 1406
rect 570 1403 596 1406
rect 660 1403 669 1406
rect 706 1403 740 1406
rect 786 1403 804 1406
rect 844 1403 853 1406
rect 914 1405 917 1416
rect 924 1413 933 1416
rect 962 1413 980 1416
rect 1085 1413 1109 1416
rect 1130 1413 1140 1416
rect 1164 1413 1173 1416
rect 1194 1413 1212 1416
rect 1226 1413 1260 1416
rect 1298 1413 1324 1416
rect 1356 1413 1381 1416
rect 1420 1413 1453 1416
rect 1514 1413 1525 1416
rect 1746 1413 1797 1416
rect 1812 1413 1837 1416
rect 1900 1413 1909 1416
rect 1916 1413 1965 1416
rect 1522 1406 1525 1413
rect 954 1403 972 1406
rect 1010 1403 1044 1406
rect 1146 1403 1156 1406
rect 1242 1403 1252 1406
rect 1298 1403 1332 1406
rect 1348 1403 1389 1406
rect 1434 1403 1460 1406
rect 1492 1403 1517 1406
rect 1522 1403 1532 1406
rect 1666 1403 1708 1406
rect 1714 1403 1732 1406
rect 1754 1403 1772 1406
rect 1804 1403 1821 1406
rect 1892 1403 1901 1406
rect 1514 1396 1517 1403
rect 578 1393 588 1396
rect 642 1393 652 1396
rect 1514 1393 1524 1396
rect 1674 1393 1700 1396
rect 1786 1393 1796 1396
rect 1874 1393 1884 1396
rect 1962 1395 1965 1413
rect 1972 1403 1981 1406
rect 1986 1405 1989 1416
rect 2132 1413 2141 1416
rect 2188 1413 2197 1416
rect 2212 1413 2221 1416
rect 2276 1413 2293 1416
rect 2564 1413 2589 1416
rect 2620 1413 2629 1416
rect 2684 1413 2709 1416
rect 2740 1413 2749 1416
rect 2012 1403 2021 1406
rect 2060 1403 2068 1406
rect 2228 1403 2237 1406
rect 2626 1403 2636 1406
rect 2746 1405 2749 1413
rect 38 1367 2794 1373
rect 498 1343 508 1346
rect 1210 1343 1220 1346
rect 1234 1343 1244 1346
rect 1858 1343 1876 1346
rect 156 1333 189 1336
rect 450 1333 460 1336
rect 474 1333 516 1336
rect 164 1323 173 1326
rect 186 1323 212 1326
rect 244 1323 277 1326
rect 332 1323 357 1326
rect 476 1323 485 1326
rect 524 1323 533 1326
rect 634 1325 637 1336
rect 690 1325 693 1336
rect 730 1326 733 1334
rect 770 1333 796 1336
rect 826 1333 860 1336
rect 890 1333 908 1336
rect 938 1333 972 1336
rect 1026 1333 1052 1336
rect 1084 1333 1125 1336
rect 716 1323 733 1326
rect 740 1323 797 1326
rect 868 1323 909 1326
rect 938 1316 941 1333
rect 1210 1326 1213 1343
rect 1234 1336 1237 1343
rect 2090 1336 2093 1346
rect 1228 1333 1237 1336
rect 1242 1333 1252 1336
rect 1258 1333 1277 1336
rect 1370 1333 1404 1336
rect 1466 1333 1484 1336
rect 1508 1333 1532 1336
rect 1562 1333 1588 1336
rect 1612 1333 1636 1336
rect 1658 1333 1676 1336
rect 1804 1333 1821 1336
rect 1828 1333 1853 1336
rect 1866 1333 1884 1336
rect 1890 1333 1924 1336
rect 1002 1323 1020 1326
rect 1026 1323 1060 1326
rect 1180 1323 1213 1326
rect 1242 1323 1245 1333
rect 1258 1325 1261 1333
rect 1274 1323 1308 1326
rect 1370 1323 1396 1326
rect 1434 1323 1460 1326
rect 1514 1323 1524 1326
rect 1570 1323 1596 1326
rect 1652 1323 1661 1326
rect 1700 1323 1709 1326
rect 1730 1323 1772 1326
rect 1940 1323 1965 1326
rect 1970 1325 1973 1336
rect 2018 1333 2028 1336
rect 2090 1333 2108 1336
rect 2362 1333 2396 1336
rect 2418 1333 2429 1336
rect 2490 1333 2524 1336
rect 1996 1323 2005 1326
rect 2026 1323 2036 1326
rect 2106 1323 2116 1326
rect 2276 1323 2333 1326
rect 2418 1325 2421 1333
rect 2442 1323 2484 1326
rect 2636 1323 2645 1326
rect 820 1313 829 1316
rect 932 1313 941 1316
rect 14 1267 2818 1273
rect 170 1213 212 1216
rect 258 1213 292 1216
rect 324 1213 333 1216
rect 508 1213 517 1216
rect 564 1213 573 1216
rect 620 1213 629 1216
rect 242 1203 300 1206
rect 700 1203 709 1206
rect 754 1203 757 1214
rect 780 1213 789 1216
rect 844 1213 853 1216
rect 866 1206 869 1214
rect 1044 1213 1053 1216
rect 1106 1206 1109 1214
rect 1228 1213 1261 1216
rect 1274 1206 1277 1214
rect 772 1203 789 1206
rect 810 1203 828 1206
rect 842 1203 853 1206
rect 866 1203 908 1206
rect 980 1203 997 1206
rect 1002 1203 1028 1206
rect 1106 1203 1124 1206
rect 1130 1203 1172 1206
rect 1194 1203 1212 1206
rect 1226 1203 1268 1206
rect 1274 1203 1292 1206
rect 1298 1203 1301 1214
rect 1354 1206 1357 1214
rect 1386 1213 1420 1216
rect 1434 1213 1460 1216
rect 1556 1213 1565 1216
rect 1644 1213 1661 1216
rect 1740 1213 1749 1216
rect 1844 1213 1869 1216
rect 1964 1213 1973 1216
rect 2012 1213 2029 1216
rect 2220 1213 2229 1216
rect 2242 1213 2284 1216
rect 2290 1213 2300 1216
rect 2484 1213 2501 1216
rect 2580 1213 2589 1216
rect 2700 1213 2717 1216
rect 1354 1203 1372 1206
rect 1394 1203 1412 1206
rect 1436 1203 1453 1206
rect 1516 1203 1548 1206
rect 1562 1203 1572 1206
rect 2266 1203 2276 1206
rect 2306 1203 2324 1206
rect 2346 1203 2396 1206
rect 682 1193 692 1196
rect 730 1193 740 1196
rect 850 1195 853 1203
rect 890 1193 900 1196
rect 1194 1193 1197 1203
rect 1234 1193 1260 1196
rect 1274 1193 1284 1196
rect 1306 1193 1340 1196
rect 38 1167 2794 1173
rect 418 1136 421 1146
rect 1106 1143 1148 1146
rect 1314 1143 1340 1146
rect 1354 1143 1364 1146
rect 1954 1136 1957 1156
rect 2466 1143 2492 1146
rect 2506 1143 2580 1146
rect 2594 1143 2636 1146
rect 2650 1143 2660 1146
rect 418 1133 468 1136
rect 1156 1133 1205 1136
rect 1338 1133 1348 1136
rect 1372 1133 1389 1136
rect 1604 1133 1637 1136
rect 1788 1133 1813 1136
rect 1948 1133 1957 1136
rect 2042 1133 2092 1136
rect 2114 1133 2156 1136
rect 2668 1133 2717 1136
rect 338 1126 356 1127
rect 164 1123 189 1126
rect 300 1124 356 1126
rect 300 1123 341 1124
rect 492 1123 533 1126
rect 538 1123 556 1126
rect 620 1123 645 1126
rect 700 1123 709 1126
rect 932 1123 949 1126
rect 1100 1123 1125 1126
rect 1202 1123 1205 1133
rect 1252 1123 1261 1126
rect 1522 1123 1556 1126
rect 1634 1123 1637 1133
rect 1754 1123 1764 1126
rect 1874 1123 1908 1126
rect 1954 1123 1996 1126
rect 2116 1123 2149 1126
rect 2228 1123 2253 1126
rect 2508 1123 2541 1126
rect 2596 1123 2605 1126
rect 2676 1123 2709 1126
rect 348 1113 357 1116
rect 1698 1113 1749 1116
rect 306 1103 364 1106
rect 14 1067 2818 1073
rect 186 1006 189 1026
rect 292 1023 341 1026
rect 380 1023 437 1026
rect 220 1013 237 1016
rect 290 1013 364 1016
rect 434 1013 444 1016
rect 476 1013 485 1016
rect 490 1013 532 1016
rect 570 1013 628 1016
rect 692 1013 741 1016
rect 788 1013 797 1016
rect 964 1013 973 1016
rect 1180 1013 1205 1016
rect 1236 1013 1277 1016
rect 1380 1013 1389 1016
rect 1532 1013 1541 1016
rect 1588 1013 1597 1016
rect 1732 1013 1741 1016
rect 1884 1013 1901 1016
rect 1914 1013 1948 1016
rect 2004 1013 2021 1016
rect 2026 1013 2036 1016
rect 2084 1013 2109 1016
rect 2324 1013 2333 1016
rect 2364 1013 2381 1016
rect 2386 1006 2389 1016
rect 2484 1013 2517 1016
rect 2530 1013 2572 1016
rect 2602 1013 2612 1016
rect 106 1003 116 1006
rect 186 1003 212 1006
rect 306 1003 356 1006
rect 380 1003 413 1006
rect 556 1003 581 1006
rect 634 1003 668 1006
rect 1476 1003 1485 1006
rect 1802 1003 1860 1006
rect 1882 1003 1940 1006
rect 1970 1003 1996 1006
rect 2052 1003 2069 1006
rect 2210 1003 2276 1006
rect 2290 1003 2316 1006
rect 2386 1003 2476 1006
rect 2594 1003 2604 1006
rect 130 993 204 996
rect 2250 993 2268 996
rect 2290 993 2308 996
rect 2370 993 2468 996
rect 38 967 2794 973
rect 242 936 245 956
rect 586 943 596 946
rect 610 943 620 946
rect 2058 943 2068 946
rect 220 933 229 936
rect 242 933 252 936
rect 266 933 292 936
rect 316 933 333 936
rect 570 933 604 936
rect 634 933 684 936
rect 706 933 716 936
rect 730 933 772 936
rect 858 933 868 936
rect 116 923 125 926
rect 172 923 189 926
rect 194 923 204 926
rect 242 923 260 926
rect 314 923 364 926
rect 370 923 380 926
rect 474 923 482 926
rect 490 923 532 926
rect 890 925 893 936
rect 914 933 924 936
rect 938 933 980 936
rect 1010 933 1052 936
rect 908 923 925 926
rect 932 923 965 926
rect 1004 923 1021 926
rect 1034 923 1044 926
rect 1076 923 1125 926
rect 1162 925 1165 936
rect 1170 933 1180 936
rect 1202 933 1244 936
rect 1178 923 1188 926
rect 1274 923 1277 934
rect 1570 933 1596 936
rect 1612 933 1629 936
rect 1986 933 2012 936
rect 2042 933 2076 936
rect 2170 933 2196 936
rect 2442 933 2460 936
rect 2618 933 2628 936
rect 2652 933 2661 936
rect 1396 923 1405 926
rect 1530 923 1548 926
rect 1740 923 1749 926
rect 1924 923 1949 926
rect 2020 923 2036 926
rect 2106 923 2124 926
rect 2298 923 2309 926
rect 2380 923 2389 926
rect 2620 923 2629 926
rect 242 916 245 923
rect 220 913 245 916
rect 268 913 285 916
rect 316 913 341 916
rect 396 913 429 916
rect 2236 913 2269 916
rect 2298 915 2301 923
rect 2652 913 2661 916
rect 802 903 820 906
rect 14 867 2818 873
rect 530 833 564 836
rect 260 823 293 826
rect 290 816 293 823
rect 116 813 133 816
rect 172 813 197 816
rect 204 813 244 816
rect 290 813 308 816
rect 412 813 421 816
rect 468 813 485 816
rect 194 805 197 813
rect 530 806 533 833
rect 1122 826 1125 856
rect 1138 833 1157 836
rect 1914 833 1932 836
rect 538 823 548 826
rect 572 823 605 826
rect 602 816 605 823
rect 626 823 637 826
rect 692 823 749 826
rect 626 816 629 823
rect 762 816 765 825
rect 794 823 813 826
rect 892 823 901 826
rect 932 823 941 826
rect 970 823 1005 826
rect 1122 823 1148 826
rect 602 813 613 816
rect 620 813 629 816
rect 634 813 652 816
rect 658 813 676 816
rect 690 813 749 816
rect 762 813 780 816
rect 210 803 236 806
rect 282 803 300 806
rect 338 803 388 806
rect 500 803 533 806
rect 610 805 613 813
rect 746 806 749 813
rect 794 806 797 823
rect 844 813 869 816
rect 890 813 924 816
rect 938 813 1004 816
rect 1100 813 1109 816
rect 1116 813 1141 816
rect 1154 815 1157 833
rect 1916 823 1925 826
rect 2116 823 2133 826
rect 2204 823 2229 826
rect 2244 823 2269 826
rect 1218 813 1244 816
rect 1276 813 1293 816
rect 1332 813 1341 816
rect 1362 813 1372 816
rect 1460 813 1469 816
rect 1636 813 1645 816
rect 1748 813 1765 816
rect 1804 813 1829 816
rect 2060 813 2077 816
rect 2084 813 2100 816
rect 2114 813 2172 816
rect 2202 813 2236 816
rect 2306 813 2349 816
rect 2356 813 2389 816
rect 2418 813 2445 816
rect 2492 813 2524 816
rect 2556 813 2565 816
rect 738 805 749 806
rect 738 803 748 805
rect 786 803 797 806
rect 866 805 869 813
rect 1074 803 1092 806
rect 1178 803 1196 806
rect 1210 803 1252 806
rect 1418 803 1436 806
rect 1538 803 1548 806
rect 1578 803 1612 806
rect 1634 803 1644 806
rect 1666 803 1700 806
rect 2074 805 2077 813
rect 2210 803 2228 806
rect 2258 803 2268 806
rect 2346 805 2349 813
rect 2396 803 2437 806
rect 2442 805 2445 813
rect 2498 803 2532 806
rect 2554 803 2596 806
rect 2626 805 2629 816
rect 2636 813 2645 816
rect 794 796 797 803
rect 482 793 492 796
rect 794 793 820 796
rect 1178 793 1188 796
rect 2370 793 2388 796
rect 38 767 2794 773
rect 1338 736 1341 746
rect 1578 743 1588 746
rect 1650 743 1660 746
rect 2266 743 2284 746
rect 2362 743 2372 746
rect 212 733 293 736
rect 298 733 316 736
rect 426 733 460 736
rect 570 733 580 736
rect 602 733 637 736
rect 668 733 685 736
rect 762 733 788 736
rect 818 733 852 736
rect 874 733 924 736
rect 948 733 957 736
rect 962 733 980 736
rect 1018 733 1052 736
rect 1076 733 1085 736
rect 1202 733 1228 736
rect 1274 733 1300 736
rect 1338 733 1372 736
rect 1386 733 1396 736
rect 340 723 349 726
rect 354 723 404 726
rect 484 723 501 726
rect 506 723 532 726
rect 562 723 572 726
rect 602 725 605 733
rect 610 723 644 726
rect 690 723 708 726
rect 762 725 765 733
rect 826 723 844 726
rect 922 723 932 726
rect 988 723 997 726
rect 1074 723 1100 726
rect 1114 723 1164 726
rect 1226 723 1253 726
rect 1260 723 1285 726
rect 1324 723 1349 726
rect 420 713 453 716
rect 812 713 837 716
rect 1386 715 1389 733
rect 1434 726 1437 734
rect 1450 733 1469 736
rect 1450 726 1453 733
rect 1404 723 1437 726
rect 1444 723 1453 726
rect 1458 723 1492 726
rect 1506 723 1556 726
rect 1570 723 1573 734
rect 1578 733 1596 736
rect 1602 733 1661 736
rect 1668 733 1701 736
rect 1754 733 1788 736
rect 1882 733 1900 736
rect 1954 733 1964 736
rect 2138 733 2148 736
rect 2178 733 2212 736
rect 2250 733 2292 736
rect 2306 733 2340 736
rect 2380 733 2429 736
rect 2450 733 2460 736
rect 2498 733 2524 736
rect 2554 733 2572 736
rect 2594 733 2604 736
rect 1602 725 1605 733
rect 1508 713 1541 716
rect 1572 713 1581 716
rect 1698 706 1701 733
rect 1738 723 1748 726
rect 1802 723 1812 726
rect 1914 723 1948 726
rect 1972 723 1981 726
rect 1986 723 2004 726
rect 2018 723 2044 726
rect 2082 723 2116 726
rect 2130 723 2156 726
rect 2178 723 2220 726
rect 2226 723 2244 726
rect 2300 723 2309 726
rect 2348 723 2373 726
rect 2434 723 2444 726
rect 2450 723 2453 733
rect 2634 726 2637 734
rect 2484 723 2516 726
rect 2548 723 2565 726
rect 2626 723 2637 726
rect 1986 716 1989 723
rect 1826 713 1852 716
rect 1876 713 1885 716
rect 1980 713 1989 716
rect 2452 713 2461 716
rect 1698 703 1724 706
rect 14 667 2818 673
rect 452 623 469 626
rect 500 623 533 626
rect 564 623 581 626
rect 794 616 797 636
rect 1698 633 1724 636
rect 2170 633 2212 636
rect 108 613 133 616
rect 164 613 173 616
rect 260 613 285 616
rect 330 613 356 616
rect 380 613 429 616
rect 514 613 548 616
rect 562 613 604 616
rect 642 613 692 616
rect 788 613 797 616
rect 802 613 828 616
rect 860 613 877 616
rect 932 613 941 616
rect 948 613 989 616
rect 1052 613 1084 616
rect 1140 613 1149 616
rect 1188 613 1213 616
rect 1362 613 1380 616
rect 1452 613 1476 616
rect 1564 613 1581 616
rect 1604 613 1613 616
rect 986 606 989 613
rect 1698 606 1701 633
rect 1810 616 1813 625
rect 1890 616 1893 625
rect 2186 623 2196 626
rect 2220 623 2253 626
rect 2466 616 2469 625
rect 1738 613 1748 616
rect 1810 613 1828 616
rect 1834 613 1876 616
rect 1890 613 1908 616
rect 2004 613 2036 616
rect 2068 613 2125 616
rect 2260 613 2285 616
rect 178 603 196 606
rect 394 603 428 606
rect 452 603 461 606
rect 466 603 476 606
rect 506 603 540 606
rect 794 603 836 606
rect 890 603 908 606
rect 978 605 989 606
rect 978 603 988 605
rect 1026 603 1036 606
rect 1100 603 1132 606
rect 1186 603 1228 606
rect 1250 603 1284 606
rect 1314 603 1324 606
rect 1362 603 1372 606
rect 1412 603 1421 606
rect 1426 603 1444 606
rect 1498 603 1524 606
rect 1610 603 1620 606
rect 1668 603 1701 606
rect 1754 603 1788 606
rect 1834 603 1868 606
rect 1914 603 1956 606
rect 1970 603 1980 606
rect 2018 603 2044 606
rect 2074 603 2092 606
rect 2242 603 2252 606
rect 2314 605 2317 616
rect 2380 613 2389 616
rect 2442 606 2445 616
rect 2450 613 2460 616
rect 2466 613 2484 616
rect 2548 613 2556 616
rect 2628 613 2637 616
rect 2716 613 2725 616
rect 2442 603 2452 606
rect 2500 603 2524 606
rect 2554 603 2564 606
rect 2690 603 2708 606
rect 170 593 188 596
rect 1018 593 1028 596
rect 1626 593 1660 596
rect 38 567 2794 573
rect 306 543 316 546
rect 194 526 197 535
rect 282 533 324 536
rect 410 533 420 536
rect 788 533 797 536
rect 802 533 828 536
rect 874 533 884 536
rect 908 533 917 536
rect 1146 533 1172 536
rect 1196 533 1205 536
rect 1210 533 1220 536
rect 1244 533 1261 536
rect 1322 533 1388 536
rect 1412 533 1429 536
rect 1434 533 1476 536
rect 1500 533 1509 536
rect 1514 533 1540 536
rect 1564 533 1573 536
rect 1578 533 1596 536
rect 1620 533 1629 536
rect 1642 533 1660 536
rect 1706 533 1764 536
rect 1786 533 1828 536
rect 1858 533 1900 536
rect 1930 533 1980 536
rect 2002 533 2036 536
rect 1434 526 1437 533
rect 2274 526 2277 545
rect 2284 533 2317 536
rect 2418 533 2484 536
rect 2554 526 2557 535
rect 2580 533 2637 536
rect 2748 533 2757 536
rect 108 523 133 526
rect 164 523 197 526
rect 204 523 220 526
rect 332 523 428 526
rect 660 523 685 526
rect 716 523 733 526
rect 738 523 772 526
rect 826 523 836 526
rect 882 523 892 526
rect 1084 523 1093 526
rect 1218 523 1228 526
rect 1250 523 1300 526
rect 1378 523 1396 526
rect 1410 523 1437 526
rect 1788 523 1805 526
rect 1852 523 1885 526
rect 1924 523 1972 526
rect 2004 523 2029 526
rect 2044 523 2061 526
rect 2066 523 2092 526
rect 2130 523 2164 526
rect 2202 523 2236 526
rect 2260 523 2277 526
rect 2492 523 2557 526
rect 2692 523 2701 526
rect 236 513 309 516
rect 444 513 453 516
rect 852 513 869 516
rect 1250 503 1253 523
rect 1308 513 1325 516
rect 1412 513 1469 516
rect 1500 513 1533 516
rect 1620 513 1653 516
rect 2052 513 2085 516
rect 14 467 2818 473
rect 890 426 893 436
rect 2178 426 2181 436
rect 884 423 893 426
rect 908 423 925 426
rect 988 423 1013 426
rect 2164 423 2181 426
rect 1010 416 1013 423
rect 164 413 181 416
rect 324 413 333 416
rect 372 413 397 416
rect 708 413 733 416
rect 796 413 868 416
rect 882 413 893 416
rect 1010 413 1028 416
rect 1148 413 1157 416
rect 1178 413 1236 416
rect 1372 413 1381 416
rect 1420 413 1445 416
rect 1490 413 1516 416
rect 1580 413 1613 416
rect 1636 413 1725 416
rect 1788 413 1845 416
rect 1860 413 1876 416
rect 1882 413 1924 416
rect 2052 413 2061 416
rect 2108 413 2125 416
rect 2162 413 2196 416
rect 2420 413 2429 416
rect 2484 413 2493 416
rect 2546 413 2556 416
rect 770 403 788 406
rect 834 403 860 406
rect 882 405 885 413
rect 954 403 964 406
rect 1010 403 1020 406
rect 1042 403 1060 406
rect 1090 403 1140 406
rect 1252 403 1277 406
rect 1490 403 1493 413
rect 1714 403 1724 406
rect 1748 403 1757 406
rect 1852 403 1861 406
rect 1906 403 1932 406
rect 2114 403 2148 406
rect 2292 403 2301 406
rect 2412 403 2437 406
rect 770 393 780 396
rect 1066 393 1132 396
rect 2298 393 2301 403
rect 2362 393 2404 396
rect 38 367 2794 373
rect 186 343 244 346
rect 386 343 420 346
rect 498 343 532 346
rect 586 336 589 346
rect 602 343 628 346
rect 690 343 732 346
rect 252 333 269 336
rect 428 333 461 336
rect 546 333 556 336
rect 586 333 636 336
rect 754 333 764 336
rect 1018 327 1021 335
rect 1450 333 1476 336
rect 1732 333 1741 336
rect 1930 333 1972 336
rect 2026 333 2060 336
rect 2202 333 2220 336
rect 260 323 269 326
rect 282 323 308 326
rect 372 323 389 326
rect 476 323 493 326
rect 564 323 597 326
rect 676 323 693 326
rect 836 323 853 326
rect 892 323 901 326
rect 956 323 981 326
rect 1012 324 1021 327
rect 2418 326 2421 335
rect 2538 333 2548 336
rect 2572 333 2589 336
rect 2620 333 2636 336
rect 1084 323 1101 326
rect 1220 323 1229 326
rect 1340 323 1365 326
rect 1420 323 1437 326
rect 1452 323 1484 326
rect 1660 323 1685 326
rect 1716 323 1725 326
rect 1740 323 1756 326
rect 1874 323 1900 326
rect 1938 323 1964 326
rect 2002 323 2020 326
rect 2140 323 2157 326
rect 2210 323 2228 326
rect 2250 323 2260 326
rect 2404 323 2421 326
rect 316 313 365 316
rect 2028 313 2053 316
rect 2076 313 2101 316
rect 2442 306 2445 325
rect 2474 313 2484 316
rect 2490 306 2493 325
rect 2514 323 2524 326
rect 2530 323 2556 326
rect 2578 323 2604 326
rect 2652 323 2661 326
rect 2700 323 2725 326
rect 2434 303 2445 306
rect 2466 303 2493 306
rect 14 267 2818 273
rect 244 223 285 226
rect 364 223 389 226
rect 484 223 493 226
rect 546 216 549 226
rect 1020 223 1037 226
rect 2548 223 2565 226
rect 180 213 228 216
rect 266 213 348 216
rect 428 213 468 216
rect 540 213 588 216
rect 636 213 676 216
rect 746 213 756 216
rect 884 213 909 216
rect 940 213 997 216
rect 1108 213 1148 216
rect 1236 213 1308 216
rect 1388 213 1460 216
rect 1844 213 1869 216
rect 1956 213 1972 216
rect 2052 213 2069 216
rect 2114 213 2148 216
rect 210 203 220 206
rect 306 203 340 206
rect 442 203 460 206
rect 642 203 668 206
rect 706 203 748 206
rect 772 203 813 206
rect 946 203 996 206
rect 1026 203 1052 206
rect 1114 203 1140 206
rect 1164 203 1181 206
rect 1274 203 1300 206
rect 1362 203 1380 206
rect 1434 203 1452 206
rect 1906 203 1948 206
rect 2282 203 2324 206
rect 2450 205 2453 216
rect 2460 213 2469 216
rect 2476 213 2532 216
rect 2506 203 2524 206
rect 2548 203 2557 206
rect 2562 205 2565 223
rect 2572 213 2605 216
rect 2644 213 2661 216
rect 2700 213 2709 216
rect 2602 203 2605 213
rect 1058 193 1092 196
rect 1170 193 1220 196
rect 1330 193 1372 196
rect 2282 193 2316 196
rect 38 167 2794 173
rect 1562 143 1580 146
rect 1850 143 1876 146
rect 2050 143 2108 146
rect 2354 143 2372 146
rect 1050 126 1053 135
rect 1588 133 1597 136
rect 1834 133 1884 136
rect 2116 133 2141 136
rect 2380 133 2397 136
rect 2420 133 2477 136
rect 2538 133 2580 136
rect 2612 133 2661 136
rect 172 123 197 126
rect 292 123 317 126
rect 412 123 437 126
rect 540 123 565 126
rect 660 123 685 126
rect 804 123 813 126
rect 956 123 981 126
rect 1012 123 1053 126
rect 1060 123 1069 126
rect 1292 123 1317 126
rect 1396 123 1413 126
rect 1500 123 1525 126
rect 1556 123 1581 126
rect 1596 123 1612 126
rect 1772 123 1797 126
rect 1828 123 1845 126
rect 1892 123 1908 126
rect 1980 123 2005 126
rect 2124 123 2141 126
rect 2236 123 2253 126
rect 2394 125 2397 133
rect 2428 123 2485 126
rect 2522 123 2532 126
rect 2588 123 2605 126
rect 14 67 2818 73
rect 38 37 2794 57
rect 14 13 2818 33
<< metal2 >>
rect 14 13 34 2627
rect 38 37 58 2603
rect 1178 2566 1181 2586
rect 322 2543 349 2546
rect 394 2543 397 2566
rect 402 2543 405 2556
rect 450 2543 461 2546
rect 186 2416 189 2426
rect 130 2393 133 2406
rect 90 1946 93 2336
rect 138 2323 141 2416
rect 162 2383 165 2406
rect 170 2403 173 2416
rect 178 2413 189 2416
rect 178 2346 181 2413
rect 186 2393 189 2406
rect 162 2343 181 2346
rect 162 2246 165 2343
rect 194 2336 197 2436
rect 250 2423 285 2426
rect 298 2423 301 2536
rect 322 2533 325 2543
rect 306 2523 325 2526
rect 330 2523 333 2536
rect 346 2533 349 2543
rect 386 2533 397 2536
rect 386 2526 389 2533
rect 450 2526 453 2543
rect 474 2533 477 2546
rect 482 2533 485 2556
rect 370 2523 389 2526
rect 322 2436 325 2516
rect 306 2433 325 2436
rect 266 2413 277 2416
rect 282 2413 285 2423
rect 210 2386 213 2406
rect 226 2403 237 2406
rect 210 2383 221 2386
rect 242 2383 245 2406
rect 258 2383 261 2396
rect 162 2243 173 2246
rect 146 2213 149 2226
rect 170 2216 173 2243
rect 178 2223 181 2336
rect 190 2333 197 2336
rect 190 2236 193 2333
rect 190 2233 197 2236
rect 154 2213 165 2216
rect 170 2213 181 2216
rect 122 2133 125 2146
rect 170 2143 173 2206
rect 178 2136 181 2213
rect 186 2143 189 2206
rect 162 2133 181 2136
rect 138 2013 141 2126
rect 162 2026 165 2133
rect 194 2116 197 2233
rect 202 2186 205 2326
rect 218 2256 221 2383
rect 242 2336 245 2346
rect 242 2333 261 2336
rect 274 2323 277 2413
rect 306 2406 309 2433
rect 210 2253 221 2256
rect 210 2226 213 2253
rect 234 2233 277 2236
rect 210 2223 221 2226
rect 234 2223 237 2233
rect 210 2203 213 2216
rect 202 2183 209 2186
rect 158 2023 165 2026
rect 186 2113 197 2116
rect 158 1966 161 2023
rect 146 1963 161 1966
rect 90 1943 109 1946
rect 106 1686 109 1943
rect 146 1836 149 1963
rect 146 1833 165 1836
rect 138 1773 141 1806
rect 146 1723 149 1816
rect 162 1813 165 1833
rect 170 1766 173 2016
rect 186 1966 189 2113
rect 206 2106 209 2183
rect 218 2156 221 2223
rect 266 2216 269 2226
rect 226 2183 229 2216
rect 258 2213 269 2216
rect 274 2213 277 2233
rect 218 2153 229 2156
rect 218 2133 221 2146
rect 202 2103 209 2106
rect 186 1963 197 1966
rect 178 1933 181 1946
rect 186 1893 189 1946
rect 194 1833 197 1963
rect 202 1836 205 2103
rect 218 1993 221 2006
rect 226 2003 229 2153
rect 242 2016 245 2206
rect 258 2123 261 2213
rect 274 2193 277 2206
rect 282 2146 285 2406
rect 298 2403 309 2406
rect 314 2383 317 2406
rect 290 2326 293 2346
rect 290 2323 297 2326
rect 294 2266 297 2323
rect 306 2276 309 2356
rect 306 2273 313 2276
rect 294 2263 301 2266
rect 298 2206 301 2263
rect 310 2226 313 2273
rect 290 2203 301 2206
rect 306 2223 313 2226
rect 290 2193 293 2203
rect 306 2196 309 2223
rect 298 2193 309 2196
rect 282 2143 293 2146
rect 266 2096 269 2116
rect 258 2093 269 2096
rect 258 2026 261 2093
rect 258 2023 269 2026
rect 238 2013 245 2016
rect 238 1966 241 2013
rect 238 1963 245 1966
rect 210 1933 213 1946
rect 242 1943 245 1963
rect 250 1933 253 2006
rect 210 1903 213 1926
rect 218 1923 245 1926
rect 202 1833 213 1836
rect 186 1813 189 1826
rect 194 1823 205 1826
rect 178 1793 181 1806
rect 194 1796 197 1823
rect 210 1816 213 1833
rect 190 1793 197 1796
rect 202 1813 213 1816
rect 170 1763 177 1766
rect 174 1686 177 1763
rect 190 1736 193 1793
rect 202 1746 205 1813
rect 210 1773 213 1806
rect 202 1743 209 1746
rect 106 1683 133 1686
rect 130 1443 133 1683
rect 170 1683 177 1686
rect 186 1733 193 1736
rect 170 1446 173 1683
rect 186 1673 189 1733
rect 194 1656 197 1726
rect 190 1653 197 1656
rect 178 1523 181 1586
rect 190 1576 193 1653
rect 206 1646 209 1743
rect 202 1643 209 1646
rect 190 1573 197 1576
rect 162 1443 173 1446
rect 138 1333 141 1366
rect 162 1346 165 1443
rect 186 1373 189 1436
rect 162 1343 173 1346
rect 130 1256 133 1326
rect 146 1273 149 1326
rect 170 1323 173 1343
rect 186 1333 189 1346
rect 194 1333 197 1573
rect 130 1253 165 1256
rect 82 1143 85 1206
rect 106 1126 109 1216
rect 122 1156 125 1246
rect 162 1213 165 1253
rect 98 1123 109 1126
rect 118 1153 125 1156
rect 98 1036 101 1123
rect 118 1106 121 1153
rect 118 1103 125 1106
rect 98 1033 109 1036
rect 90 1003 93 1016
rect 98 986 101 1016
rect 106 1003 109 1033
rect 122 1026 125 1103
rect 138 1076 141 1146
rect 138 1073 149 1076
rect 114 1023 133 1026
rect 114 996 117 1023
rect 106 993 117 996
rect 122 986 125 1016
rect 130 993 133 1023
rect 146 1016 149 1073
rect 138 1013 149 1016
rect 98 983 125 986
rect 90 656 93 936
rect 114 913 117 983
rect 138 966 141 1013
rect 162 976 165 996
rect 134 963 141 966
rect 158 973 165 976
rect 122 923 125 946
rect 134 886 137 963
rect 158 886 161 973
rect 170 896 173 1216
rect 186 1133 189 1326
rect 202 1293 205 1643
rect 218 1536 221 1836
rect 226 1733 229 1916
rect 242 1906 245 1923
rect 238 1903 245 1906
rect 238 1836 241 1903
rect 238 1833 245 1836
rect 234 1613 237 1816
rect 242 1716 245 1833
rect 250 1786 253 1926
rect 258 1923 261 1966
rect 266 1956 269 2023
rect 274 2013 277 2126
rect 266 1953 277 1956
rect 266 1913 269 1946
rect 258 1806 261 1826
rect 274 1813 277 1953
rect 282 1936 285 2136
rect 290 2123 293 2143
rect 298 2036 301 2193
rect 306 2123 309 2186
rect 314 2123 317 2206
rect 322 2166 325 2426
rect 354 2366 357 2416
rect 338 2363 357 2366
rect 338 2333 341 2363
rect 338 2213 341 2316
rect 362 2236 365 2426
rect 386 2373 389 2406
rect 394 2336 397 2526
rect 442 2523 453 2526
rect 442 2456 445 2523
rect 442 2453 453 2456
rect 450 2436 453 2453
rect 402 2423 429 2426
rect 402 2403 405 2423
rect 410 2383 413 2416
rect 394 2333 405 2336
rect 394 2313 397 2326
rect 346 2233 365 2236
rect 346 2206 349 2233
rect 330 2173 333 2206
rect 338 2203 349 2206
rect 354 2203 357 2216
rect 322 2163 329 2166
rect 326 2046 329 2163
rect 338 2133 341 2203
rect 362 2196 365 2226
rect 370 2203 373 2216
rect 378 2213 381 2306
rect 354 2193 365 2196
rect 326 2043 333 2046
rect 290 2033 301 2036
rect 290 1976 293 2033
rect 298 2023 325 2026
rect 298 2013 301 2023
rect 298 1983 301 2006
rect 306 2003 309 2016
rect 290 1973 317 1976
rect 282 1933 293 1936
rect 298 1933 301 1956
rect 306 1933 309 1946
rect 290 1916 293 1933
rect 314 1923 317 1973
rect 286 1913 293 1916
rect 286 1846 289 1913
rect 298 1903 301 1916
rect 322 1906 325 2006
rect 330 2003 333 2043
rect 314 1903 325 1906
rect 330 1936 333 1996
rect 338 1973 341 2126
rect 346 2106 349 2136
rect 354 2123 357 2193
rect 362 2133 365 2146
rect 346 2103 353 2106
rect 350 1956 353 2103
rect 362 2013 365 2036
rect 370 1986 373 2166
rect 378 2033 381 2206
rect 386 2123 389 2226
rect 394 2213 397 2286
rect 402 2196 405 2333
rect 410 2283 413 2316
rect 418 2273 421 2406
rect 426 2403 429 2423
rect 442 2386 445 2436
rect 450 2433 457 2436
rect 466 2433 469 2526
rect 434 2383 445 2386
rect 434 2276 437 2383
rect 454 2376 457 2433
rect 490 2413 493 2526
rect 498 2523 501 2536
rect 514 2433 517 2526
rect 530 2523 533 2536
rect 546 2533 549 2556
rect 562 2543 589 2546
rect 562 2533 565 2543
rect 498 2396 501 2426
rect 450 2373 457 2376
rect 482 2393 501 2396
rect 450 2306 453 2373
rect 458 2333 461 2346
rect 466 2323 469 2336
rect 450 2303 469 2306
rect 434 2273 445 2276
rect 442 2256 445 2273
rect 442 2253 453 2256
rect 410 2213 413 2236
rect 398 2193 405 2196
rect 410 2193 413 2206
rect 378 2003 381 2016
rect 386 2003 389 2106
rect 398 2046 401 2193
rect 418 2186 421 2246
rect 410 2183 421 2186
rect 398 2043 405 2046
rect 394 2013 397 2026
rect 370 1983 381 1986
rect 338 1946 341 1956
rect 350 1953 373 1956
rect 338 1943 365 1946
rect 330 1933 341 1936
rect 282 1843 289 1846
rect 314 1846 317 1903
rect 314 1843 325 1846
rect 258 1803 269 1806
rect 274 1793 277 1806
rect 250 1783 277 1786
rect 250 1733 269 1736
rect 266 1716 269 1733
rect 242 1713 253 1716
rect 250 1626 253 1713
rect 262 1713 269 1716
rect 262 1636 265 1713
rect 262 1633 269 1636
rect 242 1623 253 1626
rect 242 1596 245 1623
rect 266 1613 269 1633
rect 238 1593 245 1596
rect 218 1533 229 1536
rect 210 1433 213 1526
rect 226 1476 229 1533
rect 218 1473 229 1476
rect 218 1453 221 1473
rect 238 1456 241 1593
rect 250 1586 253 1606
rect 250 1583 261 1586
rect 238 1453 245 1456
rect 218 1403 221 1446
rect 186 1023 189 1126
rect 186 923 189 1016
rect 194 933 205 936
rect 194 913 197 926
rect 170 893 181 896
rect 134 883 141 886
rect 158 883 165 886
rect 130 803 133 816
rect 138 666 141 883
rect 162 756 165 883
rect 178 766 181 893
rect 202 876 205 933
rect 210 926 213 1376
rect 218 1333 221 1366
rect 226 1313 229 1326
rect 226 1213 229 1306
rect 218 1196 221 1206
rect 234 1203 237 1346
rect 242 1303 245 1453
rect 250 1313 253 1536
rect 258 1523 261 1583
rect 266 1426 269 1536
rect 274 1513 277 1783
rect 282 1523 285 1843
rect 290 1823 317 1826
rect 290 1813 293 1823
rect 314 1813 317 1823
rect 322 1806 325 1843
rect 290 1793 293 1806
rect 298 1803 325 1806
rect 330 1803 333 1933
rect 338 1923 357 1926
rect 338 1886 341 1906
rect 338 1883 349 1886
rect 346 1826 349 1883
rect 338 1823 349 1826
rect 362 1823 365 1943
rect 290 1723 293 1746
rect 298 1733 301 1803
rect 290 1696 293 1716
rect 306 1703 309 1726
rect 290 1693 297 1696
rect 294 1626 297 1693
rect 290 1623 297 1626
rect 290 1593 293 1623
rect 298 1543 301 1606
rect 258 1423 269 1426
rect 242 1213 245 1296
rect 258 1273 261 1423
rect 266 1393 269 1416
rect 298 1366 301 1416
rect 274 1363 301 1366
rect 274 1323 277 1363
rect 266 1226 269 1316
rect 290 1286 293 1306
rect 290 1283 297 1286
rect 266 1223 273 1226
rect 242 1196 245 1206
rect 258 1196 261 1216
rect 218 1193 245 1196
rect 242 1153 245 1193
rect 254 1193 261 1196
rect 254 1136 257 1193
rect 270 1166 273 1223
rect 218 1123 221 1136
rect 250 1133 257 1136
rect 266 1163 273 1166
rect 266 1133 269 1163
rect 250 1086 253 1133
rect 274 1093 277 1136
rect 250 1083 261 1086
rect 258 1016 261 1083
rect 282 1026 285 1276
rect 294 1156 297 1283
rect 306 1263 309 1446
rect 314 1423 317 1796
rect 338 1766 341 1823
rect 338 1763 365 1766
rect 330 1733 333 1746
rect 322 1686 325 1726
rect 330 1703 333 1726
rect 346 1713 349 1756
rect 322 1683 333 1686
rect 330 1436 333 1683
rect 354 1626 357 1726
rect 362 1696 365 1763
rect 370 1743 373 1953
rect 378 1703 381 1983
rect 386 1966 389 1986
rect 386 1963 393 1966
rect 390 1846 393 1963
rect 386 1843 393 1846
rect 386 1793 389 1843
rect 394 1813 397 1826
rect 394 1716 397 1736
rect 390 1713 397 1716
rect 362 1693 381 1696
rect 346 1623 357 1626
rect 346 1593 349 1623
rect 354 1603 357 1616
rect 362 1613 365 1636
rect 378 1623 381 1693
rect 390 1646 393 1713
rect 390 1643 397 1646
rect 370 1603 381 1606
rect 386 1603 389 1626
rect 354 1543 357 1556
rect 322 1433 333 1436
rect 314 1393 317 1406
rect 322 1393 325 1433
rect 338 1373 341 1416
rect 346 1413 349 1536
rect 226 933 229 946
rect 210 923 221 926
rect 218 906 221 923
rect 218 903 225 906
rect 202 873 213 876
rect 210 803 213 873
rect 222 826 225 903
rect 218 823 225 826
rect 154 753 165 756
rect 170 763 181 766
rect 154 686 157 753
rect 154 683 161 686
rect 138 663 149 666
rect 90 653 117 656
rect 82 593 85 606
rect 114 576 117 653
rect 130 613 133 626
rect 82 573 117 576
rect 146 576 149 663
rect 158 626 161 683
rect 158 623 165 626
rect 162 606 165 623
rect 170 613 173 763
rect 194 733 197 746
rect 162 603 173 606
rect 178 603 181 626
rect 146 573 157 576
rect 82 463 85 573
rect 130 523 133 546
rect 154 486 157 573
rect 138 483 157 486
rect 138 403 141 483
rect 170 426 173 603
rect 186 433 189 726
rect 202 723 213 726
rect 218 723 221 823
rect 234 813 237 1016
rect 254 1013 261 1016
rect 274 1023 285 1026
rect 290 1153 297 1156
rect 274 1013 277 1023
rect 290 1013 293 1153
rect 306 1143 309 1216
rect 314 1183 317 1216
rect 330 1213 333 1336
rect 354 1323 357 1406
rect 370 1403 373 1603
rect 386 1453 389 1526
rect 394 1426 397 1643
rect 378 1423 397 1426
rect 378 1336 381 1423
rect 386 1403 397 1406
rect 374 1333 381 1336
rect 346 1313 357 1316
rect 346 1166 349 1313
rect 374 1286 377 1333
rect 386 1313 389 1326
rect 362 1283 377 1286
rect 362 1236 365 1283
rect 394 1243 397 1396
rect 358 1233 365 1236
rect 358 1176 361 1233
rect 402 1213 405 2043
rect 410 1993 413 2183
rect 426 2056 429 2226
rect 434 2163 437 2206
rect 442 2143 445 2216
rect 458 2186 461 2296
rect 466 2213 469 2303
rect 474 2223 477 2336
rect 482 2323 485 2393
rect 506 2356 509 2416
rect 514 2393 517 2416
rect 522 2403 525 2446
rect 530 2403 533 2416
rect 498 2353 509 2356
rect 490 2306 493 2336
rect 486 2303 493 2306
rect 486 2236 489 2303
rect 486 2233 493 2236
rect 466 2193 469 2206
rect 458 2183 469 2186
rect 434 2133 453 2136
rect 426 2053 437 2056
rect 418 2013 421 2036
rect 434 2013 437 2053
rect 418 2003 437 2006
rect 418 1933 429 1936
rect 434 1933 437 1986
rect 410 1923 429 1926
rect 442 1916 445 2126
rect 450 2123 453 2133
rect 450 2103 453 2116
rect 418 1806 421 1916
rect 426 1903 429 1916
rect 438 1913 445 1916
rect 438 1836 441 1913
rect 438 1833 445 1836
rect 410 1803 421 1806
rect 410 1723 413 1736
rect 378 1193 381 1206
rect 358 1173 365 1176
rect 242 953 245 966
rect 254 926 257 1013
rect 266 933 269 1006
rect 290 963 293 1006
rect 254 923 261 926
rect 298 923 301 1136
rect 306 1093 309 1106
rect 306 936 309 1006
rect 306 933 317 936
rect 314 923 317 933
rect 258 816 261 923
rect 282 913 317 916
rect 314 896 317 913
rect 306 893 317 896
rect 306 846 309 893
rect 306 843 317 846
rect 258 813 269 816
rect 226 786 229 806
rect 250 803 261 806
rect 226 783 237 786
rect 210 693 213 723
rect 234 686 237 783
rect 210 683 237 686
rect 210 626 213 683
rect 210 623 217 626
rect 266 623 269 813
rect 282 803 285 836
rect 290 733 293 756
rect 298 733 301 746
rect 306 713 309 726
rect 314 636 317 843
rect 322 826 325 1166
rect 338 1163 349 1166
rect 338 1106 341 1163
rect 362 1156 365 1173
rect 354 1153 389 1156
rect 354 1113 357 1153
rect 338 1103 349 1106
rect 338 1013 341 1026
rect 330 833 333 936
rect 338 913 341 926
rect 346 836 349 1103
rect 370 1096 373 1116
rect 362 1093 373 1096
rect 362 1046 365 1093
rect 378 1056 381 1146
rect 386 1123 389 1153
rect 378 1053 389 1056
rect 362 1043 373 1046
rect 370 956 373 1043
rect 354 953 373 956
rect 354 933 357 953
rect 362 933 373 936
rect 346 833 353 836
rect 322 823 341 826
rect 322 723 325 746
rect 330 733 333 756
rect 338 733 341 823
rect 350 746 353 833
rect 362 803 365 933
rect 370 916 373 926
rect 386 916 389 1053
rect 402 1016 405 1186
rect 410 1143 413 1706
rect 418 1613 421 1776
rect 426 1563 429 1796
rect 434 1583 437 1816
rect 442 1803 445 1833
rect 442 1603 445 1796
rect 450 1746 453 2006
rect 458 1983 461 2136
rect 466 2096 469 2183
rect 474 2113 477 2206
rect 482 2203 485 2216
rect 490 2156 493 2233
rect 482 2153 493 2156
rect 482 2123 485 2153
rect 498 2146 501 2353
rect 506 2296 509 2316
rect 506 2293 513 2296
rect 510 2196 513 2293
rect 522 2203 525 2366
rect 538 2243 541 2526
rect 570 2523 573 2536
rect 578 2493 581 2536
rect 586 2533 589 2543
rect 602 2533 605 2546
rect 626 2543 653 2546
rect 546 2413 549 2426
rect 546 2303 549 2326
rect 530 2213 533 2236
rect 538 2223 549 2226
rect 506 2193 513 2196
rect 538 2193 541 2216
rect 554 2206 557 2436
rect 602 2423 605 2526
rect 626 2523 629 2543
rect 562 2313 565 2326
rect 570 2293 573 2406
rect 586 2403 589 2416
rect 610 2393 613 2406
rect 570 2213 573 2236
rect 546 2203 557 2206
rect 506 2173 509 2193
rect 490 2143 501 2146
rect 466 2093 473 2096
rect 470 1996 473 2093
rect 482 2003 485 2026
rect 466 1993 473 1996
rect 466 1976 469 1993
rect 462 1973 469 1976
rect 462 1856 465 1973
rect 474 1903 477 1976
rect 482 1923 485 1936
rect 490 1903 493 2143
rect 506 2116 509 2146
rect 502 2113 509 2116
rect 502 2036 505 2113
rect 514 2093 517 2136
rect 530 2113 533 2146
rect 538 2083 541 2156
rect 546 2126 549 2203
rect 578 2196 581 2346
rect 586 2323 605 2326
rect 618 2323 621 2336
rect 586 2306 589 2323
rect 586 2303 597 2306
rect 594 2226 597 2303
rect 554 2193 581 2196
rect 586 2223 597 2226
rect 554 2136 557 2193
rect 554 2133 565 2136
rect 546 2123 565 2126
rect 498 2033 505 2036
rect 498 1883 501 2033
rect 506 1953 509 2016
rect 458 1853 465 1856
rect 458 1806 461 1853
rect 466 1833 493 1836
rect 466 1813 469 1833
rect 482 1813 485 1826
rect 490 1813 493 1833
rect 506 1826 509 1926
rect 514 1896 517 2006
rect 522 1913 525 1936
rect 530 1923 533 1946
rect 546 1923 549 2016
rect 554 1963 557 2006
rect 562 1956 565 2123
rect 570 2093 573 2106
rect 578 2013 581 2126
rect 578 1963 581 1996
rect 586 1956 589 2223
rect 602 2193 605 2206
rect 610 2183 613 2196
rect 594 2143 605 2146
rect 594 2113 597 2143
rect 602 2123 613 2126
rect 594 2013 597 2026
rect 554 1953 565 1956
rect 582 1953 589 1956
rect 538 1903 541 1916
rect 514 1893 525 1896
rect 498 1823 509 1826
rect 522 1826 525 1893
rect 522 1823 533 1826
rect 458 1803 493 1806
rect 450 1743 477 1746
rect 450 1543 453 1736
rect 474 1733 477 1743
rect 458 1723 469 1726
rect 466 1616 469 1723
rect 482 1713 485 1746
rect 490 1713 493 1803
rect 498 1773 501 1823
rect 506 1813 525 1816
rect 506 1803 509 1813
rect 530 1796 533 1823
rect 526 1793 533 1796
rect 498 1666 501 1766
rect 506 1726 509 1746
rect 506 1723 517 1726
rect 494 1663 501 1666
rect 466 1613 477 1616
rect 458 1536 461 1606
rect 474 1573 477 1613
rect 418 1533 461 1536
rect 418 1403 421 1516
rect 426 1493 429 1526
rect 442 1446 445 1526
rect 434 1443 445 1446
rect 434 1413 437 1443
rect 418 1346 421 1366
rect 418 1343 429 1346
rect 426 1266 429 1343
rect 450 1333 453 1406
rect 458 1393 461 1496
rect 466 1356 469 1566
rect 474 1363 477 1536
rect 466 1353 477 1356
rect 466 1343 469 1353
rect 474 1343 477 1353
rect 474 1326 477 1336
rect 482 1333 485 1646
rect 494 1616 497 1663
rect 514 1656 517 1723
rect 526 1716 529 1793
rect 538 1763 541 1826
rect 554 1756 557 1953
rect 570 1863 573 1936
rect 582 1856 585 1953
rect 602 1946 605 2123
rect 618 2116 621 2206
rect 626 2123 629 2326
rect 634 2316 637 2536
rect 650 2526 653 2543
rect 690 2533 693 2546
rect 714 2533 725 2536
rect 642 2503 645 2526
rect 650 2523 661 2526
rect 658 2513 661 2523
rect 674 2513 677 2526
rect 698 2523 717 2526
rect 658 2423 669 2426
rect 658 2363 661 2423
rect 666 2353 669 2396
rect 642 2343 669 2346
rect 642 2333 645 2343
rect 634 2313 661 2316
rect 658 2266 661 2313
rect 666 2293 669 2343
rect 674 2266 677 2486
rect 682 2313 685 2416
rect 658 2263 665 2266
rect 674 2263 685 2266
rect 650 2213 653 2256
rect 634 2193 645 2196
rect 650 2193 653 2206
rect 642 2136 645 2193
rect 662 2166 665 2263
rect 658 2163 665 2166
rect 634 2133 645 2136
rect 650 2116 653 2146
rect 594 1943 605 1946
rect 610 2113 621 2116
rect 626 2113 653 2116
rect 610 1946 613 2113
rect 618 2066 621 2106
rect 650 2093 653 2106
rect 658 2086 661 2163
rect 634 2083 661 2086
rect 618 2063 625 2066
rect 622 1996 625 2063
rect 618 1993 625 1996
rect 618 1973 621 1993
rect 610 1943 621 1946
rect 594 1926 597 1943
rect 602 1933 613 1936
rect 594 1923 605 1926
rect 578 1853 585 1856
rect 570 1773 573 1806
rect 554 1753 561 1756
rect 538 1723 541 1736
rect 546 1733 549 1746
rect 526 1713 533 1716
rect 506 1653 517 1656
rect 506 1633 509 1653
rect 490 1613 497 1616
rect 522 1613 525 1636
rect 490 1516 493 1613
rect 498 1603 509 1606
rect 498 1533 501 1556
rect 506 1543 509 1566
rect 522 1553 525 1606
rect 530 1563 533 1713
rect 546 1623 549 1726
rect 558 1646 561 1753
rect 554 1643 561 1646
rect 554 1616 557 1643
rect 570 1626 573 1736
rect 578 1726 581 1853
rect 594 1826 597 1916
rect 586 1823 597 1826
rect 602 1823 605 1923
rect 610 1883 613 1926
rect 618 1823 621 1943
rect 626 1923 629 1956
rect 586 1743 589 1823
rect 626 1813 629 1916
rect 602 1803 621 1806
rect 634 1803 637 2083
rect 650 1946 653 2026
rect 658 2003 661 2016
rect 666 2013 669 2146
rect 674 2013 677 2216
rect 682 2076 685 2263
rect 690 2083 693 2406
rect 698 2403 701 2523
rect 714 2503 717 2516
rect 730 2403 733 2546
rect 746 2516 749 2536
rect 742 2513 749 2516
rect 742 2446 745 2513
rect 738 2443 745 2446
rect 738 2396 741 2443
rect 698 2393 741 2396
rect 698 2123 701 2393
rect 706 2283 709 2326
rect 714 2323 717 2376
rect 722 2333 725 2386
rect 746 2353 749 2436
rect 706 2183 709 2206
rect 706 2133 709 2166
rect 714 2143 717 2216
rect 722 2203 725 2296
rect 730 2273 733 2326
rect 738 2316 741 2336
rect 746 2333 749 2346
rect 738 2313 745 2316
rect 742 2266 745 2313
rect 738 2263 745 2266
rect 730 2203 733 2216
rect 714 2116 717 2136
rect 706 2113 717 2116
rect 682 2073 693 2076
rect 690 2013 693 2073
rect 706 2036 709 2113
rect 698 2033 709 2036
rect 642 1926 645 1946
rect 650 1943 669 1946
rect 642 1923 661 1926
rect 666 1893 669 1943
rect 674 1866 677 1926
rect 650 1863 677 1866
rect 618 1756 621 1803
rect 614 1753 621 1756
rect 578 1723 585 1726
rect 582 1646 585 1723
rect 594 1713 597 1726
rect 602 1713 605 1726
rect 614 1706 617 1753
rect 626 1733 629 1746
rect 634 1723 637 1776
rect 642 1716 645 1826
rect 634 1713 645 1716
rect 614 1703 621 1706
rect 542 1613 557 1616
rect 562 1623 573 1626
rect 578 1643 585 1646
rect 542 1556 545 1613
rect 538 1553 545 1556
rect 490 1513 501 1516
rect 498 1436 501 1513
rect 530 1496 533 1536
rect 538 1503 541 1553
rect 546 1523 549 1536
rect 522 1493 533 1496
rect 490 1433 501 1436
rect 450 1323 477 1326
rect 418 1263 429 1266
rect 418 1143 421 1263
rect 482 1223 485 1326
rect 490 1313 493 1433
rect 498 1343 501 1356
rect 458 1136 461 1216
rect 514 1213 517 1226
rect 482 1193 485 1206
rect 522 1186 525 1366
rect 530 1323 533 1416
rect 538 1403 541 1496
rect 554 1463 557 1606
rect 562 1436 565 1623
rect 570 1546 573 1616
rect 578 1603 581 1643
rect 586 1613 589 1626
rect 570 1543 589 1546
rect 570 1533 581 1536
rect 586 1526 589 1543
rect 570 1513 573 1526
rect 582 1523 589 1526
rect 554 1433 565 1436
rect 546 1386 549 1416
rect 542 1383 549 1386
rect 542 1306 545 1383
rect 554 1316 557 1433
rect 570 1413 573 1506
rect 582 1466 585 1523
rect 594 1516 597 1646
rect 602 1613 605 1636
rect 618 1603 621 1703
rect 634 1636 637 1713
rect 650 1643 653 1863
rect 666 1813 669 1846
rect 682 1836 685 2006
rect 698 2003 701 2033
rect 706 2003 709 2016
rect 674 1833 685 1836
rect 658 1733 661 1806
rect 666 1643 669 1746
rect 626 1633 637 1636
rect 626 1586 629 1633
rect 642 1613 661 1616
rect 622 1583 629 1586
rect 610 1533 613 1546
rect 622 1526 625 1583
rect 618 1523 625 1526
rect 634 1523 637 1566
rect 594 1513 605 1516
rect 578 1463 585 1466
rect 562 1393 565 1406
rect 570 1343 573 1406
rect 578 1393 581 1463
rect 578 1333 581 1356
rect 586 1323 589 1426
rect 602 1353 605 1513
rect 618 1343 621 1523
rect 642 1393 645 1586
rect 658 1553 661 1606
rect 666 1543 669 1626
rect 650 1503 653 1536
rect 658 1483 661 1536
rect 666 1416 669 1456
rect 658 1413 669 1416
rect 626 1316 629 1336
rect 634 1333 637 1376
rect 554 1313 565 1316
rect 542 1303 549 1306
rect 426 1133 461 1136
rect 426 1046 429 1133
rect 458 1106 461 1126
rect 450 1103 461 1106
rect 450 1056 453 1103
rect 450 1053 461 1056
rect 398 1013 405 1016
rect 422 1043 429 1046
rect 398 956 401 1013
rect 398 953 405 956
rect 370 913 389 916
rect 370 886 373 906
rect 394 903 397 936
rect 370 883 381 886
rect 378 836 381 883
rect 370 833 381 836
rect 370 786 373 833
rect 346 743 353 746
rect 366 783 373 786
rect 346 723 349 743
rect 298 633 317 636
rect 202 523 205 616
rect 214 556 217 623
rect 210 553 217 556
rect 234 556 237 606
rect 234 553 245 556
rect 170 423 189 426
rect 170 343 173 423
rect 178 333 181 416
rect 186 343 189 423
rect 186 213 189 326
rect 170 176 173 206
rect 210 203 213 553
rect 234 533 237 546
rect 218 413 221 436
rect 242 403 245 553
rect 282 533 285 616
rect 298 496 301 633
rect 314 613 317 626
rect 330 596 333 616
rect 322 593 333 596
rect 306 543 309 576
rect 322 516 325 593
rect 338 516 341 716
rect 354 693 357 726
rect 366 676 369 783
rect 378 683 381 816
rect 394 813 397 826
rect 402 753 405 953
rect 410 736 413 1006
rect 422 936 425 1043
rect 458 1033 461 1053
rect 434 1023 445 1026
rect 418 933 425 936
rect 418 896 421 933
rect 434 923 437 1016
rect 450 1013 461 1016
rect 450 993 453 1006
rect 442 933 445 946
rect 442 923 453 926
rect 426 913 437 916
rect 418 893 429 896
rect 426 836 429 893
rect 458 886 461 936
rect 466 933 469 1146
rect 474 1106 477 1166
rect 482 1123 485 1186
rect 514 1183 525 1186
rect 474 1103 485 1106
rect 482 1036 485 1103
rect 514 1056 517 1183
rect 530 1123 533 1186
rect 546 1163 549 1303
rect 562 1236 565 1313
rect 618 1313 629 1316
rect 618 1266 621 1313
rect 618 1263 629 1266
rect 554 1233 565 1236
rect 554 1176 557 1233
rect 570 1183 573 1216
rect 626 1213 629 1263
rect 642 1256 645 1346
rect 638 1253 645 1256
rect 554 1173 573 1176
rect 546 1133 549 1146
rect 514 1053 525 1056
rect 474 1033 485 1036
rect 474 933 477 1033
rect 514 1016 517 1036
rect 482 933 485 1016
rect 466 893 469 926
rect 474 886 477 926
rect 458 883 477 886
rect 418 833 429 836
rect 418 813 421 833
rect 458 803 461 826
rect 366 673 373 676
rect 346 603 349 616
rect 362 596 365 626
rect 370 603 373 673
rect 386 596 389 636
rect 362 593 389 596
rect 394 593 397 736
rect 406 733 413 736
rect 406 636 409 733
rect 406 633 413 636
rect 410 613 413 633
rect 362 523 365 536
rect 306 513 325 516
rect 330 513 341 516
rect 298 493 317 496
rect 266 333 269 416
rect 298 333 301 346
rect 266 306 269 326
rect 258 303 269 306
rect 258 236 261 303
rect 258 233 269 236
rect 266 213 269 233
rect 282 223 285 326
rect 314 313 317 493
rect 330 413 333 513
rect 346 376 349 466
rect 370 396 373 566
rect 386 436 389 576
rect 410 516 413 536
rect 402 513 413 516
rect 402 466 405 513
rect 402 463 413 466
rect 338 373 349 376
rect 362 393 373 396
rect 382 433 389 436
rect 338 306 341 373
rect 362 333 365 393
rect 382 386 385 433
rect 394 413 397 426
rect 382 383 389 386
rect 386 343 389 383
rect 362 313 381 316
rect 338 303 349 306
rect 170 173 229 176
rect 146 133 149 146
rect 194 123 197 166
rect 226 123 229 173
rect 242 163 245 206
rect 290 196 293 206
rect 306 203 309 226
rect 346 206 349 303
rect 386 223 389 326
rect 410 223 413 463
rect 418 343 421 736
rect 426 726 429 746
rect 426 723 437 726
rect 466 723 469 816
rect 482 813 485 926
rect 490 923 493 1016
rect 510 1013 517 1016
rect 498 806 501 966
rect 510 936 513 1013
rect 510 933 517 936
rect 514 916 517 933
rect 522 926 525 1053
rect 538 1016 541 1126
rect 570 1046 573 1173
rect 594 1156 597 1206
rect 638 1196 641 1253
rect 638 1193 645 1196
rect 658 1193 661 1413
rect 666 1393 669 1406
rect 674 1393 677 1833
rect 682 1813 685 1826
rect 690 1803 693 1986
rect 698 1933 701 1976
rect 722 1936 725 2146
rect 738 2133 741 2263
rect 754 2216 757 2536
rect 762 2523 765 2556
rect 794 2543 821 2546
rect 922 2543 925 2566
rect 1170 2563 1181 2566
rect 954 2543 973 2546
rect 794 2533 797 2543
rect 770 2473 773 2516
rect 802 2463 805 2526
rect 810 2523 813 2536
rect 818 2533 821 2543
rect 762 2413 765 2426
rect 778 2423 781 2446
rect 834 2433 837 2536
rect 858 2446 861 2526
rect 866 2523 869 2536
rect 898 2533 925 2536
rect 970 2533 973 2543
rect 978 2536 981 2546
rect 986 2543 997 2546
rect 1050 2543 1069 2546
rect 978 2533 997 2536
rect 898 2523 901 2533
rect 858 2443 869 2446
rect 866 2423 869 2443
rect 762 2323 765 2406
rect 770 2403 781 2406
rect 778 2336 781 2356
rect 774 2333 781 2336
rect 746 2213 757 2216
rect 746 2196 749 2213
rect 762 2206 765 2236
rect 774 2226 777 2333
rect 834 2326 837 2346
rect 842 2343 845 2386
rect 786 2266 789 2326
rect 826 2323 837 2326
rect 786 2263 797 2266
rect 774 2223 781 2226
rect 754 2203 765 2206
rect 746 2193 757 2196
rect 770 2193 773 2206
rect 754 2136 757 2193
rect 778 2176 781 2223
rect 786 2203 789 2216
rect 794 2206 797 2263
rect 826 2246 829 2323
rect 842 2293 845 2326
rect 826 2243 837 2246
rect 802 2223 829 2226
rect 834 2223 837 2243
rect 802 2213 805 2223
rect 810 2206 813 2216
rect 826 2206 829 2223
rect 794 2203 821 2206
rect 826 2203 837 2206
rect 750 2133 757 2136
rect 770 2173 789 2176
rect 770 2133 773 2173
rect 786 2146 789 2173
rect 786 2143 797 2146
rect 750 2036 753 2133
rect 722 1933 733 1936
rect 714 1856 717 1926
rect 714 1853 725 1856
rect 722 1813 725 1853
rect 730 1806 733 1926
rect 722 1803 733 1806
rect 690 1696 693 1726
rect 698 1713 701 1726
rect 682 1693 693 1696
rect 682 1676 685 1693
rect 682 1673 689 1676
rect 686 1556 689 1673
rect 698 1603 701 1666
rect 706 1613 709 1746
rect 714 1703 717 1736
rect 722 1666 725 1803
rect 730 1713 733 1746
rect 738 1706 741 2036
rect 750 2033 757 2036
rect 746 2003 749 2016
rect 746 1943 749 1996
rect 746 1913 749 1926
rect 746 1723 749 1826
rect 738 1703 745 1706
rect 722 1663 733 1666
rect 682 1553 689 1556
rect 682 1513 685 1553
rect 706 1546 709 1606
rect 698 1543 709 1546
rect 690 1523 693 1536
rect 698 1506 701 1543
rect 706 1533 717 1536
rect 694 1503 701 1506
rect 694 1446 697 1503
rect 690 1443 697 1446
rect 682 1376 685 1406
rect 674 1373 685 1376
rect 674 1326 677 1373
rect 690 1333 693 1443
rect 698 1393 701 1416
rect 706 1403 709 1506
rect 722 1493 725 1616
rect 730 1613 733 1663
rect 730 1583 733 1606
rect 742 1536 745 1703
rect 754 1596 757 2033
rect 762 1996 765 2126
rect 778 2026 781 2136
rect 794 2123 797 2136
rect 802 2133 805 2166
rect 770 2023 781 2026
rect 770 2006 773 2023
rect 786 2016 789 2046
rect 778 2013 789 2016
rect 794 2006 797 2016
rect 802 2013 805 2026
rect 770 2003 781 2006
rect 786 2003 797 2006
rect 802 2003 813 2006
rect 762 1993 773 1996
rect 762 1853 765 1976
rect 770 1843 773 1993
rect 778 1826 781 2003
rect 786 1913 789 1926
rect 794 1826 797 2003
rect 774 1823 781 1826
rect 786 1823 797 1826
rect 762 1706 765 1796
rect 774 1726 777 1823
rect 786 1733 789 1823
rect 774 1723 781 1726
rect 762 1703 773 1706
rect 762 1603 765 1616
rect 770 1603 773 1703
rect 778 1696 781 1723
rect 786 1713 789 1726
rect 794 1713 797 1816
rect 802 1696 805 1856
rect 810 1796 813 1976
rect 818 1943 821 2203
rect 842 2183 845 2216
rect 850 2166 853 2416
rect 882 2346 885 2516
rect 922 2396 925 2526
rect 978 2523 989 2526
rect 994 2436 997 2526
rect 1042 2446 1045 2526
rect 1050 2523 1053 2536
rect 1066 2533 1069 2543
rect 1106 2543 1141 2546
rect 1018 2443 1045 2446
rect 994 2433 1005 2436
rect 914 2393 925 2396
rect 914 2346 917 2393
rect 882 2343 889 2346
rect 914 2343 925 2346
rect 930 2343 933 2376
rect 858 2283 861 2326
rect 842 2163 853 2166
rect 858 2163 861 2226
rect 842 2096 845 2163
rect 866 2133 869 2246
rect 874 2186 877 2336
rect 886 2256 889 2343
rect 882 2253 889 2256
rect 882 2233 885 2253
rect 898 2223 901 2316
rect 906 2293 909 2326
rect 882 2206 885 2216
rect 914 2213 917 2306
rect 922 2296 925 2343
rect 938 2313 941 2386
rect 954 2326 957 2406
rect 978 2353 981 2416
rect 970 2333 973 2346
rect 954 2323 989 2326
rect 994 2306 997 2426
rect 1002 2416 1005 2433
rect 1002 2413 1009 2416
rect 1006 2306 1009 2413
rect 978 2303 997 2306
rect 1002 2303 1009 2306
rect 922 2293 933 2296
rect 930 2216 933 2293
rect 922 2213 933 2216
rect 954 2223 973 2226
rect 882 2203 909 2206
rect 874 2183 881 2186
rect 842 2093 853 2096
rect 826 1876 829 1936
rect 834 1923 837 2056
rect 842 2003 845 2076
rect 850 1973 853 2093
rect 858 1946 861 2126
rect 866 2113 869 2126
rect 878 2106 881 2183
rect 890 2113 893 2186
rect 922 2166 925 2213
rect 954 2206 957 2223
rect 970 2213 973 2223
rect 978 2206 981 2303
rect 1002 2283 1005 2303
rect 1018 2266 1021 2443
rect 1026 2403 1029 2436
rect 1050 2406 1053 2456
rect 1034 2403 1053 2406
rect 1050 2393 1053 2403
rect 1066 2366 1069 2526
rect 1098 2516 1101 2536
rect 1106 2523 1109 2543
rect 1090 2513 1101 2516
rect 1090 2426 1093 2513
rect 1090 2423 1101 2426
rect 1034 2363 1069 2366
rect 1010 2263 1021 2266
rect 986 2213 989 2236
rect 1010 2206 1013 2263
rect 954 2203 965 2206
rect 970 2203 981 2206
rect 946 2183 949 2196
rect 914 2163 925 2166
rect 874 2103 881 2106
rect 866 2013 869 2026
rect 858 1943 869 1946
rect 842 1923 853 1926
rect 842 1893 845 1923
rect 826 1873 837 1876
rect 858 1873 861 1936
rect 818 1823 821 1866
rect 834 1826 837 1873
rect 866 1836 869 1943
rect 826 1823 837 1826
rect 858 1833 869 1836
rect 826 1803 829 1823
rect 858 1813 861 1833
rect 810 1793 837 1796
rect 778 1693 789 1696
rect 786 1596 789 1693
rect 754 1593 765 1596
rect 742 1533 749 1536
rect 730 1503 733 1516
rect 746 1413 749 1533
rect 762 1476 765 1593
rect 778 1593 789 1596
rect 798 1693 805 1696
rect 810 1736 813 1766
rect 834 1736 837 1793
rect 810 1733 821 1736
rect 826 1733 837 1736
rect 770 1523 773 1536
rect 770 1483 773 1516
rect 762 1473 773 1476
rect 762 1413 765 1436
rect 674 1323 685 1326
rect 642 1173 645 1193
rect 674 1166 677 1216
rect 682 1193 685 1323
rect 698 1256 701 1336
rect 706 1326 709 1376
rect 714 1343 717 1356
rect 706 1323 717 1326
rect 694 1253 701 1256
rect 642 1163 677 1166
rect 594 1153 621 1156
rect 586 1056 589 1126
rect 594 1066 597 1136
rect 602 1123 605 1146
rect 618 1143 621 1153
rect 610 1123 613 1136
rect 642 1123 645 1163
rect 694 1156 697 1253
rect 714 1246 717 1323
rect 706 1243 717 1246
rect 706 1213 709 1243
rect 694 1153 701 1156
rect 674 1133 677 1146
rect 674 1086 677 1126
rect 698 1106 701 1153
rect 706 1123 709 1206
rect 730 1193 733 1326
rect 754 1266 757 1406
rect 770 1403 773 1473
rect 778 1386 781 1593
rect 798 1576 801 1693
rect 810 1603 813 1733
rect 826 1666 829 1733
rect 842 1703 845 1716
rect 826 1663 833 1666
rect 818 1623 821 1656
rect 798 1573 805 1576
rect 802 1546 805 1573
rect 786 1543 805 1546
rect 786 1503 789 1543
rect 818 1526 821 1616
rect 830 1606 833 1663
rect 850 1623 853 1636
rect 830 1603 845 1606
rect 834 1546 837 1603
rect 794 1523 821 1526
rect 830 1543 837 1546
rect 810 1503 813 1516
rect 786 1403 789 1426
rect 778 1383 785 1386
rect 770 1333 773 1356
rect 782 1326 785 1383
rect 778 1323 785 1326
rect 794 1323 797 1486
rect 802 1446 805 1466
rect 802 1443 809 1446
rect 806 1346 809 1443
rect 818 1396 821 1456
rect 830 1436 833 1543
rect 830 1433 837 1436
rect 826 1403 829 1416
rect 818 1393 829 1396
rect 834 1393 837 1433
rect 802 1343 809 1346
rect 802 1323 805 1343
rect 818 1326 821 1336
rect 826 1333 829 1393
rect 842 1346 845 1536
rect 850 1463 853 1596
rect 858 1533 861 1786
rect 866 1733 869 1826
rect 874 1693 877 2103
rect 914 2046 917 2163
rect 930 2123 933 2136
rect 938 2133 941 2156
rect 946 2123 949 2146
rect 962 2123 965 2203
rect 978 2153 981 2203
rect 986 2186 989 2206
rect 1010 2203 1021 2206
rect 986 2183 997 2186
rect 978 2133 981 2146
rect 978 2106 981 2126
rect 994 2106 997 2183
rect 1018 2123 1021 2203
rect 970 2103 981 2106
rect 986 2103 997 2106
rect 1018 2103 1021 2116
rect 914 2043 921 2046
rect 882 2013 893 2016
rect 882 1963 885 2006
rect 898 1936 901 2006
rect 906 2003 909 2026
rect 918 1986 921 2043
rect 918 1983 925 1986
rect 882 1853 885 1936
rect 890 1933 901 1936
rect 906 1963 917 1966
rect 890 1803 893 1933
rect 898 1813 901 1926
rect 906 1796 909 1963
rect 922 1946 925 1983
rect 890 1793 909 1796
rect 918 1943 925 1946
rect 890 1736 893 1793
rect 918 1736 921 1943
rect 886 1733 893 1736
rect 910 1733 921 1736
rect 866 1523 869 1586
rect 874 1533 877 1686
rect 886 1636 889 1733
rect 882 1633 889 1636
rect 882 1613 885 1633
rect 874 1493 877 1526
rect 850 1413 853 1436
rect 874 1413 885 1416
rect 834 1343 845 1346
rect 810 1323 821 1326
rect 754 1263 765 1266
rect 746 1233 757 1236
rect 746 1203 749 1233
rect 754 1193 757 1206
rect 762 1193 765 1263
rect 778 1246 781 1323
rect 774 1243 781 1246
rect 774 1146 777 1243
rect 786 1213 789 1236
rect 762 1126 765 1146
rect 774 1143 781 1146
rect 786 1143 789 1206
rect 698 1103 709 1106
rect 674 1083 685 1086
rect 594 1063 613 1066
rect 586 1053 605 1056
rect 570 1043 581 1046
rect 530 1013 541 1016
rect 546 1013 549 1026
rect 554 1023 573 1026
rect 530 993 533 1013
rect 554 1006 557 1023
rect 538 1003 557 1006
rect 538 933 541 966
rect 522 923 541 926
rect 514 913 525 916
rect 522 846 525 913
rect 538 906 541 923
rect 546 913 549 926
rect 554 906 557 936
rect 538 903 557 906
rect 522 843 533 846
rect 482 803 501 806
rect 482 746 485 803
rect 506 796 509 826
rect 506 793 513 796
rect 482 743 489 746
rect 426 606 429 616
rect 434 613 437 723
rect 450 703 453 716
rect 474 693 477 736
rect 486 686 489 743
rect 498 723 501 786
rect 510 736 513 793
rect 510 733 517 736
rect 522 733 525 746
rect 506 706 509 726
rect 482 683 489 686
rect 498 703 509 706
rect 466 613 469 626
rect 482 613 485 683
rect 498 626 501 703
rect 498 623 509 626
rect 426 603 453 606
rect 426 506 429 526
rect 426 503 433 506
rect 430 446 433 503
rect 426 443 433 446
rect 426 413 429 443
rect 442 423 445 536
rect 450 513 453 603
rect 458 563 461 606
rect 466 593 469 606
rect 482 603 501 606
rect 482 546 485 603
rect 506 593 509 623
rect 514 613 517 733
rect 530 726 533 843
rect 538 813 541 903
rect 562 893 565 1016
rect 570 1013 573 1023
rect 570 933 573 1006
rect 578 836 581 1043
rect 586 943 589 956
rect 594 916 597 1016
rect 554 833 581 836
rect 590 913 597 916
rect 554 783 557 833
rect 590 786 593 913
rect 590 783 597 786
rect 522 723 533 726
rect 522 586 525 723
rect 562 706 565 726
rect 570 713 573 736
rect 594 733 597 783
rect 554 703 565 706
rect 530 623 533 656
rect 554 636 557 703
rect 554 633 565 636
rect 562 613 565 633
rect 578 623 581 726
rect 586 703 589 726
rect 602 696 605 1053
rect 610 996 613 1063
rect 618 1023 677 1026
rect 618 1003 621 1023
rect 634 996 637 1006
rect 610 993 637 996
rect 610 943 613 956
rect 610 813 613 926
rect 618 876 621 966
rect 626 893 629 936
rect 634 933 637 993
rect 618 873 625 876
rect 622 806 625 873
rect 634 826 637 926
rect 658 836 661 1016
rect 674 1013 677 1023
rect 674 883 677 926
rect 682 916 685 1083
rect 706 986 709 1103
rect 754 1056 757 1126
rect 762 1123 769 1126
rect 766 1066 769 1123
rect 738 1053 757 1056
rect 762 1063 769 1066
rect 778 1066 781 1143
rect 778 1063 789 1066
rect 738 1013 741 1053
rect 762 1003 765 1063
rect 786 996 789 1063
rect 794 1013 797 1136
rect 802 1123 805 1226
rect 810 1203 813 1323
rect 826 1283 829 1326
rect 818 1213 829 1216
rect 834 1196 837 1343
rect 850 1246 853 1406
rect 874 1393 877 1406
rect 890 1333 893 1616
rect 898 1603 901 1716
rect 910 1596 913 1733
rect 906 1593 913 1596
rect 898 1523 901 1536
rect 898 1413 901 1426
rect 906 1373 909 1593
rect 922 1583 925 1726
rect 930 1716 933 2086
rect 970 2036 973 2103
rect 970 2033 981 2036
rect 938 1936 941 1996
rect 954 1963 957 2016
rect 962 1976 965 2016
rect 978 2003 981 2033
rect 986 1996 989 2103
rect 994 2023 997 2046
rect 1002 2003 1005 2026
rect 1010 2013 1013 2086
rect 978 1993 989 1996
rect 1026 1996 1029 2336
rect 1034 2253 1037 2363
rect 1042 2353 1077 2356
rect 1042 2323 1045 2353
rect 1050 2333 1053 2346
rect 1058 2293 1061 2326
rect 1050 2213 1053 2286
rect 1066 2206 1069 2336
rect 1074 2323 1077 2353
rect 1082 2253 1085 2336
rect 1090 2333 1093 2406
rect 1098 2376 1101 2423
rect 1106 2393 1109 2406
rect 1098 2373 1105 2376
rect 1102 2326 1105 2373
rect 1098 2323 1105 2326
rect 1050 2203 1069 2206
rect 1050 2196 1053 2203
rect 1082 2196 1085 2216
rect 1098 2213 1101 2323
rect 1114 2276 1117 2536
rect 1122 2513 1125 2526
rect 1138 2513 1141 2543
rect 1146 2523 1149 2546
rect 1170 2506 1173 2563
rect 1194 2513 1197 2576
rect 1210 2563 1253 2566
rect 1210 2533 1213 2563
rect 1170 2503 1181 2506
rect 1154 2423 1165 2426
rect 1138 2413 1165 2416
rect 1154 2396 1157 2406
rect 1138 2393 1157 2396
rect 1154 2373 1157 2393
rect 1162 2383 1165 2413
rect 1170 2366 1173 2426
rect 1154 2363 1173 2366
rect 1130 2283 1133 2326
rect 1138 2303 1141 2336
rect 1146 2293 1149 2326
rect 1154 2323 1157 2363
rect 1178 2306 1181 2503
rect 1202 2493 1205 2526
rect 1218 2503 1221 2526
rect 1234 2523 1237 2556
rect 1242 2506 1245 2536
rect 1250 2513 1253 2563
rect 1258 2533 1269 2536
rect 1274 2533 1277 2546
rect 1258 2523 1269 2526
rect 1242 2503 1253 2506
rect 1250 2466 1253 2503
rect 1258 2473 1261 2523
rect 1282 2466 1285 2556
rect 1250 2463 1285 2466
rect 1170 2303 1181 2306
rect 1114 2273 1149 2276
rect 1106 2203 1109 2216
rect 1034 2193 1053 2196
rect 1066 2193 1085 2196
rect 1034 2086 1037 2136
rect 1042 2103 1045 2126
rect 1034 2083 1045 2086
rect 1026 1993 1037 1996
rect 962 1973 969 1976
rect 938 1933 949 1936
rect 938 1733 941 1806
rect 946 1773 949 1866
rect 930 1713 937 1716
rect 934 1606 937 1713
rect 930 1603 937 1606
rect 914 1506 917 1536
rect 922 1523 925 1576
rect 914 1503 921 1506
rect 918 1436 921 1503
rect 930 1463 933 1603
rect 914 1433 921 1436
rect 914 1413 917 1433
rect 930 1393 933 1416
rect 898 1333 917 1336
rect 930 1333 933 1386
rect 842 1243 853 1246
rect 842 1203 845 1243
rect 850 1223 877 1226
rect 850 1213 853 1223
rect 858 1203 861 1216
rect 818 1193 837 1196
rect 818 1066 821 1193
rect 842 1173 845 1196
rect 850 1133 853 1146
rect 874 1123 877 1223
rect 890 1193 893 1206
rect 898 1166 901 1333
rect 906 1316 909 1326
rect 914 1323 917 1333
rect 906 1313 933 1316
rect 938 1306 941 1586
rect 946 1326 949 1766
rect 954 1723 957 1926
rect 966 1756 969 1973
rect 978 1793 981 1993
rect 986 1913 989 1926
rect 962 1753 969 1756
rect 962 1713 965 1753
rect 994 1746 997 1966
rect 1002 1923 1005 1946
rect 1026 1933 1029 1986
rect 1018 1913 1021 1926
rect 1034 1916 1037 1993
rect 1042 1986 1045 2083
rect 1066 2013 1069 2193
rect 1090 2136 1093 2196
rect 1130 2153 1133 2196
rect 1106 2143 1125 2146
rect 1090 2133 1097 2136
rect 1106 2133 1109 2143
rect 1122 2136 1125 2143
rect 1042 1983 1049 1986
rect 1046 1926 1049 1983
rect 1030 1913 1037 1916
rect 1042 1923 1049 1926
rect 1002 1813 1005 1826
rect 994 1743 1001 1746
rect 970 1656 973 1736
rect 954 1653 973 1656
rect 954 1593 957 1653
rect 970 1613 973 1646
rect 978 1613 981 1726
rect 986 1683 989 1736
rect 998 1676 1001 1743
rect 994 1673 1001 1676
rect 954 1523 957 1546
rect 962 1533 965 1606
rect 970 1516 973 1606
rect 978 1536 981 1606
rect 994 1603 997 1673
rect 978 1533 989 1536
rect 954 1513 973 1516
rect 954 1403 957 1513
rect 978 1503 981 1526
rect 962 1413 965 1446
rect 986 1423 989 1533
rect 994 1523 997 1596
rect 1002 1533 1005 1616
rect 1010 1593 1013 1906
rect 1030 1836 1033 1913
rect 1030 1833 1037 1836
rect 1018 1813 1021 1826
rect 1018 1723 1021 1806
rect 1026 1783 1029 1816
rect 1026 1733 1029 1746
rect 1026 1583 1029 1606
rect 994 1413 997 1456
rect 946 1323 957 1326
rect 978 1323 981 1336
rect 922 1303 941 1306
rect 922 1226 925 1303
rect 922 1223 929 1226
rect 914 1183 917 1216
rect 926 1176 929 1223
rect 946 1213 949 1316
rect 954 1306 957 1323
rect 954 1303 961 1306
rect 958 1236 961 1303
rect 986 1286 989 1406
rect 1002 1403 1005 1506
rect 1010 1473 1013 1536
rect 1018 1523 1021 1576
rect 1026 1516 1029 1546
rect 1022 1513 1029 1516
rect 1022 1466 1025 1513
rect 1034 1503 1037 1833
rect 1042 1763 1045 1923
rect 1050 1803 1053 1906
rect 1058 1876 1061 2006
rect 1074 1996 1077 2126
rect 1082 2093 1085 2126
rect 1094 2086 1097 2133
rect 1090 2083 1097 2086
rect 1090 2006 1093 2083
rect 1090 2003 1097 2006
rect 1066 1993 1077 1996
rect 1066 1896 1069 1993
rect 1074 1913 1077 1986
rect 1082 1973 1085 1996
rect 1094 1946 1097 2003
rect 1090 1943 1097 1946
rect 1066 1893 1077 1896
rect 1058 1873 1065 1876
rect 1062 1816 1065 1873
rect 1058 1813 1065 1816
rect 1042 1743 1045 1756
rect 1050 1733 1053 1786
rect 1058 1726 1061 1813
rect 1074 1796 1077 1893
rect 1090 1813 1093 1943
rect 1106 1923 1109 2126
rect 1114 2123 1117 2136
rect 1122 2133 1133 2136
rect 1138 2123 1141 2216
rect 1146 2116 1149 2273
rect 1170 2236 1173 2303
rect 1170 2233 1181 2236
rect 1154 2143 1157 2216
rect 1178 2206 1181 2233
rect 1186 2213 1189 2416
rect 1234 2413 1237 2446
rect 1250 2413 1253 2463
rect 1274 2446 1277 2463
rect 1290 2453 1293 2526
rect 1306 2453 1309 2536
rect 1330 2466 1333 2536
rect 1362 2516 1365 2536
rect 1314 2463 1333 2466
rect 1354 2513 1365 2516
rect 1314 2446 1317 2463
rect 1270 2443 1277 2446
rect 1282 2443 1317 2446
rect 1194 2353 1197 2406
rect 1258 2373 1261 2416
rect 1270 2396 1273 2443
rect 1282 2403 1285 2443
rect 1306 2403 1309 2436
rect 1330 2413 1333 2456
rect 1354 2426 1357 2513
rect 1354 2423 1365 2426
rect 1354 2396 1357 2406
rect 1270 2393 1277 2396
rect 1242 2336 1245 2346
rect 1202 2266 1205 2336
rect 1218 2333 1245 2336
rect 1226 2323 1237 2326
rect 1226 2273 1229 2323
rect 1202 2263 1253 2266
rect 1178 2203 1189 2206
rect 1162 2116 1165 2136
rect 1122 2113 1149 2116
rect 1158 2113 1165 2116
rect 1170 2133 1181 2136
rect 1122 1956 1125 2113
rect 1138 1993 1141 2016
rect 1146 2003 1149 2066
rect 1158 2046 1161 2113
rect 1158 2043 1165 2046
rect 1154 2003 1157 2026
rect 1162 2013 1165 2043
rect 1170 2036 1173 2133
rect 1186 2116 1189 2203
rect 1202 2126 1205 2206
rect 1210 2203 1213 2216
rect 1226 2213 1229 2226
rect 1218 2183 1221 2206
rect 1242 2156 1245 2206
rect 1250 2203 1253 2263
rect 1258 2216 1261 2336
rect 1274 2316 1277 2393
rect 1322 2393 1357 2396
rect 1282 2333 1285 2346
rect 1322 2323 1325 2393
rect 1330 2333 1341 2336
rect 1346 2333 1349 2346
rect 1274 2313 1285 2316
rect 1282 2216 1285 2313
rect 1330 2283 1333 2326
rect 1354 2293 1357 2326
rect 1258 2213 1265 2216
rect 1234 2133 1237 2156
rect 1242 2153 1253 2156
rect 1202 2123 1237 2126
rect 1178 2103 1181 2116
rect 1186 2113 1205 2116
rect 1170 2033 1181 2036
rect 1114 1953 1125 1956
rect 1066 1793 1077 1796
rect 1066 1736 1069 1793
rect 1090 1783 1093 1806
rect 1066 1733 1077 1736
rect 1058 1723 1069 1726
rect 1058 1696 1061 1716
rect 1050 1693 1061 1696
rect 1050 1636 1053 1693
rect 1050 1633 1061 1636
rect 1042 1613 1053 1616
rect 1058 1606 1061 1633
rect 1042 1586 1045 1606
rect 1050 1603 1061 1606
rect 1042 1583 1049 1586
rect 1046 1496 1049 1583
rect 1066 1546 1069 1723
rect 1074 1613 1077 1733
rect 1074 1583 1077 1606
rect 1082 1603 1085 1776
rect 1106 1726 1109 1806
rect 1114 1756 1117 1953
rect 1170 1946 1173 2033
rect 1122 1906 1125 1936
rect 1130 1916 1133 1936
rect 1138 1923 1141 1946
rect 1154 1943 1173 1946
rect 1130 1913 1141 1916
rect 1122 1903 1141 1906
rect 1122 1813 1125 1846
rect 1138 1826 1141 1903
rect 1154 1876 1157 1943
rect 1154 1873 1165 1876
rect 1162 1853 1165 1873
rect 1170 1856 1173 1936
rect 1186 1873 1189 1916
rect 1170 1853 1181 1856
rect 1178 1836 1181 1853
rect 1178 1833 1185 1836
rect 1134 1823 1141 1826
rect 1114 1753 1125 1756
rect 1114 1733 1117 1746
rect 1090 1706 1093 1726
rect 1098 1723 1109 1726
rect 1122 1713 1125 1753
rect 1134 1746 1137 1823
rect 1154 1816 1157 1826
rect 1146 1813 1157 1816
rect 1162 1813 1165 1826
rect 1146 1753 1149 1813
rect 1154 1783 1157 1806
rect 1170 1793 1173 1806
rect 1182 1766 1185 1833
rect 1178 1763 1185 1766
rect 1178 1746 1181 1763
rect 1194 1746 1197 1976
rect 1202 1763 1205 2113
rect 1234 2096 1237 2116
rect 1226 2093 1237 2096
rect 1226 2046 1229 2093
rect 1226 2043 1237 2046
rect 1234 2023 1237 2043
rect 1210 1946 1213 2016
rect 1234 1946 1237 2016
rect 1210 1943 1221 1946
rect 1226 1943 1237 1946
rect 1210 1813 1213 1936
rect 1218 1866 1221 1943
rect 1242 1926 1245 2146
rect 1250 1963 1253 2153
rect 1262 2086 1265 2213
rect 1258 2083 1265 2086
rect 1274 2213 1285 2216
rect 1306 2213 1309 2276
rect 1354 2246 1357 2266
rect 1346 2243 1357 2246
rect 1314 2213 1317 2226
rect 1258 2063 1261 2083
rect 1258 1973 1261 2006
rect 1274 1996 1277 2213
rect 1290 2153 1293 2196
rect 1306 2186 1309 2206
rect 1314 2196 1317 2206
rect 1330 2203 1333 2216
rect 1314 2193 1333 2196
rect 1306 2183 1325 2186
rect 1298 2083 1301 2136
rect 1306 2066 1309 2136
rect 1322 2133 1325 2183
rect 1330 2153 1333 2193
rect 1298 2063 1309 2066
rect 1282 2013 1285 2026
rect 1298 2016 1301 2063
rect 1298 2013 1309 2016
rect 1314 2013 1317 2126
rect 1330 2046 1333 2146
rect 1346 2056 1349 2243
rect 1362 2216 1365 2423
rect 1370 2413 1373 2526
rect 1378 2523 1381 2566
rect 1418 2543 1445 2546
rect 1370 2303 1373 2346
rect 1378 2293 1381 2416
rect 1386 2413 1389 2436
rect 1394 2353 1397 2516
rect 1358 2213 1365 2216
rect 1358 2146 1361 2213
rect 1378 2206 1381 2276
rect 1386 2223 1389 2236
rect 1370 2153 1373 2206
rect 1378 2203 1385 2206
rect 1358 2143 1365 2146
rect 1362 2066 1365 2143
rect 1382 2136 1385 2203
rect 1394 2143 1397 2336
rect 1382 2133 1397 2136
rect 1362 2063 1373 2066
rect 1346 2053 1365 2056
rect 1322 2043 1333 2046
rect 1274 1993 1285 1996
rect 1306 1993 1309 2013
rect 1226 1883 1229 1926
rect 1238 1923 1245 1926
rect 1250 1943 1269 1946
rect 1218 1863 1225 1866
rect 1222 1786 1225 1863
rect 1238 1826 1241 1923
rect 1238 1823 1245 1826
rect 1218 1783 1225 1786
rect 1134 1743 1141 1746
rect 1090 1703 1101 1706
rect 1098 1636 1101 1703
rect 1090 1633 1101 1636
rect 1090 1603 1093 1633
rect 1098 1556 1101 1616
rect 1018 1463 1025 1466
rect 1042 1493 1049 1496
rect 1058 1543 1069 1546
rect 1094 1553 1101 1556
rect 1010 1393 1013 1406
rect 994 1313 997 1326
rect 1002 1323 1005 1336
rect 1010 1293 1013 1336
rect 954 1233 961 1236
rect 970 1283 989 1286
rect 954 1206 957 1233
rect 938 1203 957 1206
rect 962 1186 965 1216
rect 970 1193 973 1283
rect 986 1186 989 1216
rect 1018 1213 1021 1463
rect 1042 1426 1045 1493
rect 1058 1466 1061 1543
rect 1066 1483 1069 1536
rect 1082 1503 1085 1536
rect 1094 1506 1097 1553
rect 1106 1513 1109 1546
rect 1094 1503 1101 1506
rect 1058 1463 1077 1466
rect 1034 1423 1045 1426
rect 1026 1333 1029 1366
rect 1026 1313 1029 1326
rect 1034 1296 1037 1423
rect 1074 1416 1077 1463
rect 1050 1376 1053 1416
rect 1058 1413 1069 1416
rect 1074 1413 1093 1416
rect 1042 1373 1053 1376
rect 1042 1333 1045 1373
rect 1050 1316 1053 1366
rect 1066 1333 1069 1406
rect 1074 1363 1077 1406
rect 1050 1313 1061 1316
rect 1074 1313 1077 1326
rect 1030 1293 1037 1296
rect 1030 1206 1033 1293
rect 962 1183 989 1186
rect 890 1163 901 1166
rect 922 1173 929 1176
rect 890 1086 893 1163
rect 890 1083 901 1086
rect 810 1063 821 1066
rect 810 1046 813 1063
rect 806 1043 813 1046
rect 698 983 709 986
rect 778 993 789 996
rect 698 963 701 983
rect 690 943 709 946
rect 690 923 693 943
rect 698 916 701 936
rect 706 933 709 943
rect 682 913 701 916
rect 706 913 709 926
rect 722 923 725 966
rect 730 896 733 946
rect 778 906 781 993
rect 806 986 809 1043
rect 890 1036 893 1056
rect 882 1033 893 1036
rect 806 983 813 986
rect 714 893 733 896
rect 770 903 781 906
rect 658 833 709 836
rect 634 823 661 826
rect 658 816 661 823
rect 618 803 625 806
rect 618 726 621 803
rect 586 693 605 696
rect 586 606 589 693
rect 498 583 525 586
rect 546 603 565 606
rect 582 603 589 606
rect 498 566 501 583
rect 474 543 485 546
rect 494 563 501 566
rect 474 456 477 543
rect 494 506 497 563
rect 546 536 549 603
rect 514 523 517 536
rect 546 533 553 536
rect 494 503 501 506
rect 498 486 501 503
rect 538 486 541 526
rect 498 483 525 486
rect 474 453 485 456
rect 442 403 445 416
rect 466 346 469 416
rect 458 343 469 346
rect 458 333 461 343
rect 482 336 485 453
rect 522 413 525 483
rect 534 483 541 486
rect 534 416 537 483
rect 550 476 553 533
rect 546 473 553 476
rect 534 413 541 416
rect 498 343 501 366
rect 466 333 485 336
rect 538 333 541 413
rect 546 333 549 473
rect 562 403 565 526
rect 582 506 585 603
rect 594 523 597 686
rect 610 656 613 726
rect 618 723 625 726
rect 602 653 613 656
rect 602 613 605 653
rect 622 636 625 723
rect 622 633 629 636
rect 610 613 621 616
rect 610 603 621 606
rect 626 593 629 633
rect 634 613 637 816
rect 658 813 693 816
rect 642 796 645 806
rect 666 803 677 806
rect 690 796 693 806
rect 642 793 693 796
rect 650 733 669 736
rect 642 613 645 726
rect 650 723 661 726
rect 666 693 669 733
rect 674 703 677 726
rect 682 613 685 786
rect 690 613 693 726
rect 698 723 701 826
rect 706 683 709 833
rect 698 603 701 636
rect 706 613 709 656
rect 714 603 717 893
rect 722 883 733 886
rect 722 783 725 816
rect 722 613 725 706
rect 634 523 637 536
rect 582 503 589 506
rect 586 486 589 503
rect 586 483 645 486
rect 586 343 589 416
rect 642 413 645 483
rect 666 436 669 486
rect 658 433 669 436
rect 658 386 661 433
rect 682 423 685 526
rect 730 523 733 883
rect 770 846 773 903
rect 770 843 781 846
rect 746 823 757 826
rect 754 813 757 823
rect 738 726 741 806
rect 762 746 765 826
rect 778 813 781 843
rect 786 823 789 946
rect 794 906 797 926
rect 802 913 805 966
rect 810 923 813 983
rect 794 903 805 906
rect 826 826 829 916
rect 842 913 845 1016
rect 858 933 861 986
rect 882 966 885 1033
rect 882 963 893 966
rect 882 933 885 946
rect 890 933 893 963
rect 898 933 901 1083
rect 922 993 925 1173
rect 994 1146 997 1206
rect 938 1126 941 1146
rect 962 1143 997 1146
rect 934 1123 941 1126
rect 934 1046 937 1123
rect 946 1053 949 1126
rect 934 1043 941 1046
rect 938 1003 941 1043
rect 970 1013 973 1136
rect 978 1123 981 1136
rect 1002 1056 1005 1206
rect 1030 1203 1037 1206
rect 1034 1186 1037 1203
rect 1042 1193 1045 1296
rect 1058 1236 1061 1313
rect 1082 1296 1085 1376
rect 1050 1233 1061 1236
rect 1074 1293 1085 1296
rect 1050 1203 1053 1233
rect 1058 1196 1061 1216
rect 1050 1193 1061 1196
rect 1034 1183 1045 1186
rect 1018 1133 1021 1146
rect 1042 1123 1045 1183
rect 1050 1116 1053 1193
rect 1074 1186 1077 1293
rect 1090 1276 1093 1413
rect 1098 1396 1101 1503
rect 1114 1436 1117 1626
rect 1138 1623 1141 1743
rect 1162 1713 1165 1746
rect 1170 1743 1189 1746
rect 1194 1743 1201 1746
rect 1170 1733 1173 1743
rect 1178 1733 1181 1743
rect 1186 1733 1189 1743
rect 1122 1523 1125 1546
rect 1138 1523 1141 1606
rect 1162 1603 1165 1616
rect 1170 1613 1173 1726
rect 1178 1626 1181 1676
rect 1186 1633 1189 1716
rect 1198 1636 1201 1743
rect 1218 1723 1221 1783
rect 1226 1683 1229 1726
rect 1194 1633 1201 1636
rect 1178 1623 1189 1626
rect 1122 1476 1125 1516
rect 1162 1506 1165 1556
rect 1170 1523 1173 1546
rect 1146 1503 1165 1506
rect 1170 1503 1173 1516
rect 1122 1473 1133 1476
rect 1106 1433 1117 1436
rect 1106 1413 1109 1433
rect 1098 1393 1105 1396
rect 1086 1273 1093 1276
rect 1086 1216 1089 1273
rect 1102 1266 1105 1393
rect 1098 1263 1105 1266
rect 1086 1213 1093 1216
rect 1098 1213 1101 1263
rect 1090 1193 1093 1213
rect 1098 1203 1109 1206
rect 1074 1183 1085 1186
rect 1082 1166 1085 1183
rect 1082 1163 1093 1166
rect 1042 1113 1053 1116
rect 1002 1053 1009 1056
rect 1006 1006 1009 1053
rect 1002 1003 1009 1006
rect 810 823 829 826
rect 794 813 845 816
rect 770 803 789 806
rect 746 743 765 746
rect 754 733 781 736
rect 738 723 765 726
rect 738 523 741 666
rect 746 596 749 686
rect 754 613 757 696
rect 778 636 781 733
rect 794 723 797 813
rect 826 803 837 806
rect 810 733 813 746
rect 818 716 821 736
rect 858 733 861 926
rect 874 916 877 926
rect 914 916 917 936
rect 938 933 941 986
rect 954 936 957 996
rect 950 933 957 936
rect 874 913 917 916
rect 922 876 925 926
rect 914 873 925 876
rect 874 813 893 816
rect 866 803 877 806
rect 866 733 869 766
rect 874 733 877 803
rect 810 713 821 716
rect 826 713 829 726
rect 810 646 813 713
rect 834 693 837 716
rect 810 643 821 646
rect 778 633 797 636
rect 818 626 821 643
rect 762 623 821 626
rect 762 603 765 623
rect 746 593 753 596
rect 750 516 753 593
rect 770 536 773 616
rect 778 603 781 616
rect 794 603 797 623
rect 802 603 805 616
rect 762 523 765 536
rect 770 533 781 536
rect 778 516 781 533
rect 750 513 765 516
rect 778 513 789 516
rect 754 456 757 476
rect 750 453 757 456
rect 682 403 685 416
rect 658 383 669 386
rect 602 343 605 366
rect 666 333 669 383
rect 690 343 693 366
rect 730 356 733 416
rect 750 406 753 453
rect 762 413 765 513
rect 794 483 797 536
rect 802 523 805 536
rect 826 523 829 676
rect 858 626 861 726
rect 858 623 869 626
rect 842 583 845 616
rect 850 593 853 606
rect 850 473 853 536
rect 866 513 869 623
rect 874 613 877 726
rect 874 523 877 536
rect 882 523 885 766
rect 890 726 893 806
rect 898 793 901 826
rect 914 816 917 873
rect 906 813 917 816
rect 890 723 897 726
rect 894 656 897 723
rect 906 716 909 813
rect 914 736 917 806
rect 914 733 925 736
rect 922 723 925 733
rect 906 713 917 716
rect 890 653 897 656
rect 914 656 917 713
rect 914 653 925 656
rect 890 603 893 653
rect 898 613 901 636
rect 914 613 917 626
rect 922 603 925 653
rect 930 603 933 926
rect 938 823 941 856
rect 950 826 953 933
rect 962 826 965 926
rect 970 906 973 926
rect 986 923 989 956
rect 994 933 997 946
rect 970 903 981 906
rect 950 823 957 826
rect 962 823 973 826
rect 938 713 941 816
rect 946 713 949 806
rect 954 803 957 823
rect 978 756 981 903
rect 1002 823 1005 1003
rect 1018 996 1021 1016
rect 1018 993 1029 996
rect 1010 933 1013 986
rect 1026 946 1029 993
rect 1042 986 1045 1113
rect 1058 1003 1061 1146
rect 1090 1086 1093 1163
rect 1106 1143 1109 1203
rect 1114 1193 1117 1426
rect 1122 1413 1125 1466
rect 1130 1413 1133 1473
rect 1130 1383 1133 1406
rect 1146 1403 1149 1476
rect 1162 1426 1165 1486
rect 1158 1423 1165 1426
rect 1122 1333 1125 1366
rect 1158 1356 1161 1423
rect 1158 1353 1165 1356
rect 1130 1333 1133 1346
rect 1146 1333 1157 1336
rect 1138 1303 1141 1326
rect 1122 1213 1141 1216
rect 1122 1183 1125 1213
rect 1130 1136 1133 1206
rect 1138 1163 1141 1213
rect 1146 1183 1149 1333
rect 1154 1283 1157 1316
rect 1162 1213 1165 1353
rect 1170 1293 1173 1416
rect 1170 1203 1173 1286
rect 1082 1083 1093 1086
rect 1106 1133 1133 1136
rect 1082 1013 1085 1083
rect 1106 1056 1109 1133
rect 1122 1106 1125 1126
rect 1122 1103 1133 1106
rect 1098 1053 1109 1056
rect 1042 983 1049 986
rect 1018 943 1029 946
rect 1018 923 1021 943
rect 1046 926 1049 983
rect 1010 823 1013 836
rect 970 753 981 756
rect 938 613 941 706
rect 954 606 957 736
rect 962 733 965 746
rect 970 616 973 753
rect 978 743 1005 746
rect 978 703 981 743
rect 938 603 957 606
rect 966 613 973 616
rect 906 513 909 586
rect 966 556 969 613
rect 966 553 973 556
rect 890 433 901 436
rect 750 403 757 406
rect 770 403 773 426
rect 730 353 741 356
rect 738 333 741 353
rect 754 333 757 403
rect 770 363 773 396
rect 802 393 805 406
rect 834 346 837 406
rect 834 343 841 346
rect 434 213 437 326
rect 474 313 485 316
rect 346 203 357 206
rect 290 193 349 196
rect 266 133 269 146
rect 314 123 317 176
rect 346 123 349 193
rect 354 143 357 203
rect 362 173 365 206
rect 418 176 421 206
rect 442 203 445 226
rect 490 223 493 326
rect 546 223 549 326
rect 562 313 573 316
rect 594 296 597 326
rect 594 293 605 296
rect 602 223 605 293
rect 642 213 645 326
rect 674 313 685 316
rect 690 223 693 326
rect 746 216 749 326
rect 770 223 773 326
rect 778 313 781 326
rect 810 226 813 336
rect 838 296 841 343
rect 850 323 853 426
rect 890 413 893 426
rect 898 413 901 433
rect 914 406 917 536
rect 946 513 949 536
rect 970 533 973 553
rect 970 433 973 526
rect 978 523 981 606
rect 986 596 989 736
rect 994 733 997 743
rect 994 703 997 726
rect 1002 693 1005 726
rect 1010 686 1013 776
rect 994 683 1013 686
rect 994 613 997 683
rect 1002 623 1013 626
rect 986 593 993 596
rect 990 506 993 593
rect 1010 566 1013 606
rect 1018 593 1021 826
rect 1034 816 1037 926
rect 1046 923 1053 926
rect 1058 923 1061 996
rect 1066 933 1069 946
rect 1030 813 1037 816
rect 1030 716 1033 813
rect 1030 713 1037 716
rect 1026 603 1029 696
rect 1034 643 1037 713
rect 1042 633 1045 806
rect 1050 683 1053 923
rect 1098 916 1101 1053
rect 1130 1046 1133 1103
rect 1126 1043 1133 1046
rect 1126 976 1129 1043
rect 1122 973 1129 976
rect 1122 923 1125 973
rect 1138 953 1141 1016
rect 1154 1003 1157 1146
rect 1162 1123 1165 1136
rect 1178 986 1181 1606
rect 1186 1553 1189 1623
rect 1186 1423 1189 1546
rect 1186 1213 1189 1386
rect 1194 1206 1197 1633
rect 1202 1543 1205 1616
rect 1210 1523 1213 1676
rect 1218 1603 1221 1656
rect 1234 1633 1237 1806
rect 1242 1796 1245 1823
rect 1250 1813 1253 1943
rect 1258 1916 1261 1936
rect 1266 1933 1269 1943
rect 1258 1913 1269 1916
rect 1266 1846 1269 1913
rect 1258 1843 1269 1846
rect 1242 1793 1249 1796
rect 1218 1593 1229 1596
rect 1226 1583 1229 1593
rect 1234 1576 1237 1616
rect 1246 1606 1249 1793
rect 1258 1743 1261 1843
rect 1266 1823 1293 1826
rect 1290 1813 1293 1823
rect 1258 1623 1261 1736
rect 1266 1633 1269 1806
rect 1282 1783 1285 1806
rect 1246 1603 1269 1606
rect 1274 1603 1277 1726
rect 1282 1693 1285 1706
rect 1226 1573 1237 1576
rect 1202 1503 1205 1516
rect 1202 1476 1205 1496
rect 1226 1483 1229 1573
rect 1234 1533 1237 1566
rect 1266 1543 1269 1603
rect 1274 1543 1277 1596
rect 1250 1516 1253 1536
rect 1250 1513 1257 1516
rect 1202 1473 1213 1476
rect 1210 1426 1213 1473
rect 1202 1423 1213 1426
rect 1202 1223 1205 1423
rect 1226 1413 1229 1476
rect 1242 1403 1245 1506
rect 1254 1396 1257 1513
rect 1266 1493 1269 1526
rect 1274 1503 1277 1536
rect 1250 1393 1257 1396
rect 1226 1333 1229 1366
rect 1210 1303 1213 1326
rect 1226 1323 1237 1326
rect 1226 1283 1229 1323
rect 1242 1316 1245 1326
rect 1234 1313 1245 1316
rect 1202 1213 1221 1216
rect 1218 1206 1221 1213
rect 1186 1193 1189 1206
rect 1194 1203 1213 1206
rect 1218 1203 1229 1206
rect 1194 1183 1197 1196
rect 1202 1013 1205 1126
rect 1210 1106 1213 1203
rect 1226 1173 1229 1196
rect 1234 1193 1237 1313
rect 1250 1226 1253 1393
rect 1266 1376 1269 1406
rect 1262 1373 1269 1376
rect 1262 1286 1265 1373
rect 1274 1333 1277 1456
rect 1282 1403 1285 1656
rect 1290 1583 1293 1796
rect 1298 1523 1301 1966
rect 1314 1903 1317 1916
rect 1322 1883 1325 2043
rect 1306 1823 1325 1826
rect 1306 1813 1309 1823
rect 1306 1753 1309 1806
rect 1314 1733 1317 1816
rect 1322 1793 1325 1823
rect 1330 1726 1333 2006
rect 1338 1993 1341 2026
rect 1354 1973 1357 2026
rect 1362 2013 1365 2053
rect 1370 2003 1373 2063
rect 1338 1903 1341 1926
rect 1346 1923 1357 1926
rect 1338 1856 1341 1876
rect 1338 1853 1345 1856
rect 1342 1766 1345 1853
rect 1354 1803 1357 1816
rect 1362 1793 1365 1996
rect 1370 1883 1373 1926
rect 1378 1873 1381 2106
rect 1386 2093 1389 2126
rect 1378 1823 1381 1866
rect 1386 1786 1389 2086
rect 1394 1873 1397 2133
rect 1402 1966 1405 2536
rect 1418 2533 1421 2543
rect 1426 2473 1429 2526
rect 1434 2503 1437 2536
rect 1442 2533 1445 2543
rect 1474 2533 1493 2536
rect 1506 2533 1509 2556
rect 1410 2403 1413 2456
rect 1410 2333 1413 2366
rect 1418 2306 1421 2426
rect 1434 2346 1437 2416
rect 1442 2403 1453 2406
rect 1450 2373 1453 2403
rect 1458 2383 1461 2516
rect 1474 2423 1477 2516
rect 1482 2513 1485 2526
rect 1434 2343 1469 2346
rect 1474 2343 1477 2416
rect 1482 2403 1485 2436
rect 1490 2426 1493 2533
rect 1538 2526 1541 2546
rect 1546 2533 1549 2546
rect 1498 2473 1501 2526
rect 1506 2523 1541 2526
rect 1506 2493 1509 2523
rect 1522 2426 1525 2456
rect 1546 2446 1549 2516
rect 1554 2503 1557 2536
rect 1586 2533 1589 2556
rect 1570 2466 1573 2526
rect 1578 2493 1581 2526
rect 1602 2473 1605 2536
rect 1570 2463 1597 2466
rect 1546 2443 1565 2446
rect 1490 2423 1525 2426
rect 1554 2416 1557 2436
rect 1530 2413 1557 2416
rect 1530 2406 1533 2413
rect 1506 2403 1533 2406
rect 1490 2343 1533 2346
rect 1410 2303 1421 2306
rect 1426 2303 1429 2326
rect 1410 2153 1413 2303
rect 1418 2223 1421 2296
rect 1418 2136 1421 2216
rect 1434 2143 1437 2336
rect 1442 2293 1445 2326
rect 1450 2323 1453 2336
rect 1450 2213 1453 2286
rect 1410 2133 1421 2136
rect 1410 2093 1413 2133
rect 1418 2083 1421 2126
rect 1410 1983 1413 2016
rect 1418 1986 1421 2076
rect 1426 2023 1429 2126
rect 1442 2096 1445 2136
rect 1450 2113 1453 2146
rect 1442 2093 1449 2096
rect 1434 2016 1437 2056
rect 1446 2036 1449 2093
rect 1446 2033 1453 2036
rect 1426 1993 1429 2016
rect 1434 2013 1445 2016
rect 1434 1986 1437 2006
rect 1418 1983 1437 1986
rect 1402 1963 1409 1966
rect 1406 1866 1409 1963
rect 1306 1723 1333 1726
rect 1338 1763 1345 1766
rect 1362 1783 1389 1786
rect 1402 1863 1409 1866
rect 1306 1516 1309 1723
rect 1314 1696 1317 1716
rect 1314 1693 1321 1696
rect 1318 1626 1321 1693
rect 1338 1656 1341 1763
rect 1346 1733 1349 1746
rect 1314 1623 1321 1626
rect 1330 1653 1341 1656
rect 1314 1603 1317 1623
rect 1314 1576 1317 1596
rect 1314 1573 1321 1576
rect 1290 1513 1309 1516
rect 1274 1293 1277 1326
rect 1290 1306 1293 1513
rect 1318 1506 1321 1573
rect 1298 1413 1301 1506
rect 1314 1503 1321 1506
rect 1330 1526 1333 1653
rect 1338 1536 1341 1606
rect 1354 1593 1357 1636
rect 1362 1606 1365 1783
rect 1370 1723 1381 1726
rect 1370 1713 1373 1723
rect 1386 1646 1389 1736
rect 1402 1653 1405 1863
rect 1418 1823 1421 1976
rect 1434 1886 1437 1976
rect 1442 1933 1445 1946
rect 1450 1943 1453 2033
rect 1426 1883 1437 1886
rect 1426 1816 1429 1883
rect 1418 1813 1429 1816
rect 1418 1743 1421 1813
rect 1426 1723 1429 1806
rect 1386 1643 1397 1646
rect 1370 1613 1373 1636
rect 1362 1603 1373 1606
rect 1378 1603 1381 1626
rect 1370 1546 1373 1603
rect 1370 1543 1377 1546
rect 1338 1533 1349 1536
rect 1330 1523 1349 1526
rect 1314 1406 1317 1503
rect 1298 1393 1301 1406
rect 1314 1403 1325 1406
rect 1298 1333 1309 1336
rect 1314 1316 1317 1386
rect 1322 1333 1325 1403
rect 1330 1376 1333 1523
rect 1346 1493 1349 1516
rect 1362 1476 1365 1536
rect 1374 1486 1377 1543
rect 1386 1533 1389 1616
rect 1394 1613 1397 1643
rect 1402 1623 1429 1626
rect 1402 1603 1405 1623
rect 1410 1543 1413 1606
rect 1418 1526 1421 1546
rect 1414 1523 1421 1526
rect 1354 1473 1365 1476
rect 1370 1483 1377 1486
rect 1338 1383 1341 1416
rect 1354 1396 1357 1473
rect 1370 1463 1373 1483
rect 1354 1393 1365 1396
rect 1330 1373 1349 1376
rect 1330 1333 1341 1336
rect 1346 1326 1349 1373
rect 1338 1323 1349 1326
rect 1314 1313 1325 1316
rect 1354 1313 1357 1326
rect 1290 1303 1317 1306
rect 1262 1283 1269 1286
rect 1246 1223 1253 1226
rect 1266 1226 1269 1283
rect 1314 1236 1317 1303
rect 1362 1296 1365 1393
rect 1370 1366 1373 1426
rect 1378 1373 1381 1416
rect 1386 1413 1389 1426
rect 1402 1413 1405 1506
rect 1414 1456 1417 1523
rect 1414 1453 1421 1456
rect 1370 1363 1381 1366
rect 1370 1333 1373 1356
rect 1378 1326 1381 1363
rect 1386 1346 1389 1406
rect 1394 1393 1397 1406
rect 1410 1403 1413 1436
rect 1418 1426 1421 1453
rect 1426 1446 1429 1616
rect 1434 1453 1437 1876
rect 1442 1816 1445 1866
rect 1458 1826 1461 2236
rect 1466 2096 1469 2343
rect 1482 2316 1485 2336
rect 1478 2313 1485 2316
rect 1478 2246 1481 2313
rect 1478 2243 1485 2246
rect 1474 2113 1477 2226
rect 1482 2123 1485 2243
rect 1466 2093 1477 2096
rect 1474 2036 1477 2093
rect 1466 2033 1477 2036
rect 1466 1986 1469 2033
rect 1490 2016 1493 2343
rect 1538 2336 1541 2406
rect 1506 2333 1541 2336
rect 1506 2253 1509 2326
rect 1538 2316 1541 2333
rect 1522 2293 1525 2316
rect 1534 2313 1541 2316
rect 1534 2266 1537 2313
rect 1546 2273 1549 2336
rect 1562 2316 1565 2443
rect 1570 2373 1573 2416
rect 1578 2403 1581 2456
rect 1586 2413 1589 2446
rect 1578 2323 1581 2386
rect 1562 2313 1573 2316
rect 1534 2263 1541 2266
rect 1506 2223 1517 2226
rect 1498 2116 1501 2206
rect 1530 2123 1533 2216
rect 1498 2113 1509 2116
rect 1506 2026 1509 2113
rect 1530 2103 1533 2116
rect 1506 2023 1533 2026
rect 1482 2013 1501 2016
rect 1482 1993 1485 2013
rect 1466 1983 1485 1986
rect 1474 1906 1477 1926
rect 1470 1903 1477 1906
rect 1470 1846 1473 1903
rect 1470 1843 1477 1846
rect 1458 1823 1469 1826
rect 1442 1813 1461 1816
rect 1442 1783 1445 1806
rect 1466 1796 1469 1823
rect 1474 1813 1477 1843
rect 1482 1806 1485 1983
rect 1490 1976 1493 2006
rect 1498 1993 1501 2013
rect 1506 1993 1509 2016
rect 1490 1973 1497 1976
rect 1462 1793 1469 1796
rect 1474 1803 1485 1806
rect 1494 1806 1497 1973
rect 1514 1963 1517 2006
rect 1522 1956 1525 2016
rect 1506 1953 1525 1956
rect 1506 1813 1509 1953
rect 1514 1936 1517 1946
rect 1514 1933 1525 1936
rect 1530 1916 1533 2023
rect 1538 1993 1541 2263
rect 1570 2236 1573 2313
rect 1586 2303 1589 2346
rect 1570 2233 1581 2236
rect 1546 2213 1557 2216
rect 1554 2193 1557 2206
rect 1562 2203 1565 2216
rect 1570 2173 1573 2206
rect 1578 2166 1581 2233
rect 1586 2196 1589 2216
rect 1594 2213 1597 2463
rect 1610 2386 1613 2576
rect 1618 2526 1621 2536
rect 1626 2533 1629 2556
rect 1650 2533 1653 2556
rect 1618 2523 1629 2526
rect 1626 2513 1629 2523
rect 1666 2503 1669 2546
rect 1698 2513 1701 2536
rect 1706 2533 1709 2546
rect 1738 2543 1741 2586
rect 1730 2533 1741 2536
rect 1730 2526 1733 2533
rect 1706 2503 1709 2526
rect 1714 2523 1733 2526
rect 1618 2403 1621 2436
rect 1610 2383 1621 2386
rect 1618 2326 1621 2383
rect 1602 2256 1605 2326
rect 1610 2323 1621 2326
rect 1610 2303 1613 2323
rect 1642 2256 1645 2406
rect 1658 2346 1661 2416
rect 1666 2396 1669 2486
rect 1690 2423 1693 2446
rect 1674 2403 1693 2406
rect 1666 2393 1677 2396
rect 1698 2393 1701 2466
rect 1602 2253 1613 2256
rect 1586 2193 1593 2196
rect 1546 2163 1581 2166
rect 1546 2116 1549 2163
rect 1570 2133 1573 2146
rect 1578 2133 1581 2156
rect 1546 2113 1553 2116
rect 1550 2046 1553 2113
rect 1546 2043 1553 2046
rect 1546 1973 1549 2043
rect 1554 2013 1557 2026
rect 1522 1913 1533 1916
rect 1522 1836 1525 1913
rect 1522 1833 1533 1836
rect 1494 1803 1501 1806
rect 1450 1733 1453 1766
rect 1462 1726 1465 1793
rect 1474 1736 1477 1803
rect 1482 1793 1493 1796
rect 1498 1746 1501 1803
rect 1522 1796 1525 1816
rect 1530 1813 1533 1833
rect 1538 1813 1541 1926
rect 1546 1883 1549 1926
rect 1554 1836 1557 1946
rect 1546 1833 1557 1836
rect 1546 1823 1549 1833
rect 1554 1813 1557 1826
rect 1538 1803 1557 1806
rect 1498 1743 1505 1746
rect 1474 1733 1485 1736
rect 1442 1563 1445 1716
rect 1450 1706 1453 1726
rect 1462 1723 1469 1726
rect 1450 1703 1457 1706
rect 1454 1576 1457 1703
rect 1466 1613 1469 1723
rect 1474 1653 1477 1726
rect 1466 1583 1469 1606
rect 1450 1573 1457 1576
rect 1450 1556 1453 1573
rect 1474 1563 1477 1616
rect 1442 1553 1453 1556
rect 1426 1443 1437 1446
rect 1418 1423 1429 1426
rect 1386 1343 1397 1346
rect 1354 1293 1365 1296
rect 1370 1323 1381 1326
rect 1314 1233 1325 1236
rect 1266 1223 1309 1226
rect 1246 1156 1249 1223
rect 1246 1153 1253 1156
rect 1226 1133 1229 1146
rect 1210 1103 1229 1106
rect 1178 983 1193 986
rect 1138 933 1141 946
rect 1146 933 1157 936
rect 1162 933 1165 956
rect 1098 913 1109 916
rect 1066 813 1069 826
rect 1074 763 1077 856
rect 1098 806 1101 866
rect 1106 856 1109 913
rect 1106 853 1125 856
rect 1106 813 1109 853
rect 1098 803 1109 806
rect 1082 733 1085 756
rect 1090 733 1093 746
rect 1058 723 1077 726
rect 1074 703 1077 716
rect 1098 673 1101 803
rect 1122 796 1125 846
rect 1106 793 1125 796
rect 1106 636 1109 793
rect 1130 776 1133 926
rect 1146 913 1149 926
rect 1170 913 1173 936
rect 1178 903 1181 926
rect 1138 783 1141 836
rect 1146 793 1149 826
rect 1162 806 1165 836
rect 1170 823 1173 846
rect 1190 806 1193 983
rect 1202 886 1205 946
rect 1226 936 1229 1103
rect 1250 953 1253 1153
rect 1258 1123 1261 1216
rect 1274 1193 1277 1216
rect 1298 1163 1301 1206
rect 1306 1193 1309 1223
rect 1322 1166 1325 1233
rect 1354 1226 1357 1293
rect 1370 1263 1373 1323
rect 1354 1223 1365 1226
rect 1346 1203 1357 1206
rect 1314 1163 1325 1166
rect 1314 1143 1317 1163
rect 1354 1143 1357 1203
rect 1362 1193 1365 1223
rect 1378 1163 1381 1316
rect 1386 1213 1389 1336
rect 1394 1286 1397 1343
rect 1418 1333 1421 1356
rect 1426 1343 1429 1423
rect 1434 1403 1437 1443
rect 1410 1293 1413 1326
rect 1426 1286 1429 1326
rect 1434 1323 1437 1336
rect 1394 1283 1429 1286
rect 1434 1223 1437 1296
rect 1394 1203 1397 1216
rect 1426 1213 1437 1216
rect 1426 1196 1429 1213
rect 1418 1193 1429 1196
rect 1306 1026 1309 1126
rect 1338 1036 1341 1136
rect 1354 1126 1357 1136
rect 1354 1123 1381 1126
rect 1266 1023 1309 1026
rect 1330 1033 1341 1036
rect 1258 936 1261 976
rect 1222 933 1229 936
rect 1242 933 1261 936
rect 1202 883 1213 886
rect 1162 803 1181 806
rect 1190 803 1197 806
rect 1126 773 1133 776
rect 1178 773 1181 796
rect 1114 713 1117 726
rect 1126 666 1129 773
rect 1138 726 1141 746
rect 1170 743 1181 746
rect 1170 726 1173 743
rect 1186 733 1189 756
rect 1138 723 1149 726
rect 1146 676 1149 723
rect 1138 673 1149 676
rect 1162 723 1173 726
rect 1126 663 1133 666
rect 1074 633 1109 636
rect 1074 603 1077 633
rect 1098 593 1101 626
rect 1122 566 1125 646
rect 1130 606 1133 663
rect 1138 653 1141 673
rect 1130 603 1141 606
rect 1010 563 1017 566
rect 1122 563 1129 566
rect 990 503 997 506
rect 890 403 917 406
rect 898 323 901 396
rect 922 356 925 426
rect 970 413 973 426
rect 914 353 925 356
rect 914 323 917 353
rect 778 223 813 226
rect 834 293 841 296
rect 746 213 757 216
rect 418 173 469 176
rect 386 133 389 146
rect 434 123 437 156
rect 466 123 469 173
rect 482 153 485 206
rect 530 173 533 206
rect 578 203 589 206
rect 602 196 605 206
rect 562 193 605 196
rect 514 133 517 146
rect 562 123 565 193
rect 594 123 597 176
rect 626 163 629 206
rect 634 203 645 206
rect 690 166 693 206
rect 706 193 709 206
rect 682 163 693 166
rect 634 133 637 146
rect 682 123 685 163
rect 714 123 717 166
rect 746 113 749 136
rect 754 123 757 213
rect 778 133 781 223
rect 810 123 813 206
rect 834 203 837 293
rect 858 203 861 316
rect 906 183 909 216
rect 930 133 933 336
rect 954 226 957 406
rect 986 366 989 406
rect 994 386 997 503
rect 1014 486 1017 563
rect 1026 523 1029 536
rect 1010 483 1017 486
rect 1010 403 1013 483
rect 994 383 1005 386
rect 978 363 989 366
rect 978 323 981 363
rect 1002 286 1005 383
rect 1026 323 1029 426
rect 1034 413 1037 426
rect 1034 386 1037 406
rect 1042 403 1045 436
rect 1034 383 1041 386
rect 1050 383 1053 396
rect 1038 316 1041 383
rect 946 223 957 226
rect 994 283 1005 286
rect 1034 313 1041 316
rect 1058 313 1061 536
rect 1066 413 1069 426
rect 1090 403 1093 526
rect 1126 516 1129 563
rect 1138 523 1141 603
rect 1146 533 1149 616
rect 1154 603 1157 616
rect 1162 593 1165 723
rect 1178 626 1181 726
rect 1194 723 1197 803
rect 1202 663 1205 876
rect 1210 803 1213 883
rect 1222 866 1225 933
rect 1234 876 1237 926
rect 1242 896 1245 933
rect 1250 916 1253 926
rect 1266 923 1269 1023
rect 1274 976 1277 1016
rect 1274 973 1293 976
rect 1290 956 1293 973
rect 1274 916 1277 926
rect 1250 913 1277 916
rect 1282 896 1285 956
rect 1290 953 1297 956
rect 1242 893 1269 896
rect 1234 873 1245 876
rect 1222 863 1229 866
rect 1178 623 1205 626
rect 1170 546 1173 616
rect 1178 573 1181 606
rect 1186 593 1189 606
rect 1202 596 1205 623
rect 1210 613 1213 796
rect 1218 713 1221 816
rect 1226 723 1229 863
rect 1242 796 1245 873
rect 1258 813 1261 866
rect 1266 806 1269 893
rect 1278 893 1285 896
rect 1278 826 1281 893
rect 1294 886 1297 953
rect 1314 933 1317 1016
rect 1330 986 1333 1033
rect 1354 1003 1357 1016
rect 1386 1013 1389 1136
rect 1418 1123 1421 1193
rect 1434 1026 1437 1136
rect 1442 1133 1445 1553
rect 1450 1533 1453 1546
rect 1450 1473 1453 1526
rect 1458 1423 1461 1536
rect 1466 1493 1469 1526
rect 1450 1406 1453 1416
rect 1450 1403 1461 1406
rect 1466 1403 1469 1416
rect 1458 1396 1461 1403
rect 1474 1396 1477 1536
rect 1450 1363 1453 1396
rect 1458 1393 1477 1396
rect 1482 1393 1485 1733
rect 1490 1673 1493 1736
rect 1502 1656 1505 1743
rect 1498 1653 1505 1656
rect 1490 1603 1493 1626
rect 1490 1543 1493 1566
rect 1490 1523 1493 1536
rect 1498 1533 1501 1653
rect 1506 1613 1509 1636
rect 1514 1613 1517 1796
rect 1522 1793 1529 1796
rect 1526 1706 1529 1793
rect 1538 1726 1541 1756
rect 1546 1733 1549 1746
rect 1554 1736 1557 1803
rect 1562 1753 1565 2126
rect 1570 2123 1581 2126
rect 1590 2116 1593 2193
rect 1586 2113 1593 2116
rect 1570 1953 1573 2016
rect 1586 2013 1589 2113
rect 1602 2013 1605 2246
rect 1610 2223 1613 2253
rect 1618 2253 1645 2256
rect 1654 2343 1661 2346
rect 1610 2186 1613 2216
rect 1618 2196 1621 2253
rect 1642 2236 1645 2246
rect 1626 2233 1645 2236
rect 1654 2236 1657 2343
rect 1666 2253 1669 2336
rect 1674 2323 1677 2393
rect 1706 2373 1709 2416
rect 1714 2346 1717 2476
rect 1722 2413 1733 2416
rect 1682 2343 1717 2346
rect 1654 2233 1661 2236
rect 1626 2213 1629 2233
rect 1634 2213 1637 2226
rect 1642 2223 1645 2233
rect 1626 2203 1637 2206
rect 1618 2193 1629 2196
rect 1610 2183 1617 2186
rect 1614 2086 1617 2183
rect 1614 2083 1621 2086
rect 1610 2013 1613 2066
rect 1594 1973 1597 2006
rect 1570 1933 1589 1936
rect 1602 1933 1605 1956
rect 1586 1916 1589 1933
rect 1610 1916 1613 2006
rect 1586 1913 1597 1916
rect 1570 1813 1573 1846
rect 1570 1796 1573 1806
rect 1578 1796 1581 1886
rect 1594 1846 1597 1913
rect 1586 1843 1597 1846
rect 1606 1913 1613 1916
rect 1606 1846 1609 1913
rect 1606 1843 1613 1846
rect 1586 1816 1589 1843
rect 1586 1813 1597 1816
rect 1594 1803 1597 1813
rect 1570 1793 1597 1796
rect 1554 1733 1565 1736
rect 1538 1723 1545 1726
rect 1526 1703 1533 1706
rect 1530 1646 1533 1703
rect 1522 1643 1533 1646
rect 1542 1646 1545 1723
rect 1542 1643 1549 1646
rect 1506 1603 1517 1606
rect 1522 1546 1525 1643
rect 1506 1543 1525 1546
rect 1458 1356 1461 1386
rect 1450 1353 1461 1356
rect 1450 1333 1453 1353
rect 1458 1326 1461 1346
rect 1450 1323 1461 1326
rect 1450 1203 1453 1323
rect 1466 1283 1469 1393
rect 1490 1323 1493 1476
rect 1498 1413 1501 1466
rect 1506 1323 1509 1543
rect 1514 1503 1517 1536
rect 1522 1513 1525 1526
rect 1530 1473 1533 1616
rect 1538 1613 1541 1626
rect 1538 1533 1541 1546
rect 1546 1516 1549 1643
rect 1554 1563 1557 1676
rect 1570 1656 1573 1726
rect 1578 1673 1581 1793
rect 1562 1653 1573 1656
rect 1562 1573 1565 1653
rect 1570 1603 1581 1606
rect 1586 1596 1589 1736
rect 1594 1733 1597 1793
rect 1602 1783 1605 1826
rect 1610 1766 1613 1843
rect 1606 1763 1613 1766
rect 1594 1703 1597 1726
rect 1606 1666 1609 1763
rect 1618 1693 1621 2083
rect 1626 1933 1629 2193
rect 1634 2156 1637 2203
rect 1642 2163 1645 2216
rect 1650 2203 1653 2216
rect 1634 2153 1645 2156
rect 1626 1793 1629 1806
rect 1634 1716 1637 2126
rect 1642 2113 1645 2153
rect 1650 2133 1653 2176
rect 1658 2116 1661 2233
rect 1666 2213 1669 2246
rect 1674 2176 1677 2306
rect 1682 2186 1685 2343
rect 1738 2336 1741 2526
rect 1746 2513 1749 2546
rect 1754 2426 1757 2566
rect 1750 2423 1757 2426
rect 1750 2356 1753 2423
rect 1770 2416 1773 2556
rect 1954 2543 1997 2546
rect 1874 2533 1893 2536
rect 1914 2533 1925 2536
rect 1954 2533 1957 2543
rect 1978 2533 1989 2536
rect 1994 2533 1997 2543
rect 2042 2533 2061 2536
rect 2066 2533 2077 2536
rect 2082 2533 2085 2546
rect 2154 2543 2189 2546
rect 1794 2436 1797 2526
rect 1834 2523 1869 2526
rect 1810 2486 1813 2506
rect 1786 2433 1797 2436
rect 1806 2483 1813 2486
rect 1762 2413 1773 2416
rect 1750 2353 1757 2356
rect 1690 2316 1693 2336
rect 1714 2333 1741 2336
rect 1754 2333 1757 2353
rect 1690 2313 1697 2316
rect 1694 2196 1697 2313
rect 1706 2203 1709 2296
rect 1694 2193 1709 2196
rect 1682 2183 1693 2186
rect 1674 2173 1685 2176
rect 1654 2113 1661 2116
rect 1642 1966 1645 2076
rect 1654 2016 1657 2113
rect 1666 2016 1669 2136
rect 1674 2023 1677 2126
rect 1682 2073 1685 2173
rect 1690 2166 1693 2183
rect 1690 2163 1697 2166
rect 1694 2066 1697 2163
rect 1690 2063 1697 2066
rect 1654 2013 1661 2016
rect 1666 2013 1677 2016
rect 1658 1996 1661 2013
rect 1666 2003 1677 2006
rect 1658 1993 1677 1996
rect 1642 1963 1661 1966
rect 1658 1946 1661 1963
rect 1658 1943 1665 1946
rect 1650 1906 1653 1926
rect 1646 1903 1653 1906
rect 1646 1836 1649 1903
rect 1662 1896 1665 1943
rect 1674 1913 1677 1993
rect 1690 1956 1693 2063
rect 1698 2013 1701 2026
rect 1706 2003 1709 2193
rect 1714 2146 1717 2333
rect 1722 2213 1725 2286
rect 1730 2173 1733 2326
rect 1762 2316 1765 2413
rect 1770 2383 1773 2406
rect 1778 2343 1781 2416
rect 1786 2396 1789 2433
rect 1794 2413 1797 2426
rect 1806 2416 1809 2483
rect 1818 2423 1821 2516
rect 1826 2503 1829 2516
rect 1834 2496 1837 2523
rect 1826 2493 1837 2496
rect 1842 2513 1853 2516
rect 1806 2413 1813 2416
rect 1826 2413 1829 2493
rect 1842 2483 1845 2513
rect 1858 2506 1861 2516
rect 1850 2503 1861 2506
rect 1834 2443 1853 2446
rect 1834 2433 1837 2443
rect 1842 2423 1845 2436
rect 1850 2433 1853 2443
rect 1786 2393 1793 2396
rect 1754 2313 1765 2316
rect 1754 2246 1757 2313
rect 1754 2243 1765 2246
rect 1738 2206 1741 2226
rect 1738 2203 1749 2206
rect 1738 2183 1741 2196
rect 1746 2173 1749 2203
rect 1714 2143 1741 2146
rect 1714 2103 1717 2126
rect 1714 2003 1717 2016
rect 1690 1953 1697 1956
rect 1682 1933 1685 1946
rect 1694 1906 1697 1953
rect 1706 1923 1717 1926
rect 1722 1923 1725 2126
rect 1730 2003 1733 2136
rect 1738 2066 1741 2143
rect 1746 2083 1749 2146
rect 1738 2063 1745 2066
rect 1742 1996 1745 2063
rect 1738 1993 1745 1996
rect 1658 1893 1665 1896
rect 1690 1903 1697 1906
rect 1714 1906 1717 1923
rect 1730 1906 1733 1946
rect 1714 1903 1733 1906
rect 1646 1833 1653 1836
rect 1630 1713 1637 1716
rect 1602 1663 1609 1666
rect 1570 1593 1589 1596
rect 1570 1556 1573 1593
rect 1578 1583 1589 1586
rect 1578 1563 1581 1583
rect 1594 1576 1597 1626
rect 1602 1603 1605 1663
rect 1610 1596 1613 1656
rect 1618 1613 1621 1646
rect 1630 1636 1633 1713
rect 1630 1633 1637 1636
rect 1634 1613 1637 1633
rect 1586 1573 1597 1576
rect 1602 1593 1613 1596
rect 1554 1553 1573 1556
rect 1554 1533 1557 1553
rect 1562 1523 1581 1526
rect 1538 1493 1541 1516
rect 1546 1513 1565 1516
rect 1514 1323 1517 1416
rect 1522 1383 1525 1456
rect 1530 1423 1557 1426
rect 1530 1346 1533 1423
rect 1538 1403 1541 1416
rect 1554 1413 1557 1423
rect 1562 1406 1565 1513
rect 1578 1506 1581 1523
rect 1574 1503 1581 1506
rect 1574 1436 1577 1503
rect 1574 1433 1581 1436
rect 1546 1393 1549 1406
rect 1554 1403 1565 1406
rect 1570 1403 1573 1416
rect 1522 1343 1533 1346
rect 1522 1316 1525 1343
rect 1546 1336 1549 1346
rect 1506 1273 1509 1316
rect 1514 1313 1525 1316
rect 1530 1333 1549 1336
rect 1530 1316 1533 1333
rect 1530 1313 1537 1316
rect 1474 1203 1477 1266
rect 1514 1253 1517 1313
rect 1490 1203 1493 1226
rect 1514 1223 1517 1246
rect 1490 1133 1493 1146
rect 1498 1136 1501 1216
rect 1522 1203 1525 1296
rect 1534 1236 1537 1313
rect 1530 1233 1537 1236
rect 1530 1173 1533 1233
rect 1546 1216 1549 1326
rect 1538 1213 1549 1216
rect 1538 1186 1541 1213
rect 1554 1206 1557 1403
rect 1562 1333 1565 1386
rect 1578 1376 1581 1433
rect 1586 1393 1589 1573
rect 1594 1523 1597 1536
rect 1594 1443 1597 1516
rect 1602 1506 1605 1593
rect 1602 1503 1609 1506
rect 1606 1436 1609 1503
rect 1602 1433 1609 1436
rect 1602 1416 1605 1433
rect 1594 1413 1605 1416
rect 1570 1323 1573 1376
rect 1578 1373 1585 1376
rect 1582 1316 1585 1373
rect 1578 1313 1585 1316
rect 1562 1223 1565 1256
rect 1578 1226 1581 1313
rect 1578 1223 1589 1226
rect 1594 1223 1597 1413
rect 1602 1373 1605 1406
rect 1610 1393 1613 1416
rect 1610 1273 1613 1316
rect 1618 1293 1621 1606
rect 1626 1543 1629 1606
rect 1626 1466 1629 1536
rect 1634 1523 1637 1576
rect 1642 1473 1645 1816
rect 1626 1463 1637 1466
rect 1626 1413 1629 1426
rect 1626 1363 1629 1406
rect 1634 1403 1637 1463
rect 1650 1443 1653 1833
rect 1658 1823 1661 1893
rect 1690 1883 1693 1903
rect 1698 1856 1701 1876
rect 1666 1793 1669 1816
rect 1674 1783 1677 1806
rect 1658 1616 1661 1726
rect 1666 1723 1669 1736
rect 1674 1666 1677 1776
rect 1682 1716 1685 1856
rect 1698 1853 1705 1856
rect 1690 1723 1693 1836
rect 1702 1756 1705 1853
rect 1730 1826 1733 1896
rect 1738 1873 1741 1993
rect 1754 1936 1757 2216
rect 1762 2123 1765 2243
rect 1770 2213 1773 2226
rect 1778 2206 1781 2326
rect 1790 2286 1793 2393
rect 1802 2293 1805 2336
rect 1786 2283 1793 2286
rect 1786 2263 1789 2283
rect 1810 2266 1813 2413
rect 1858 2406 1861 2426
rect 1866 2413 1869 2523
rect 1874 2406 1877 2533
rect 1882 2453 1885 2516
rect 1858 2403 1877 2406
rect 1882 2393 1885 2426
rect 1890 2423 1893 2526
rect 1818 2273 1821 2336
rect 1826 2303 1829 2316
rect 1810 2263 1821 2266
rect 1770 2183 1773 2206
rect 1778 2203 1789 2206
rect 1786 2146 1789 2203
rect 1770 2056 1773 2146
rect 1786 2143 1797 2146
rect 1786 2103 1789 2126
rect 1766 2053 1773 2056
rect 1766 1966 1769 2053
rect 1766 1963 1773 1966
rect 1754 1933 1761 1936
rect 1746 1863 1749 1926
rect 1746 1826 1749 1836
rect 1722 1823 1733 1826
rect 1738 1823 1749 1826
rect 1714 1793 1717 1806
rect 1698 1753 1705 1756
rect 1682 1713 1693 1716
rect 1674 1663 1685 1666
rect 1658 1613 1677 1616
rect 1658 1593 1661 1606
rect 1682 1603 1685 1663
rect 1690 1613 1693 1706
rect 1698 1573 1701 1753
rect 1706 1713 1709 1736
rect 1722 1703 1725 1823
rect 1758 1816 1761 1933
rect 1730 1743 1733 1806
rect 1738 1733 1741 1816
rect 1758 1813 1765 1816
rect 1658 1493 1661 1556
rect 1706 1546 1709 1636
rect 1746 1616 1749 1766
rect 1762 1763 1765 1813
rect 1770 1803 1773 1963
rect 1778 1903 1781 2046
rect 1786 1953 1789 1996
rect 1794 1933 1797 2143
rect 1802 2133 1805 2206
rect 1810 2066 1813 2246
rect 1818 2186 1821 2263
rect 1826 2213 1829 2236
rect 1826 2193 1829 2206
rect 1834 2203 1837 2386
rect 1858 2333 1861 2346
rect 1842 2323 1853 2326
rect 1858 2313 1861 2326
rect 1898 2323 1901 2426
rect 1914 2403 1917 2533
rect 1922 2503 1925 2526
rect 1930 2413 1933 2496
rect 1922 2316 1925 2336
rect 1938 2333 1941 2346
rect 1946 2333 1949 2426
rect 1938 2323 1949 2326
rect 1922 2313 1949 2316
rect 1842 2223 1869 2226
rect 1818 2183 1837 2186
rect 1818 2103 1821 2136
rect 1802 2063 1813 2066
rect 1802 2013 1805 2063
rect 1810 2036 1813 2056
rect 1810 2033 1817 2036
rect 1786 1863 1789 1926
rect 1802 1866 1805 2006
rect 1814 1956 1817 2033
rect 1826 2016 1829 2136
rect 1834 2123 1837 2183
rect 1842 2123 1845 2136
rect 1850 2023 1853 2046
rect 1826 2013 1849 2016
rect 1826 1973 1829 2006
rect 1810 1953 1817 1956
rect 1810 1933 1813 1953
rect 1834 1936 1837 2006
rect 1846 1946 1849 2013
rect 1846 1943 1853 1946
rect 1826 1933 1837 1936
rect 1826 1886 1829 1933
rect 1850 1926 1853 1943
rect 1858 1933 1861 2216
rect 1866 2213 1869 2223
rect 1866 2196 1869 2206
rect 1882 2203 1885 2226
rect 1914 2213 1917 2226
rect 1922 2196 1925 2206
rect 1866 2193 1925 2196
rect 1930 2156 1933 2216
rect 1938 2203 1941 2276
rect 1946 2193 1949 2313
rect 1930 2153 1949 2156
rect 1914 2143 1933 2146
rect 1930 2136 1933 2143
rect 1866 2043 1877 2046
rect 1874 2013 1877 2043
rect 1882 2006 1885 2136
rect 1914 2123 1917 2136
rect 1930 2133 1941 2136
rect 1946 2133 1949 2153
rect 1898 2093 1901 2116
rect 1930 2063 1933 2126
rect 1938 2093 1941 2133
rect 1954 2076 1957 2526
rect 1978 2483 1981 2526
rect 1994 2513 1997 2526
rect 2058 2523 2061 2533
rect 2082 2516 2085 2526
rect 2010 2513 2085 2516
rect 1962 2433 1965 2446
rect 1962 2403 1965 2426
rect 1970 2413 1973 2436
rect 1994 2433 1997 2476
rect 2034 2436 2037 2506
rect 1962 2316 1965 2336
rect 1962 2313 1973 2316
rect 1970 2226 1973 2313
rect 1986 2273 1989 2426
rect 1994 2406 1997 2426
rect 1994 2403 2013 2406
rect 2002 2303 2005 2326
rect 2010 2323 2013 2403
rect 2018 2316 2021 2436
rect 2026 2433 2037 2436
rect 2026 2333 2029 2433
rect 2034 2416 2037 2426
rect 2050 2423 2069 2426
rect 2034 2413 2061 2416
rect 2058 2386 2061 2406
rect 2066 2393 2069 2423
rect 2074 2386 2077 2446
rect 2098 2413 2101 2536
rect 2154 2533 2157 2543
rect 2138 2496 2141 2526
rect 2114 2493 2141 2496
rect 2114 2476 2117 2493
rect 2110 2473 2117 2476
rect 2082 2393 2085 2406
rect 2058 2383 2077 2386
rect 2110 2386 2113 2473
rect 2162 2466 2165 2536
rect 2122 2463 2165 2466
rect 2110 2383 2117 2386
rect 2034 2333 2037 2376
rect 2010 2313 2021 2316
rect 2018 2273 2021 2313
rect 1962 2223 1973 2226
rect 1962 2133 1965 2223
rect 1986 2206 1989 2256
rect 2026 2243 2029 2316
rect 1978 2203 1989 2206
rect 1994 2203 1997 2226
rect 1970 2183 1973 2196
rect 1978 2146 1981 2203
rect 1986 2183 1989 2196
rect 1970 2143 1981 2146
rect 1946 2073 1957 2076
rect 1890 2013 1893 2056
rect 1866 2003 1885 2006
rect 1842 1886 1845 1926
rect 1850 1923 1861 1926
rect 1850 1903 1853 1916
rect 1826 1883 1837 1886
rect 1842 1883 1849 1886
rect 1802 1863 1829 1866
rect 1786 1853 1821 1856
rect 1786 1796 1789 1853
rect 1794 1843 1813 1846
rect 1794 1833 1797 1843
rect 1778 1793 1789 1796
rect 1794 1793 1797 1816
rect 1754 1743 1789 1746
rect 1778 1706 1781 1726
rect 1786 1713 1789 1743
rect 1802 1736 1805 1836
rect 1810 1823 1813 1843
rect 1818 1813 1821 1853
rect 1826 1806 1829 1863
rect 1818 1803 1829 1806
rect 1818 1746 1821 1803
rect 1818 1743 1825 1746
rect 1802 1733 1813 1736
rect 1794 1723 1805 1726
rect 1770 1703 1781 1706
rect 1770 1646 1773 1703
rect 1794 1663 1797 1723
rect 1810 1656 1813 1733
rect 1794 1653 1813 1656
rect 1770 1643 1789 1646
rect 1714 1583 1717 1616
rect 1674 1543 1709 1546
rect 1666 1463 1669 1536
rect 1674 1533 1677 1543
rect 1690 1533 1701 1536
rect 1714 1533 1717 1546
rect 1682 1506 1685 1526
rect 1678 1503 1685 1506
rect 1678 1416 1681 1503
rect 1690 1426 1693 1533
rect 1722 1526 1725 1616
rect 1746 1613 1757 1616
rect 1746 1606 1749 1613
rect 1738 1603 1749 1606
rect 1754 1603 1765 1606
rect 1770 1596 1773 1626
rect 1778 1613 1781 1636
rect 1762 1593 1773 1596
rect 1786 1593 1789 1643
rect 1794 1603 1797 1653
rect 1822 1646 1825 1743
rect 1818 1643 1825 1646
rect 1818 1616 1821 1643
rect 1834 1626 1837 1883
rect 1846 1746 1849 1883
rect 1846 1743 1853 1746
rect 1802 1613 1821 1616
rect 1826 1623 1837 1626
rect 1826 1613 1829 1623
rect 1698 1463 1701 1526
rect 1706 1523 1725 1526
rect 1706 1513 1709 1523
rect 1730 1503 1733 1536
rect 1738 1496 1741 1576
rect 1730 1493 1741 1496
rect 1690 1423 1697 1426
rect 1642 1413 1653 1416
rect 1650 1356 1653 1413
rect 1658 1366 1661 1416
rect 1678 1413 1685 1416
rect 1666 1373 1669 1406
rect 1674 1366 1677 1396
rect 1658 1363 1677 1366
rect 1650 1353 1661 1356
rect 1626 1323 1629 1346
rect 1650 1333 1653 1346
rect 1658 1333 1661 1353
rect 1682 1336 1685 1413
rect 1694 1376 1697 1423
rect 1714 1413 1717 1426
rect 1730 1406 1733 1493
rect 1746 1486 1749 1536
rect 1762 1523 1765 1593
rect 1770 1523 1773 1546
rect 1738 1483 1749 1486
rect 1738 1413 1741 1483
rect 1746 1413 1749 1426
rect 1714 1386 1717 1406
rect 1730 1403 1741 1406
rect 1690 1373 1697 1376
rect 1706 1383 1717 1386
rect 1690 1353 1693 1373
rect 1706 1343 1709 1383
rect 1722 1373 1725 1396
rect 1674 1333 1685 1336
rect 1714 1333 1717 1346
rect 1562 1213 1581 1216
rect 1554 1203 1565 1206
rect 1586 1196 1589 1223
rect 1582 1193 1589 1196
rect 1538 1183 1549 1186
rect 1498 1133 1509 1136
rect 1450 1106 1453 1126
rect 1474 1123 1501 1126
rect 1506 1106 1509 1133
rect 1426 1023 1437 1026
rect 1446 1103 1453 1106
rect 1498 1103 1509 1106
rect 1446 1026 1449 1103
rect 1446 1023 1453 1026
rect 1426 1013 1429 1023
rect 1330 983 1341 986
rect 1338 923 1341 983
rect 1434 943 1437 1016
rect 1450 1006 1453 1023
rect 1458 1013 1461 1096
rect 1498 1036 1501 1103
rect 1514 1056 1517 1136
rect 1522 1123 1525 1146
rect 1546 1116 1549 1183
rect 1582 1136 1585 1193
rect 1594 1143 1597 1216
rect 1658 1213 1661 1326
rect 1674 1316 1677 1333
rect 1670 1313 1677 1316
rect 1670 1256 1673 1313
rect 1666 1253 1673 1256
rect 1682 1253 1685 1326
rect 1706 1323 1725 1326
rect 1730 1323 1733 1336
rect 1666 1206 1669 1253
rect 1618 1146 1621 1206
rect 1658 1203 1669 1206
rect 1618 1143 1625 1146
rect 1538 1113 1549 1116
rect 1514 1053 1525 1056
rect 1522 1046 1525 1053
rect 1522 1043 1533 1046
rect 1490 1033 1501 1036
rect 1450 1003 1461 1006
rect 1290 883 1297 886
rect 1278 823 1285 826
rect 1282 806 1285 823
rect 1290 813 1293 883
rect 1306 813 1309 846
rect 1266 803 1277 806
rect 1282 803 1293 806
rect 1314 803 1317 836
rect 1354 826 1357 886
rect 1350 823 1357 826
rect 1242 793 1269 796
rect 1242 736 1245 756
rect 1238 733 1245 736
rect 1250 736 1253 776
rect 1250 733 1261 736
rect 1218 613 1221 686
rect 1238 646 1241 733
rect 1238 643 1245 646
rect 1234 613 1237 626
rect 1202 593 1237 596
rect 1170 543 1189 546
rect 1186 526 1189 543
rect 1126 513 1141 516
rect 1138 446 1141 513
rect 1178 473 1181 526
rect 1186 523 1197 526
rect 1194 513 1197 523
rect 1130 443 1141 446
rect 1066 366 1069 396
rect 1130 376 1133 443
rect 1154 433 1181 436
rect 1154 413 1157 433
rect 1154 383 1157 406
rect 1162 403 1165 416
rect 1130 373 1141 376
rect 1066 363 1085 366
rect 1082 346 1085 363
rect 1082 343 1089 346
rect 946 206 949 223
rect 994 213 997 283
rect 1034 223 1037 313
rect 1086 296 1089 343
rect 1082 293 1089 296
rect 1002 213 1061 216
rect 1058 206 1061 213
rect 938 203 949 206
rect 1018 196 1021 206
rect 978 193 1021 196
rect 858 113 861 126
rect 978 123 981 193
rect 1026 183 1029 206
rect 1058 203 1069 206
rect 1042 193 1061 196
rect 1066 123 1069 203
rect 1082 193 1085 293
rect 1098 203 1101 326
rect 1138 323 1141 373
rect 1154 293 1157 336
rect 1162 223 1165 326
rect 1170 313 1173 426
rect 1178 413 1181 433
rect 1202 383 1205 536
rect 1210 533 1213 546
rect 1218 523 1221 586
rect 1234 526 1237 593
rect 1242 573 1245 643
rect 1250 613 1253 726
rect 1250 546 1253 606
rect 1242 543 1253 546
rect 1234 523 1245 526
rect 1242 513 1245 523
rect 1250 423 1253 506
rect 1210 393 1213 406
rect 1226 336 1229 406
rect 1194 313 1197 336
rect 1226 333 1241 336
rect 1226 276 1229 326
rect 1238 286 1241 333
rect 1258 293 1261 536
rect 1266 516 1269 793
rect 1274 773 1277 803
rect 1274 733 1277 746
rect 1282 703 1285 726
rect 1290 696 1293 803
rect 1330 766 1333 806
rect 1338 793 1341 816
rect 1330 763 1341 766
rect 1314 733 1317 756
rect 1338 743 1341 763
rect 1350 746 1353 823
rect 1350 743 1357 746
rect 1306 716 1309 726
rect 1306 713 1341 716
rect 1282 693 1293 696
rect 1282 633 1285 693
rect 1290 613 1293 686
rect 1298 623 1309 626
rect 1290 603 1309 606
rect 1290 533 1293 603
rect 1314 543 1317 606
rect 1322 533 1325 646
rect 1338 626 1341 713
rect 1346 703 1349 726
rect 1338 623 1349 626
rect 1330 583 1333 616
rect 1346 566 1349 606
rect 1338 563 1349 566
rect 1266 513 1277 516
rect 1274 446 1277 513
rect 1266 443 1277 446
rect 1266 366 1269 443
rect 1274 376 1277 406
rect 1290 403 1293 426
rect 1314 376 1317 416
rect 1322 413 1325 516
rect 1338 506 1341 563
rect 1354 513 1357 743
rect 1362 703 1365 816
rect 1370 796 1373 846
rect 1378 803 1381 826
rect 1386 813 1389 876
rect 1402 813 1405 926
rect 1434 883 1437 936
rect 1458 923 1461 1003
rect 1482 986 1485 1006
rect 1478 983 1485 986
rect 1490 986 1493 1033
rect 1506 993 1509 1006
rect 1490 983 1501 986
rect 1370 793 1389 796
rect 1386 733 1389 793
rect 1394 773 1397 806
rect 1418 803 1421 826
rect 1418 726 1421 746
rect 1378 723 1389 726
rect 1410 723 1421 726
rect 1362 613 1365 636
rect 1362 573 1365 606
rect 1338 503 1349 506
rect 1346 456 1349 503
rect 1330 453 1349 456
rect 1274 373 1317 376
rect 1330 366 1333 453
rect 1266 363 1277 366
rect 1274 323 1277 363
rect 1282 363 1333 366
rect 1282 333 1285 363
rect 1238 283 1245 286
rect 1218 273 1229 276
rect 1218 226 1221 273
rect 1218 223 1229 226
rect 1098 113 1101 136
rect 1106 123 1109 216
rect 1114 193 1117 206
rect 1170 193 1173 206
rect 1154 133 1157 146
rect 1178 123 1181 206
rect 1226 203 1229 223
rect 1242 193 1245 283
rect 1290 226 1293 326
rect 1298 313 1301 326
rect 1314 313 1317 336
rect 1338 313 1341 416
rect 1370 386 1373 716
rect 1378 523 1381 676
rect 1386 603 1389 696
rect 1410 666 1413 723
rect 1426 673 1429 816
rect 1434 713 1437 726
rect 1410 663 1421 666
rect 1394 613 1397 626
rect 1410 623 1413 646
rect 1418 603 1421 663
rect 1426 603 1429 656
rect 1442 573 1445 856
rect 1466 813 1469 946
rect 1478 906 1481 983
rect 1498 966 1501 983
rect 1498 963 1505 966
rect 1478 903 1485 906
rect 1482 883 1485 903
rect 1502 886 1505 963
rect 1498 883 1505 886
rect 1498 866 1501 883
rect 1490 863 1501 866
rect 1450 773 1453 806
rect 1490 776 1493 863
rect 1514 833 1517 926
rect 1530 923 1533 1043
rect 1538 1013 1541 1113
rect 1570 993 1573 1136
rect 1582 1133 1589 1136
rect 1586 1026 1589 1133
rect 1610 1123 1613 1136
rect 1622 1096 1625 1143
rect 1618 1093 1625 1096
rect 1618 1076 1621 1093
rect 1582 1023 1589 1026
rect 1610 1073 1621 1076
rect 1582 976 1585 1023
rect 1594 976 1597 1016
rect 1610 993 1613 1073
rect 1634 1013 1637 1126
rect 1658 1056 1661 1203
rect 1698 1113 1701 1216
rect 1714 1056 1717 1206
rect 1738 1126 1741 1403
rect 1754 1373 1757 1446
rect 1762 1366 1765 1476
rect 1754 1363 1765 1366
rect 1746 1213 1749 1326
rect 1754 1316 1757 1363
rect 1770 1356 1773 1496
rect 1762 1353 1773 1356
rect 1762 1333 1765 1353
rect 1754 1313 1761 1316
rect 1758 1206 1761 1313
rect 1778 1256 1781 1536
rect 1786 1393 1789 1556
rect 1794 1413 1797 1546
rect 1802 1543 1805 1613
rect 1810 1523 1813 1606
rect 1818 1603 1829 1606
rect 1802 1406 1805 1506
rect 1826 1496 1829 1596
rect 1834 1563 1837 1616
rect 1842 1546 1845 1726
rect 1850 1653 1853 1743
rect 1858 1686 1861 1923
rect 1866 1706 1869 1956
rect 1898 1933 1901 2016
rect 1922 1996 1925 2016
rect 1914 1993 1925 1996
rect 1914 1946 1917 1993
rect 1914 1943 1925 1946
rect 1874 1903 1877 1916
rect 1874 1713 1877 1806
rect 1882 1793 1885 1816
rect 1890 1803 1893 1826
rect 1898 1816 1901 1866
rect 1906 1843 1909 1926
rect 1922 1923 1925 1943
rect 1922 1853 1925 1916
rect 1898 1813 1925 1816
rect 1906 1766 1909 1806
rect 1922 1793 1925 1813
rect 1930 1796 1933 2056
rect 1946 1966 1949 2073
rect 1962 2003 1965 2096
rect 1946 1963 1957 1966
rect 1938 1803 1941 1946
rect 1946 1913 1949 1936
rect 1954 1846 1957 1963
rect 1962 1923 1965 1996
rect 1970 1946 1973 2143
rect 1978 2123 1981 2136
rect 1986 2133 1989 2146
rect 1994 2053 1997 2136
rect 2018 2133 2021 2186
rect 2010 2123 2021 2126
rect 1986 2026 1989 2036
rect 1994 2033 2005 2036
rect 1978 2013 1981 2026
rect 1986 2023 2005 2026
rect 2010 2023 2013 2123
rect 2026 2083 2029 2216
rect 2042 2146 2045 2356
rect 2058 2323 2061 2383
rect 2114 2353 2117 2383
rect 2066 2333 2093 2336
rect 2034 2143 2045 2146
rect 2050 2133 2053 2146
rect 2058 2126 2061 2226
rect 2074 2213 2077 2266
rect 2066 2203 2077 2206
rect 2082 2193 2085 2206
rect 2090 2193 2093 2333
rect 2106 2293 2109 2316
rect 2122 2303 2125 2463
rect 2170 2403 2173 2526
rect 2186 2523 2189 2543
rect 2210 2533 2213 2556
rect 2138 2316 2141 2336
rect 2170 2333 2173 2346
rect 2066 2133 2069 2156
rect 2058 2123 2069 2126
rect 1970 1943 1981 1946
rect 1970 1906 1973 1936
rect 1946 1843 1957 1846
rect 1966 1903 1973 1906
rect 1946 1813 1949 1843
rect 1966 1826 1969 1903
rect 1954 1823 1969 1826
rect 1954 1813 1957 1823
rect 1962 1803 1965 1816
rect 1970 1796 1973 1806
rect 1930 1793 1973 1796
rect 1882 1733 1885 1746
rect 1898 1733 1901 1766
rect 1906 1763 1933 1766
rect 1922 1746 1925 1756
rect 1906 1743 1925 1746
rect 1890 1723 1901 1726
rect 1906 1723 1909 1743
rect 1866 1703 1909 1706
rect 1914 1703 1917 1736
rect 1858 1683 1869 1686
rect 1866 1626 1869 1683
rect 1858 1623 1869 1626
rect 1898 1623 1901 1636
rect 1850 1583 1853 1616
rect 1834 1543 1845 1546
rect 1850 1533 1853 1546
rect 1858 1543 1861 1623
rect 1890 1613 1901 1616
rect 1890 1606 1893 1613
rect 1866 1556 1869 1606
rect 1874 1603 1893 1606
rect 1866 1553 1885 1556
rect 1822 1493 1829 1496
rect 1794 1403 1805 1406
rect 1794 1343 1797 1403
rect 1810 1313 1813 1466
rect 1822 1426 1825 1493
rect 1822 1423 1829 1426
rect 1818 1343 1821 1406
rect 1826 1396 1829 1423
rect 1834 1413 1837 1486
rect 1850 1463 1853 1526
rect 1858 1506 1861 1536
rect 1874 1523 1877 1546
rect 1882 1533 1885 1553
rect 1898 1506 1901 1606
rect 1906 1593 1909 1703
rect 1922 1686 1925 1743
rect 1918 1683 1925 1686
rect 1918 1616 1921 1683
rect 1914 1613 1921 1616
rect 1914 1563 1917 1613
rect 1922 1536 1925 1606
rect 1906 1533 1925 1536
rect 1858 1503 1869 1506
rect 1842 1403 1845 1446
rect 1850 1413 1853 1456
rect 1866 1436 1869 1503
rect 1858 1433 1869 1436
rect 1890 1503 1901 1506
rect 1826 1393 1845 1396
rect 1818 1326 1821 1336
rect 1818 1323 1837 1326
rect 1778 1253 1785 1256
rect 1754 1203 1761 1206
rect 1754 1156 1757 1203
rect 1782 1186 1785 1253
rect 1842 1246 1845 1393
rect 1858 1343 1861 1433
rect 1866 1393 1869 1416
rect 1874 1373 1877 1396
rect 1850 1313 1853 1336
rect 1842 1243 1853 1246
rect 1778 1183 1785 1186
rect 1778 1163 1781 1183
rect 1754 1153 1781 1156
rect 1770 1133 1773 1146
rect 1650 1053 1661 1056
rect 1706 1053 1717 1056
rect 1730 1123 1741 1126
rect 1730 1056 1733 1123
rect 1730 1053 1741 1056
rect 1650 1006 1653 1053
rect 1674 1013 1693 1016
rect 1650 1003 1661 1006
rect 1658 983 1661 1003
rect 1674 976 1677 1013
rect 1706 993 1709 1053
rect 1738 1013 1741 1053
rect 1582 973 1589 976
rect 1594 973 1621 976
rect 1586 956 1589 973
rect 1586 953 1605 956
rect 1562 923 1565 936
rect 1570 876 1573 946
rect 1586 906 1589 926
rect 1586 903 1593 906
rect 1570 873 1581 876
rect 1522 833 1565 836
rect 1490 773 1501 776
rect 1450 713 1453 766
rect 1458 713 1461 726
rect 1458 563 1461 626
rect 1466 593 1469 736
rect 1482 733 1485 756
rect 1498 733 1501 773
rect 1506 733 1509 826
rect 1514 813 1525 816
rect 1530 763 1533 826
rect 1538 813 1549 816
rect 1562 813 1565 833
rect 1538 753 1541 806
rect 1546 783 1549 813
rect 1562 793 1565 806
rect 1578 803 1581 873
rect 1590 796 1593 903
rect 1602 826 1605 953
rect 1618 923 1621 973
rect 1642 973 1677 976
rect 1602 823 1613 826
rect 1586 793 1593 796
rect 1570 743 1581 746
rect 1546 733 1581 736
rect 1498 723 1509 726
rect 1554 723 1573 726
rect 1538 713 1549 716
rect 1410 536 1413 556
rect 1386 533 1413 536
rect 1410 523 1413 533
rect 1378 393 1381 416
rect 1394 403 1397 416
rect 1426 396 1429 536
rect 1466 443 1469 516
rect 1474 506 1477 706
rect 1482 523 1485 666
rect 1522 656 1525 676
rect 1518 653 1525 656
rect 1490 623 1493 636
rect 1518 606 1521 653
rect 1530 613 1533 626
rect 1538 623 1549 626
rect 1490 533 1493 606
rect 1498 593 1501 606
rect 1518 603 1525 606
rect 1474 503 1485 506
rect 1482 436 1485 503
rect 1474 433 1485 436
rect 1410 393 1429 396
rect 1370 383 1397 386
rect 1290 223 1325 226
rect 1258 163 1261 206
rect 1274 193 1277 206
rect 1314 203 1325 206
rect 1266 133 1269 146
rect 1234 113 1237 126
rect 1314 123 1317 203
rect 1330 193 1333 206
rect 1362 203 1365 326
rect 1394 323 1397 383
rect 1410 333 1413 393
rect 1434 336 1437 346
rect 1418 333 1437 336
rect 1442 333 1445 416
rect 1474 413 1477 433
rect 1450 333 1453 376
rect 1418 296 1421 333
rect 1490 326 1493 406
rect 1506 403 1509 536
rect 1514 533 1517 556
rect 1522 463 1525 603
rect 1538 543 1541 623
rect 1546 593 1549 606
rect 1554 603 1557 723
rect 1578 693 1581 716
rect 1546 523 1549 576
rect 1530 513 1541 516
rect 1562 493 1565 516
rect 1570 476 1573 536
rect 1578 533 1581 616
rect 1586 586 1589 793
rect 1594 606 1597 746
rect 1602 643 1605 816
rect 1610 633 1613 823
rect 1610 613 1613 626
rect 1594 603 1613 606
rect 1586 583 1593 586
rect 1590 506 1593 583
rect 1610 563 1613 596
rect 1618 556 1621 816
rect 1626 773 1629 966
rect 1642 813 1645 973
rect 1674 933 1677 946
rect 1658 893 1661 926
rect 1682 916 1685 976
rect 1690 966 1693 986
rect 1690 963 1697 966
rect 1674 913 1685 916
rect 1674 826 1677 913
rect 1694 906 1697 963
rect 1706 913 1709 926
rect 1690 903 1697 906
rect 1674 823 1681 826
rect 1634 733 1637 806
rect 1650 753 1653 816
rect 1642 736 1645 746
rect 1650 736 1653 746
rect 1642 733 1653 736
rect 1642 723 1645 733
rect 1650 706 1653 726
rect 1626 703 1653 706
rect 1658 703 1661 736
rect 1626 613 1629 703
rect 1650 676 1653 703
rect 1666 683 1669 806
rect 1678 746 1681 823
rect 1678 743 1685 746
rect 1674 676 1677 726
rect 1650 673 1677 676
rect 1682 666 1685 743
rect 1658 663 1685 666
rect 1626 593 1629 606
rect 1602 553 1621 556
rect 1602 523 1605 553
rect 1626 506 1629 536
rect 1590 503 1597 506
rect 1562 473 1573 476
rect 1562 426 1565 473
rect 1498 333 1501 356
rect 1426 313 1429 326
rect 1410 293 1421 296
rect 1410 203 1413 293
rect 1434 226 1437 326
rect 1482 306 1485 326
rect 1490 323 1501 326
rect 1506 323 1509 336
rect 1522 333 1525 426
rect 1498 313 1501 323
rect 1514 306 1517 326
rect 1482 303 1517 306
rect 1434 223 1477 226
rect 1418 166 1421 206
rect 1434 193 1437 206
rect 1346 123 1349 166
rect 1370 133 1373 146
rect 1410 123 1413 166
rect 1418 163 1453 166
rect 1474 163 1477 206
rect 1450 123 1453 163
rect 1474 133 1477 146
rect 1522 123 1525 166
rect 1538 123 1541 426
rect 1562 423 1573 426
rect 1570 403 1573 423
rect 1586 403 1589 426
rect 1594 383 1597 503
rect 1618 503 1629 506
rect 1618 436 1621 503
rect 1642 473 1645 636
rect 1650 503 1653 516
rect 1658 473 1661 663
rect 1674 613 1677 636
rect 1666 486 1669 526
rect 1674 523 1677 606
rect 1682 546 1685 596
rect 1690 583 1693 903
rect 1714 836 1717 946
rect 1722 923 1725 986
rect 1730 926 1733 996
rect 1730 923 1741 926
rect 1746 923 1749 1116
rect 1754 953 1757 1126
rect 1778 973 1781 1153
rect 1794 1123 1797 1216
rect 1810 1106 1813 1186
rect 1818 1173 1821 1206
rect 1850 1196 1853 1243
rect 1866 1213 1869 1336
rect 1890 1333 1893 1503
rect 1914 1456 1917 1526
rect 1914 1453 1925 1456
rect 1906 1413 1909 1426
rect 1914 1413 1917 1446
rect 1898 1393 1901 1406
rect 1890 1216 1893 1326
rect 1906 1303 1909 1406
rect 1914 1313 1917 1326
rect 1922 1226 1925 1453
rect 1930 1436 1933 1763
rect 1938 1723 1941 1793
rect 1978 1786 1981 1943
rect 1986 1926 1989 2016
rect 2018 1943 2021 2036
rect 2042 2026 2045 2116
rect 2066 2026 2069 2123
rect 2098 2116 2101 2136
rect 2090 2113 2101 2116
rect 2090 2046 2093 2113
rect 2090 2043 2101 2046
rect 2098 2026 2101 2043
rect 2042 2023 2061 2026
rect 2066 2023 2077 2026
rect 2026 2013 2045 2016
rect 2026 1996 2029 2013
rect 2066 2003 2069 2016
rect 2026 1993 2033 1996
rect 2030 1936 2033 1993
rect 1986 1923 1997 1926
rect 1986 1803 1989 1836
rect 1954 1783 1981 1786
rect 1954 1716 1957 1783
rect 1946 1713 1957 1716
rect 1938 1453 1941 1596
rect 1946 1576 1949 1713
rect 1970 1606 1973 1746
rect 1978 1723 1981 1736
rect 1954 1603 1973 1606
rect 1954 1593 1957 1603
rect 1946 1573 1953 1576
rect 1950 1446 1953 1573
rect 1962 1533 1965 1596
rect 1962 1496 1965 1526
rect 1970 1503 1973 1526
rect 1978 1523 1981 1656
rect 1986 1613 1989 1766
rect 1994 1753 1997 1816
rect 2002 1803 2005 1936
rect 2018 1916 2021 1936
rect 2014 1913 2021 1916
rect 2026 1933 2033 1936
rect 2014 1826 2017 1913
rect 2014 1823 2021 1826
rect 2010 1793 2013 1806
rect 1994 1623 1997 1646
rect 2002 1616 2005 1766
rect 2018 1733 2021 1823
rect 2026 1616 2029 1933
rect 2042 1926 2045 1946
rect 2050 1943 2053 1956
rect 2042 1923 2049 1926
rect 2034 1813 2037 1916
rect 2046 1806 2049 1923
rect 2042 1803 2049 1806
rect 2058 1803 2061 1996
rect 2074 1923 2077 2023
rect 2086 2023 2101 2026
rect 2086 1966 2089 2023
rect 2082 1963 2089 1966
rect 2082 1943 2085 1963
rect 2098 1946 2101 2006
rect 2106 1986 2109 2266
rect 2122 2213 2125 2226
rect 2130 2213 2133 2316
rect 2138 2313 2149 2316
rect 2146 2226 2149 2313
rect 2178 2293 2181 2416
rect 2186 2323 2189 2366
rect 2194 2333 2197 2346
rect 2202 2343 2205 2406
rect 2226 2336 2229 2416
rect 2202 2333 2229 2336
rect 2218 2293 2221 2326
rect 2142 2223 2149 2226
rect 2170 2223 2213 2226
rect 2114 1993 2117 2136
rect 2122 2013 2125 2196
rect 2130 2133 2133 2166
rect 2142 2156 2145 2223
rect 2170 2213 2173 2223
rect 2178 2213 2197 2216
rect 2154 2163 2157 2206
rect 2170 2193 2173 2206
rect 2178 2203 2181 2213
rect 2138 2153 2145 2156
rect 2130 2103 2133 2126
rect 2138 2096 2141 2153
rect 2146 2113 2149 2136
rect 2138 2093 2149 2096
rect 2130 1993 2133 2076
rect 2146 2026 2149 2093
rect 2138 2023 2149 2026
rect 2106 1983 2125 1986
rect 2094 1943 2101 1946
rect 2082 1893 2085 1936
rect 2042 1736 2045 1803
rect 2066 1756 2069 1816
rect 2082 1813 2085 1836
rect 2058 1753 2069 1756
rect 2042 1733 2053 1736
rect 2058 1723 2061 1753
rect 2034 1683 2037 1716
rect 1994 1613 2005 1616
rect 2018 1613 2029 1616
rect 1994 1536 1997 1613
rect 1986 1533 1997 1536
rect 2010 1526 2013 1536
rect 2002 1523 2013 1526
rect 2002 1516 2005 1523
rect 1978 1496 1981 1516
rect 1962 1493 1981 1496
rect 1986 1513 2005 1516
rect 1946 1443 1953 1446
rect 1930 1433 1937 1436
rect 1934 1366 1937 1433
rect 1930 1363 1937 1366
rect 1930 1313 1933 1363
rect 1938 1333 1941 1346
rect 1946 1303 1949 1443
rect 1970 1436 1973 1466
rect 1962 1433 1973 1436
rect 1962 1356 1965 1433
rect 1978 1413 1981 1426
rect 1986 1413 1989 1513
rect 2010 1503 2013 1516
rect 2018 1463 2021 1613
rect 2026 1583 2029 1606
rect 2034 1593 2037 1606
rect 2026 1523 2029 1566
rect 1978 1383 1981 1406
rect 1994 1393 1997 1416
rect 2010 1413 2013 1426
rect 1962 1353 1973 1356
rect 1962 1323 1965 1336
rect 1970 1333 1973 1353
rect 1922 1223 1949 1226
rect 1882 1213 1893 1216
rect 1834 1193 1853 1196
rect 1802 1103 1813 1106
rect 1802 1036 1805 1103
rect 1826 1056 1829 1126
rect 1834 1106 1837 1193
rect 1842 1133 1845 1156
rect 1850 1123 1853 1146
rect 1834 1103 1845 1106
rect 1822 1053 1829 1056
rect 1802 1033 1813 1036
rect 1786 956 1789 1016
rect 1762 953 1789 956
rect 1714 833 1725 836
rect 1706 773 1709 816
rect 1714 746 1717 816
rect 1722 803 1725 833
rect 1730 793 1733 816
rect 1738 803 1741 923
rect 1762 813 1765 953
rect 1802 943 1805 1006
rect 1810 963 1813 1033
rect 1786 856 1789 936
rect 1810 923 1813 936
rect 1822 916 1825 1053
rect 1842 1046 1845 1103
rect 1834 1043 1845 1046
rect 1822 913 1829 916
rect 1826 893 1829 913
rect 1834 886 1837 1043
rect 1866 1026 1869 1136
rect 1882 1133 1885 1213
rect 1874 1113 1877 1126
rect 1898 1096 1901 1216
rect 1890 1093 1901 1096
rect 1890 1036 1893 1093
rect 1890 1033 1901 1036
rect 1858 1023 1869 1026
rect 1850 963 1853 1016
rect 1858 1003 1861 1023
rect 1866 1013 1885 1016
rect 1898 1013 1901 1033
rect 1874 993 1877 1006
rect 1882 1003 1885 1013
rect 1858 896 1861 956
rect 1914 946 1917 1166
rect 1922 1133 1925 1146
rect 1930 1136 1933 1216
rect 1938 1153 1941 1206
rect 1946 1146 1949 1223
rect 1962 1206 1965 1316
rect 1978 1233 1981 1336
rect 1994 1303 1997 1346
rect 2002 1323 2005 1366
rect 2018 1333 2021 1406
rect 2034 1386 2037 1546
rect 2042 1493 2045 1626
rect 2058 1583 2061 1626
rect 2074 1613 2077 1806
rect 2082 1743 2085 1806
rect 2094 1746 2097 1943
rect 2106 1756 2109 1936
rect 2114 1923 2117 1946
rect 2122 1763 2125 1983
rect 2130 1926 2133 1946
rect 2138 1936 2141 2023
rect 2162 1946 2165 2176
rect 2170 2103 2173 2136
rect 2154 1943 2165 1946
rect 2138 1933 2149 1936
rect 2130 1923 2141 1926
rect 2138 1856 2141 1923
rect 2130 1853 2141 1856
rect 2106 1753 2125 1756
rect 2094 1743 2101 1746
rect 2082 1723 2085 1736
rect 2090 1703 2093 1726
rect 2090 1593 2093 1606
rect 2074 1533 2077 1556
rect 2066 1523 2077 1526
rect 2082 1523 2085 1536
rect 2058 1423 2061 1436
rect 2066 1416 2069 1523
rect 2074 1503 2077 1516
rect 2042 1413 2069 1416
rect 2034 1383 2045 1386
rect 2074 1383 2077 1416
rect 2090 1413 2093 1586
rect 2098 1453 2101 1743
rect 2106 1593 2109 1726
rect 2114 1613 2117 1746
rect 2122 1696 2125 1753
rect 2130 1743 2133 1853
rect 2138 1813 2141 1846
rect 2138 1713 2141 1806
rect 2146 1766 2149 1933
rect 2154 1916 2157 1943
rect 2178 1936 2181 1946
rect 2162 1933 2181 1936
rect 2154 1913 2161 1916
rect 2158 1836 2161 1913
rect 2170 1863 2173 1926
rect 2154 1833 2161 1836
rect 2154 1786 2157 1833
rect 2162 1803 2165 1816
rect 2178 1796 2181 1816
rect 2174 1793 2181 1796
rect 2154 1783 2165 1786
rect 2146 1763 2153 1766
rect 2150 1706 2153 1763
rect 2146 1703 2153 1706
rect 2122 1693 2133 1696
rect 2130 1606 2133 1693
rect 2146 1613 2149 1703
rect 2162 1626 2165 1783
rect 2174 1636 2177 1793
rect 2174 1633 2181 1636
rect 2158 1623 2165 1626
rect 2122 1603 2133 1606
rect 2106 1533 2109 1556
rect 2106 1433 2109 1526
rect 2114 1463 2117 1516
rect 2122 1503 2125 1603
rect 2158 1546 2161 1623
rect 2158 1543 2165 1546
rect 2146 1513 2149 1526
rect 2138 1413 2141 1486
rect 2154 1456 2157 1526
rect 2162 1513 2165 1543
rect 2150 1453 2157 1456
rect 2026 1306 2029 1326
rect 2022 1303 2029 1306
rect 2022 1236 2025 1303
rect 2042 1276 2045 1383
rect 2090 1343 2093 1406
rect 2106 1336 2109 1406
rect 2150 1396 2153 1453
rect 2034 1273 2045 1276
rect 2082 1333 2109 1336
rect 2130 1393 2153 1396
rect 2034 1256 2037 1273
rect 2034 1253 2053 1256
rect 2022 1233 2029 1236
rect 1970 1213 1973 1226
rect 2026 1213 2029 1233
rect 1954 1183 1957 1206
rect 1962 1203 1973 1206
rect 1962 1176 1965 1196
rect 1954 1173 1965 1176
rect 1954 1153 1957 1173
rect 1970 1156 1973 1203
rect 1986 1173 1989 1206
rect 2018 1173 2021 1196
rect 2050 1176 2053 1253
rect 2058 1216 2061 1226
rect 2058 1213 2069 1216
rect 2082 1193 2085 1333
rect 2106 1213 2109 1326
rect 2130 1266 2133 1393
rect 2170 1356 2173 1616
rect 2178 1593 2181 1633
rect 2178 1533 2181 1586
rect 2186 1526 2189 2206
rect 2210 1943 2213 2223
rect 2242 2203 2245 2556
rect 2258 2486 2261 2526
rect 2290 2523 2293 2546
rect 2306 2533 2309 2556
rect 2346 2486 2349 2526
rect 2258 2483 2285 2486
rect 2282 2413 2285 2483
rect 2338 2483 2349 2486
rect 2354 2486 2357 2556
rect 2386 2523 2389 2536
rect 2402 2533 2405 2556
rect 2570 2543 2597 2546
rect 2450 2523 2453 2536
rect 2482 2503 2485 2526
rect 2354 2483 2365 2486
rect 2338 2366 2341 2483
rect 2362 2403 2365 2483
rect 2274 2363 2317 2366
rect 2338 2363 2373 2366
rect 2410 2363 2413 2416
rect 2450 2413 2453 2466
rect 2274 2333 2277 2363
rect 2226 2123 2229 2166
rect 2218 2113 2245 2116
rect 2218 2023 2237 2026
rect 2218 2013 2221 2023
rect 2242 2013 2245 2113
rect 2258 2096 2261 2116
rect 2254 2093 2261 2096
rect 2226 1936 2229 1996
rect 2254 1946 2257 2093
rect 2266 2036 2269 2136
rect 2274 2133 2277 2306
rect 2290 2276 2293 2346
rect 2314 2323 2317 2363
rect 2290 2273 2309 2276
rect 2290 2193 2293 2216
rect 2306 2206 2309 2273
rect 2322 2213 2325 2306
rect 2354 2236 2357 2336
rect 2370 2323 2373 2363
rect 2458 2343 2461 2406
rect 2498 2393 2501 2536
rect 2514 2533 2525 2536
rect 2506 2523 2525 2526
rect 2522 2503 2525 2516
rect 2522 2363 2525 2406
rect 2530 2403 2533 2536
rect 2570 2533 2573 2543
rect 2578 2533 2589 2536
rect 2562 2523 2573 2526
rect 2578 2523 2589 2526
rect 2570 2516 2573 2523
rect 2570 2513 2581 2516
rect 2538 2423 2541 2436
rect 2578 2413 2581 2513
rect 2586 2503 2589 2523
rect 2594 2496 2597 2543
rect 2602 2503 2605 2536
rect 2610 2506 2613 2526
rect 2634 2506 2637 2526
rect 2610 2503 2637 2506
rect 2594 2493 2629 2496
rect 2626 2436 2629 2493
rect 2626 2433 2637 2436
rect 2394 2246 2397 2336
rect 2394 2243 2401 2246
rect 2346 2233 2357 2236
rect 2306 2203 2325 2206
rect 2322 2133 2325 2203
rect 2346 2176 2349 2233
rect 2370 2183 2373 2206
rect 2398 2196 2401 2243
rect 2410 2213 2413 2326
rect 2418 2313 2421 2326
rect 2458 2286 2461 2336
rect 2506 2323 2509 2336
rect 2538 2313 2541 2326
rect 2442 2283 2485 2286
rect 2394 2193 2401 2196
rect 2346 2173 2357 2176
rect 2354 2156 2357 2173
rect 2354 2153 2365 2156
rect 2282 2116 2285 2126
rect 2274 2113 2285 2116
rect 2266 2033 2277 2036
rect 2254 1943 2261 1946
rect 2226 1933 2233 1936
rect 2202 1923 2213 1926
rect 2194 1733 2197 1826
rect 2210 1813 2213 1896
rect 2218 1763 2221 1926
rect 2230 1866 2233 1933
rect 2226 1863 2233 1866
rect 2226 1813 2229 1863
rect 2242 1846 2245 1916
rect 2250 1913 2253 1926
rect 2234 1843 2245 1846
rect 2194 1623 2197 1656
rect 2202 1603 2205 1716
rect 2210 1696 2213 1726
rect 2218 1713 2221 1756
rect 2226 1733 2229 1746
rect 2234 1716 2237 1806
rect 2226 1713 2237 1716
rect 2242 1713 2245 1726
rect 2226 1696 2229 1713
rect 2250 1706 2253 1806
rect 2234 1703 2253 1706
rect 2210 1693 2217 1696
rect 2226 1693 2237 1696
rect 2214 1626 2217 1693
rect 2210 1623 2217 1626
rect 2210 1593 2213 1623
rect 2226 1613 2229 1626
rect 2218 1583 2221 1606
rect 2194 1533 2205 1536
rect 2234 1533 2237 1693
rect 2258 1633 2261 1943
rect 2266 1933 2269 2026
rect 2274 1833 2277 2033
rect 2282 1993 2285 2113
rect 2306 2086 2309 2126
rect 2346 2086 2349 2126
rect 2306 2083 2349 2086
rect 2362 2076 2365 2153
rect 2394 2113 2397 2193
rect 2354 2073 2365 2076
rect 2282 1923 2285 1936
rect 2290 1913 2301 1916
rect 2282 1833 2285 1846
rect 2266 1803 2269 1816
rect 2266 1703 2269 1746
rect 2274 1683 2277 1816
rect 2282 1803 2285 1826
rect 2290 1753 2293 1913
rect 2306 1836 2309 1926
rect 2322 1913 2325 1936
rect 2314 1893 2317 1906
rect 2330 1836 2333 1926
rect 2282 1703 2285 1726
rect 2290 1693 2293 1716
rect 2298 1686 2301 1836
rect 2306 1833 2333 1836
rect 2306 1813 2309 1826
rect 2306 1703 2309 1726
rect 2294 1683 2301 1686
rect 2258 1613 2269 1616
rect 2282 1613 2285 1636
rect 2294 1626 2297 1683
rect 2290 1623 2297 1626
rect 2258 1593 2261 1606
rect 2258 1533 2261 1546
rect 2178 1523 2189 1526
rect 2178 1403 2181 1523
rect 2194 1513 2205 1516
rect 2186 1396 2189 1506
rect 2210 1483 2213 1526
rect 2266 1523 2269 1613
rect 2290 1533 2293 1623
rect 2306 1613 2309 1626
rect 2298 1583 2301 1606
rect 2274 1446 2277 1466
rect 2274 1443 2281 1446
rect 2194 1413 2213 1416
rect 2218 1413 2237 1416
rect 2186 1393 2197 1396
rect 2202 1373 2205 1406
rect 2162 1353 2173 1356
rect 2162 1306 2165 1353
rect 2194 1333 2197 1356
rect 2210 1346 2213 1413
rect 2218 1393 2221 1406
rect 2226 1356 2229 1413
rect 2234 1393 2237 1406
rect 2250 1363 2253 1406
rect 2278 1396 2281 1443
rect 2290 1413 2293 1516
rect 2314 1446 2317 1766
rect 2322 1646 2325 1826
rect 2330 1723 2333 1833
rect 2338 1736 2341 1896
rect 2346 1823 2349 2006
rect 2354 1833 2357 2073
rect 2370 1943 2373 2006
rect 2362 1913 2373 1916
rect 2362 1843 2365 1913
rect 2370 1893 2373 1906
rect 2378 1856 2381 1926
rect 2394 1913 2397 1926
rect 2410 1856 2413 2016
rect 2418 2013 2421 2206
rect 2434 1993 2437 2146
rect 2442 1996 2445 2283
rect 2466 2236 2469 2276
rect 2462 2233 2469 2236
rect 2450 2203 2453 2216
rect 2462 2166 2465 2233
rect 2482 2203 2485 2283
rect 2546 2256 2549 2396
rect 2610 2343 2613 2396
rect 2578 2333 2589 2336
rect 2602 2333 2621 2336
rect 2546 2253 2553 2256
rect 2530 2196 2533 2216
rect 2550 2206 2553 2253
rect 2562 2213 2565 2276
rect 2570 2256 2573 2326
rect 2594 2313 2597 2326
rect 2570 2253 2589 2256
rect 2586 2216 2589 2253
rect 2594 2223 2605 2226
rect 2522 2193 2533 2196
rect 2546 2203 2553 2206
rect 2462 2163 2469 2166
rect 2466 2143 2469 2163
rect 2450 2133 2469 2136
rect 2450 2113 2453 2126
rect 2450 2003 2453 2016
rect 2474 2003 2477 2186
rect 2522 2146 2525 2193
rect 2498 2133 2501 2146
rect 2522 2143 2533 2146
rect 2498 2013 2501 2126
rect 2514 2006 2517 2126
rect 2530 2053 2533 2143
rect 2546 2136 2549 2203
rect 2570 2183 2573 2206
rect 2542 2133 2549 2136
rect 2542 2026 2545 2133
rect 2554 2096 2557 2126
rect 2554 2093 2565 2096
rect 2562 2046 2565 2093
rect 2578 2063 2581 2216
rect 2586 2213 2597 2216
rect 2594 2193 2597 2206
rect 2602 2203 2605 2216
rect 2594 2123 2597 2146
rect 2602 2133 2605 2146
rect 2610 2133 2613 2333
rect 2626 2326 2629 2416
rect 2634 2353 2637 2433
rect 2642 2343 2645 2526
rect 2658 2483 2661 2536
rect 2650 2413 2653 2426
rect 2666 2413 2669 2436
rect 2674 2383 2677 2536
rect 2682 2506 2685 2526
rect 2682 2503 2689 2506
rect 2698 2503 2701 2516
rect 2706 2513 2741 2516
rect 2626 2323 2669 2326
rect 2626 2296 2629 2316
rect 2666 2313 2669 2323
rect 2626 2293 2637 2296
rect 2634 2246 2637 2293
rect 2626 2243 2637 2246
rect 2626 2223 2629 2243
rect 2618 2133 2621 2146
rect 2618 2113 2621 2126
rect 2634 2123 2637 2216
rect 2650 2213 2653 2226
rect 2642 2166 2645 2206
rect 2658 2183 2661 2206
rect 2642 2163 2653 2166
rect 2642 2133 2645 2146
rect 2650 2136 2653 2163
rect 2666 2143 2669 2216
rect 2674 2193 2677 2356
rect 2686 2306 2689 2503
rect 2706 2413 2709 2513
rect 2738 2413 2741 2426
rect 2698 2343 2701 2406
rect 2754 2393 2757 2406
rect 2706 2333 2709 2356
rect 2706 2323 2717 2326
rect 2686 2303 2701 2306
rect 2698 2246 2701 2303
rect 2698 2243 2709 2246
rect 2706 2223 2709 2243
rect 2682 2203 2685 2216
rect 2690 2176 2693 2216
rect 2690 2173 2701 2176
rect 2650 2133 2661 2136
rect 2666 2133 2677 2136
rect 2554 2043 2565 2046
rect 2542 2023 2549 2026
rect 2498 2003 2517 2006
rect 2546 2006 2549 2023
rect 2554 2013 2557 2043
rect 2570 2013 2573 2026
rect 2578 2016 2581 2056
rect 2642 2026 2645 2126
rect 2586 2023 2613 2026
rect 2578 2013 2589 2016
rect 2594 2013 2605 2016
rect 2610 2013 2613 2023
rect 2546 2003 2565 2006
rect 2586 2003 2589 2013
rect 2626 2006 2629 2026
rect 2642 2023 2653 2026
rect 2658 2023 2661 2133
rect 2674 2096 2677 2133
rect 2698 2113 2701 2173
rect 2722 2156 2725 2386
rect 2738 2306 2741 2326
rect 2738 2303 2749 2306
rect 2746 2246 2749 2303
rect 2738 2243 2749 2246
rect 2738 2226 2741 2243
rect 2738 2223 2749 2226
rect 2714 2153 2725 2156
rect 2714 2096 2717 2153
rect 2730 2113 2733 2146
rect 2674 2093 2685 2096
rect 2714 2093 2733 2096
rect 2442 1993 2453 1996
rect 2450 1856 2453 1993
rect 2474 1946 2477 1996
rect 2474 1943 2485 1946
rect 2482 1866 2485 1943
rect 2498 1923 2501 2003
rect 2530 1893 2533 1926
rect 2538 1923 2541 1936
rect 2546 1923 2549 2003
rect 2602 1993 2605 2006
rect 2618 1956 2621 2006
rect 2626 2003 2645 2006
rect 2602 1953 2621 1956
rect 2602 1933 2605 1953
rect 2610 1943 2637 1946
rect 2610 1933 2613 1943
rect 2474 1863 2485 1866
rect 2378 1853 2389 1856
rect 2410 1853 2417 1856
rect 2362 1833 2381 1836
rect 2362 1823 2373 1826
rect 2354 1813 2365 1816
rect 2338 1733 2357 1736
rect 2338 1716 2341 1733
rect 2330 1713 2341 1716
rect 2346 1653 2349 1716
rect 2362 1703 2365 1813
rect 2378 1746 2381 1833
rect 2386 1753 2389 1853
rect 2394 1843 2405 1846
rect 2402 1826 2405 1843
rect 2398 1823 2405 1826
rect 2398 1776 2401 1823
rect 2414 1786 2417 1853
rect 2434 1853 2469 1856
rect 2434 1803 2437 1853
rect 2466 1806 2469 1853
rect 2474 1813 2477 1863
rect 2514 1813 2517 1826
rect 2530 1806 2533 1856
rect 2554 1853 2557 1916
rect 2562 1836 2565 1926
rect 2570 1903 2573 1916
rect 2586 1913 2589 1926
rect 2538 1813 2541 1826
rect 2546 1813 2549 1826
rect 2466 1803 2477 1806
rect 2530 1803 2541 1806
rect 2414 1783 2429 1786
rect 2398 1773 2405 1776
rect 2370 1743 2381 1746
rect 2370 1723 2373 1743
rect 2378 1733 2397 1736
rect 2394 1713 2397 1733
rect 2402 1723 2405 1773
rect 2410 1703 2413 1726
rect 2418 1703 2421 1716
rect 2426 1696 2429 1783
rect 2418 1693 2429 1696
rect 2322 1643 2365 1646
rect 2322 1576 2325 1616
rect 2330 1613 2333 1626
rect 2330 1593 2333 1606
rect 2322 1573 2341 1576
rect 2338 1486 2341 1573
rect 2322 1483 2341 1486
rect 2322 1463 2325 1483
rect 2314 1443 2321 1446
rect 2362 1443 2365 1643
rect 2378 1613 2381 1626
rect 2402 1603 2405 1626
rect 2274 1393 2281 1396
rect 2226 1353 2237 1356
rect 2210 1343 2229 1346
rect 2218 1323 2221 1336
rect 2226 1306 2229 1343
rect 2162 1303 2173 1306
rect 2122 1263 2133 1266
rect 2170 1286 2173 1303
rect 2222 1303 2229 1306
rect 2170 1283 2205 1286
rect 2122 1196 2125 1263
rect 2098 1193 2125 1196
rect 2050 1173 2061 1176
rect 1970 1153 1981 1156
rect 1946 1143 1973 1146
rect 1930 1133 1941 1136
rect 1930 1116 1933 1126
rect 1938 1123 1941 1133
rect 1954 1116 1957 1126
rect 1930 1113 1957 1116
rect 1962 1096 1965 1136
rect 1954 1093 1965 1096
rect 1954 1016 1957 1093
rect 1954 1013 1965 1016
rect 1962 993 1965 1013
rect 1970 1003 1973 1143
rect 1978 986 1981 1153
rect 2010 1136 2013 1166
rect 1986 1133 2013 1136
rect 2034 1133 2037 1146
rect 2042 1133 2045 1156
rect 1986 1106 1989 1133
rect 2058 1126 2061 1173
rect 1994 1123 2021 1126
rect 2050 1123 2061 1126
rect 2082 1123 2085 1186
rect 1986 1103 1997 1106
rect 1994 1026 1997 1103
rect 1986 1023 1997 1026
rect 1986 1003 1989 1023
rect 1962 983 1981 986
rect 1914 943 1933 946
rect 1866 913 1869 926
rect 1898 923 1901 936
rect 1930 896 1933 943
rect 1946 923 1949 946
rect 1858 893 1869 896
rect 1834 883 1845 886
rect 1778 853 1789 856
rect 1770 756 1773 776
rect 1766 753 1773 756
rect 1698 743 1717 746
rect 1698 556 1701 743
rect 1706 713 1709 736
rect 1714 733 1749 736
rect 1754 733 1757 746
rect 1714 723 1717 733
rect 1730 693 1733 716
rect 1738 713 1741 726
rect 1746 626 1749 733
rect 1766 666 1769 753
rect 1778 676 1781 853
rect 1826 756 1829 816
rect 1842 773 1845 883
rect 1866 836 1869 893
rect 1922 893 1933 896
rect 1858 833 1869 836
rect 1858 813 1861 833
rect 1890 816 1893 846
rect 1866 813 1893 816
rect 1906 833 1917 836
rect 1906 813 1909 833
rect 1922 826 1925 893
rect 1962 836 1965 983
rect 1970 926 1973 966
rect 2002 943 2005 966
rect 1978 933 1989 936
rect 2018 926 2021 1016
rect 2026 1013 2029 1026
rect 1970 923 1981 926
rect 2010 923 2021 926
rect 2010 856 2013 923
rect 2026 856 2029 936
rect 2042 933 2045 946
rect 2010 853 2021 856
rect 2026 853 2045 856
rect 1954 833 1965 836
rect 1922 823 1933 826
rect 1866 806 1869 813
rect 1850 803 1869 806
rect 1826 753 1841 756
rect 1794 733 1813 736
rect 1794 723 1797 733
rect 1802 676 1805 726
rect 1778 673 1785 676
rect 1766 663 1773 666
rect 1706 573 1709 626
rect 1730 623 1749 626
rect 1714 613 1741 616
rect 1730 563 1733 613
rect 1738 583 1741 606
rect 1698 553 1717 556
rect 1746 553 1749 623
rect 1754 603 1757 626
rect 1682 543 1709 546
rect 1682 533 1685 543
rect 1690 533 1701 536
rect 1706 533 1709 543
rect 1714 536 1717 553
rect 1714 533 1725 536
rect 1690 493 1693 526
rect 1706 486 1709 526
rect 1666 483 1709 486
rect 1706 463 1709 483
rect 1722 456 1725 533
rect 1754 523 1757 536
rect 1706 436 1709 456
rect 1618 433 1629 436
rect 1554 353 1565 356
rect 1562 323 1565 353
rect 1610 336 1613 416
rect 1626 403 1629 433
rect 1698 433 1709 436
rect 1714 453 1725 456
rect 1714 433 1717 453
rect 1642 403 1645 426
rect 1698 376 1701 433
rect 1722 423 1749 426
rect 1722 413 1725 423
rect 1698 373 1705 376
rect 1714 373 1717 406
rect 1602 333 1613 336
rect 1634 333 1637 346
rect 1602 306 1605 333
rect 1610 323 1621 326
rect 1682 323 1685 336
rect 1602 303 1621 306
rect 1618 223 1621 303
rect 1702 276 1705 373
rect 1722 336 1725 346
rect 1690 273 1705 276
rect 1714 333 1725 336
rect 1602 213 1613 216
rect 1562 143 1565 206
rect 1594 193 1597 206
rect 1594 133 1597 146
rect 1578 86 1581 126
rect 1602 86 1605 136
rect 1610 123 1613 213
rect 1618 163 1621 206
rect 1690 176 1693 273
rect 1714 203 1717 333
rect 1730 326 1733 416
rect 1738 333 1741 346
rect 1722 316 1725 326
rect 1730 323 1741 326
rect 1746 316 1749 336
rect 1754 333 1757 406
rect 1762 373 1765 646
rect 1770 573 1773 663
rect 1782 606 1785 673
rect 1794 673 1805 676
rect 1794 613 1797 673
rect 1818 626 1821 726
rect 1826 703 1829 716
rect 1838 646 1841 753
rect 1838 643 1845 646
rect 1818 623 1829 626
rect 1826 606 1829 623
rect 1834 613 1837 626
rect 1842 613 1845 643
rect 1782 603 1797 606
rect 1778 533 1781 546
rect 1786 533 1789 596
rect 1770 513 1773 526
rect 1770 396 1773 416
rect 1778 403 1781 476
rect 1794 396 1797 603
rect 1810 583 1813 606
rect 1802 496 1805 576
rect 1818 543 1821 606
rect 1826 603 1837 606
rect 1842 533 1845 546
rect 1850 533 1853 803
rect 1882 756 1885 806
rect 1882 753 1901 756
rect 1858 723 1861 736
rect 1866 733 1885 736
rect 1866 703 1869 733
rect 1890 726 1893 746
rect 1874 723 1893 726
rect 1858 533 1861 596
rect 1866 526 1869 616
rect 1818 513 1821 526
rect 1802 493 1813 496
rect 1770 393 1797 396
rect 1722 313 1749 316
rect 1690 173 1733 176
rect 1650 133 1653 156
rect 1674 123 1677 146
rect 1730 123 1733 173
rect 1746 133 1749 156
rect 1778 153 1781 393
rect 1810 376 1813 493
rect 1834 443 1837 526
rect 1842 523 1853 526
rect 1858 523 1869 526
rect 1874 523 1877 723
rect 1882 703 1885 716
rect 1898 696 1901 753
rect 1906 713 1909 726
rect 1914 723 1917 786
rect 1922 696 1925 816
rect 1890 693 1901 696
rect 1914 693 1925 696
rect 1890 626 1893 693
rect 1882 623 1893 626
rect 1914 626 1917 693
rect 1914 623 1925 626
rect 1882 586 1885 623
rect 1890 593 1893 606
rect 1882 583 1893 586
rect 1842 506 1845 523
rect 1842 503 1849 506
rect 1846 436 1849 503
rect 1842 433 1849 436
rect 1842 413 1845 433
rect 1858 403 1861 523
rect 1842 393 1853 396
rect 1802 373 1813 376
rect 1802 353 1805 373
rect 1802 323 1805 346
rect 1794 163 1813 166
rect 1794 123 1797 163
rect 1810 136 1813 163
rect 1818 153 1821 206
rect 1810 133 1837 136
rect 1842 123 1845 386
rect 1850 306 1853 393
rect 1866 383 1869 406
rect 1858 323 1861 376
rect 1874 323 1877 466
rect 1882 413 1885 526
rect 1890 523 1893 583
rect 1898 533 1901 606
rect 1914 586 1917 606
rect 1922 596 1925 623
rect 1930 603 1933 823
rect 1938 743 1941 826
rect 1954 786 1957 833
rect 1954 783 1965 786
rect 1938 693 1941 736
rect 1954 703 1957 736
rect 1962 723 1965 783
rect 1978 746 1981 806
rect 2002 793 2005 816
rect 2010 746 2013 776
rect 1978 743 2013 746
rect 1994 733 2005 736
rect 1954 643 1973 646
rect 1922 593 1941 596
rect 1906 583 1917 586
rect 1914 533 1917 546
rect 1906 493 1909 526
rect 1922 523 1925 566
rect 1898 396 1901 436
rect 1890 393 1901 396
rect 1890 326 1893 393
rect 1906 346 1909 406
rect 1930 346 1933 536
rect 1938 513 1941 593
rect 1954 586 1957 643
rect 1962 613 1965 636
rect 1970 623 1973 643
rect 1970 593 1973 606
rect 1954 583 1973 586
rect 1962 426 1965 526
rect 1970 516 1973 583
rect 1978 533 1981 726
rect 2010 716 2013 743
rect 2002 713 2013 716
rect 1986 613 1989 656
rect 2002 596 2005 713
rect 2018 603 2021 853
rect 2042 776 2045 853
rect 2050 813 2053 1123
rect 2098 1026 2101 1193
rect 2106 1133 2109 1176
rect 2130 1166 2133 1236
rect 2170 1226 2173 1283
rect 2170 1223 2177 1226
rect 2154 1213 2165 1216
rect 2130 1163 2137 1166
rect 2114 1133 2117 1146
rect 2066 1003 2069 1026
rect 2074 1023 2101 1026
rect 2074 1003 2077 1023
rect 2058 943 2061 966
rect 2082 906 2085 926
rect 2074 903 2085 906
rect 2074 836 2077 903
rect 2074 833 2085 836
rect 2082 813 2085 833
rect 2026 773 2045 776
rect 2026 716 2029 773
rect 2050 733 2053 746
rect 2058 723 2061 806
rect 2066 716 2069 736
rect 2074 723 2077 736
rect 2026 713 2037 716
rect 2034 646 2037 713
rect 2026 643 2037 646
rect 2058 713 2069 716
rect 2002 593 2013 596
rect 2010 576 2013 593
rect 2010 573 2017 576
rect 1986 543 2005 546
rect 1986 523 1989 543
rect 1994 523 1997 536
rect 2002 533 2005 543
rect 2014 526 2017 573
rect 2010 523 2017 526
rect 1970 513 1989 516
rect 1962 423 1969 426
rect 1938 413 1949 416
rect 1906 343 1933 346
rect 1906 333 1909 343
rect 1890 323 1901 326
rect 1850 303 1861 306
rect 1858 236 1861 303
rect 1850 233 1861 236
rect 1850 143 1853 233
rect 1866 176 1869 216
rect 1898 213 1901 323
rect 1914 313 1917 326
rect 1922 323 1925 336
rect 1930 333 1933 343
rect 1882 203 1909 206
rect 1882 176 1885 203
rect 1930 186 1933 326
rect 1938 323 1941 356
rect 1946 346 1949 406
rect 1954 383 1957 416
rect 1966 366 1969 423
rect 1978 413 1981 436
rect 1986 406 1989 513
rect 2010 436 2013 523
rect 2026 443 2029 643
rect 2034 613 2037 626
rect 2050 536 2053 616
rect 2058 593 2061 713
rect 2082 703 2085 726
rect 2090 646 2093 896
rect 2106 836 2109 1016
rect 2122 1003 2125 1156
rect 2134 1116 2137 1163
rect 2154 1146 2157 1213
rect 2146 1143 2157 1146
rect 2146 1123 2149 1143
rect 2162 1123 2165 1176
rect 2174 1116 2177 1223
rect 2186 1133 2189 1216
rect 2202 1213 2205 1283
rect 2222 1236 2225 1303
rect 2222 1233 2229 1236
rect 2226 1213 2229 1233
rect 2194 1203 2205 1206
rect 2210 1173 2213 1206
rect 2202 1133 2205 1156
rect 2134 1113 2149 1116
rect 2146 1066 2149 1113
rect 2170 1113 2177 1116
rect 2146 1063 2157 1066
rect 2146 1013 2149 1026
rect 2154 1006 2157 1063
rect 2170 1056 2173 1113
rect 2146 1003 2157 1006
rect 2166 1053 2173 1056
rect 2130 853 2133 936
rect 2138 913 2141 926
rect 2146 896 2149 1003
rect 2166 976 2169 1053
rect 2202 1013 2205 1126
rect 2210 1003 2213 1016
rect 2166 973 2173 976
rect 2170 933 2173 973
rect 2234 943 2237 1353
rect 2274 1273 2277 1393
rect 2242 1213 2245 1236
rect 2282 1213 2293 1216
rect 2298 1206 2301 1416
rect 2318 1376 2321 1443
rect 2418 1426 2421 1693
rect 2474 1686 2477 1803
rect 2538 1766 2541 1803
rect 2554 1796 2557 1836
rect 2562 1833 2573 1836
rect 2562 1823 2565 1833
rect 2570 1803 2573 1826
rect 2578 1796 2581 1846
rect 2554 1793 2581 1796
rect 2586 1823 2597 1826
rect 2538 1763 2545 1766
rect 2498 1706 2501 1726
rect 2498 1703 2509 1706
rect 2474 1683 2485 1686
rect 2482 1666 2485 1683
rect 2482 1663 2489 1666
rect 2442 1613 2445 1626
rect 2486 1576 2489 1663
rect 2506 1646 2509 1703
rect 2542 1686 2545 1763
rect 2586 1736 2589 1823
rect 2554 1723 2557 1736
rect 2578 1733 2589 1736
rect 2498 1643 2509 1646
rect 2538 1683 2545 1686
rect 2498 1613 2501 1643
rect 2514 1603 2517 1616
rect 2522 1603 2525 1616
rect 2482 1573 2489 1576
rect 2482 1483 2485 1573
rect 2530 1523 2533 1606
rect 2538 1583 2541 1683
rect 2546 1603 2549 1626
rect 2546 1536 2549 1596
rect 2554 1546 2557 1616
rect 2562 1613 2565 1726
rect 2602 1716 2605 1926
rect 2626 1916 2629 1936
rect 2634 1923 2637 1943
rect 2642 1933 2645 2003
rect 2650 1983 2653 2023
rect 2666 2016 2669 2066
rect 2682 2036 2685 2093
rect 2658 2013 2669 2016
rect 2674 2033 2685 2036
rect 2674 2016 2677 2033
rect 2674 2013 2717 2016
rect 2658 1953 2661 2013
rect 2674 2006 2677 2013
rect 2666 2003 2677 2006
rect 2682 1983 2685 1996
rect 2650 1943 2677 1946
rect 2658 1933 2669 1936
rect 2666 1916 2669 1926
rect 2626 1913 2669 1916
rect 2626 1833 2637 1836
rect 2618 1813 2621 1826
rect 2626 1806 2629 1833
rect 2642 1823 2645 1846
rect 2658 1823 2661 1856
rect 2634 1813 2669 1816
rect 2618 1803 2629 1806
rect 2674 1803 2677 1943
rect 2714 1933 2717 1996
rect 2722 1933 2725 1946
rect 2730 1933 2733 2093
rect 2738 1993 2741 2006
rect 2690 1903 2693 1926
rect 2706 1913 2709 1926
rect 2682 1803 2701 1806
rect 2706 1803 2709 1816
rect 2610 1733 2613 1746
rect 2618 1733 2621 1803
rect 2650 1743 2669 1746
rect 2650 1733 2653 1743
rect 2682 1733 2685 1803
rect 2722 1756 2725 1926
rect 2730 1903 2733 1926
rect 2746 1846 2749 2016
rect 2730 1843 2749 1846
rect 2730 1813 2733 1843
rect 2722 1753 2733 1756
rect 2706 1743 2725 1746
rect 2602 1713 2629 1716
rect 2666 1713 2669 1726
rect 2690 1723 2693 1736
rect 2706 1733 2709 1743
rect 2730 1733 2733 1753
rect 2738 1713 2741 1726
rect 2602 1613 2613 1616
rect 2554 1543 2573 1546
rect 2546 1533 2565 1536
rect 2594 1533 2597 1606
rect 2618 1573 2621 1626
rect 2626 1613 2629 1713
rect 2642 1623 2669 1626
rect 2642 1613 2645 1623
rect 2650 1613 2669 1616
rect 2626 1583 2629 1606
rect 2642 1546 2645 1606
rect 2634 1543 2645 1546
rect 2634 1533 2637 1543
rect 2562 1523 2565 1533
rect 2414 1423 2421 1426
rect 2314 1373 2321 1376
rect 2314 1276 2317 1373
rect 2330 1346 2333 1416
rect 2346 1363 2349 1406
rect 2370 1376 2373 1416
rect 2354 1373 2373 1376
rect 2414 1356 2417 1423
rect 2414 1353 2421 1356
rect 2330 1343 2349 1346
rect 2330 1333 2341 1336
rect 2330 1283 2333 1326
rect 2338 1313 2341 1326
rect 2314 1273 2333 1276
rect 2314 1213 2325 1216
rect 2266 1193 2269 1206
rect 2290 1203 2301 1206
rect 2250 1086 2253 1126
rect 2282 1123 2285 1186
rect 2298 1146 2301 1203
rect 2306 1163 2309 1206
rect 2330 1196 2333 1273
rect 2346 1213 2349 1343
rect 2362 1206 2365 1346
rect 2386 1253 2389 1326
rect 2402 1323 2405 1336
rect 2410 1296 2413 1336
rect 2418 1326 2421 1353
rect 2426 1333 2429 1416
rect 2442 1363 2445 1406
rect 2466 1393 2469 1416
rect 2418 1323 2429 1326
rect 2402 1293 2413 1296
rect 2402 1236 2405 1293
rect 2386 1213 2389 1236
rect 2402 1233 2413 1236
rect 2322 1193 2333 1196
rect 2298 1143 2309 1146
rect 2250 1083 2293 1086
rect 2250 963 2253 996
rect 2202 933 2253 936
rect 2142 893 2149 896
rect 2106 833 2125 836
rect 2106 813 2117 816
rect 2106 733 2109 813
rect 2114 793 2117 806
rect 2122 783 2125 833
rect 2130 803 2133 826
rect 2142 776 2145 893
rect 2142 773 2149 776
rect 2130 733 2133 746
rect 2138 733 2141 756
rect 2114 723 2133 726
rect 2090 643 2101 646
rect 2130 643 2133 716
rect 2042 533 2053 536
rect 2042 446 2045 533
rect 2042 443 2053 446
rect 2010 433 2029 436
rect 1986 403 1997 406
rect 1962 363 1969 366
rect 1962 346 1965 363
rect 2026 356 2029 433
rect 2026 353 2037 356
rect 1946 343 1989 346
rect 1946 323 1949 343
rect 1978 323 1981 336
rect 1986 333 1989 343
rect 1986 323 1997 326
rect 1986 306 1989 323
rect 1978 303 1989 306
rect 1978 246 1981 303
rect 1978 243 1989 246
rect 1986 206 1989 243
rect 1938 193 1941 206
rect 1962 203 1989 206
rect 1866 173 1885 176
rect 1898 183 1933 186
rect 1898 133 1901 183
rect 1930 173 1933 183
rect 1954 123 1957 136
rect 2002 123 2005 326
rect 2010 313 2013 336
rect 2018 333 2029 336
rect 2034 326 2037 353
rect 2026 323 2037 326
rect 2026 123 2029 323
rect 2050 313 2053 443
rect 2058 413 2061 526
rect 2066 523 2069 626
rect 2074 603 2077 636
rect 2082 513 2085 616
rect 2098 576 2101 643
rect 2146 636 2149 773
rect 2154 733 2157 926
rect 2202 923 2205 933
rect 2186 913 2213 916
rect 2162 793 2165 806
rect 2162 636 2165 786
rect 2170 733 2173 856
rect 2186 803 2189 913
rect 2218 896 2221 926
rect 2210 893 2221 896
rect 2210 826 2213 893
rect 2226 836 2229 906
rect 2250 886 2253 933
rect 2266 903 2269 916
rect 2274 893 2277 936
rect 2282 923 2285 1016
rect 2290 1003 2293 1083
rect 2306 1056 2309 1143
rect 2322 1106 2325 1193
rect 2338 1113 2341 1206
rect 2346 1203 2365 1206
rect 2346 1143 2349 1203
rect 2402 1193 2405 1216
rect 2362 1133 2365 1156
rect 2322 1103 2333 1106
rect 2298 1053 2309 1056
rect 2298 1033 2301 1053
rect 2330 1026 2333 1103
rect 2322 1023 2333 1026
rect 2290 963 2293 996
rect 2290 933 2301 936
rect 2306 933 2309 946
rect 2250 883 2261 886
rect 2226 833 2253 836
rect 2202 823 2213 826
rect 2226 823 2245 826
rect 2178 733 2181 756
rect 2194 746 2197 816
rect 2202 793 2205 823
rect 2210 783 2213 806
rect 2194 743 2237 746
rect 2170 643 2173 716
rect 2178 693 2181 726
rect 2146 633 2157 636
rect 2162 633 2173 636
rect 2090 573 2101 576
rect 2090 393 2093 573
rect 2098 533 2101 556
rect 2106 533 2117 536
rect 2106 426 2109 526
rect 2122 523 2125 616
rect 2130 523 2133 626
rect 2138 613 2149 616
rect 2138 593 2141 606
rect 2154 573 2157 633
rect 2162 603 2165 616
rect 2170 593 2173 633
rect 2186 623 2189 736
rect 2194 686 2197 743
rect 2210 733 2229 736
rect 2234 733 2237 743
rect 2250 736 2253 833
rect 2242 733 2253 736
rect 2226 723 2229 733
rect 2258 716 2261 883
rect 2266 823 2293 826
rect 2194 683 2205 686
rect 2202 613 2205 683
rect 2226 636 2229 716
rect 2250 713 2261 716
rect 2250 646 2253 713
rect 2266 683 2269 746
rect 2210 633 2229 636
rect 2234 643 2253 646
rect 2226 606 2229 626
rect 2170 533 2173 546
rect 2098 423 2109 426
rect 2066 213 2069 326
rect 2098 313 2101 423
rect 2114 403 2117 416
rect 2122 413 2125 446
rect 2114 333 2117 346
rect 2154 323 2157 416
rect 2162 413 2165 436
rect 2178 433 2181 526
rect 2186 513 2189 536
rect 2194 523 2197 606
rect 2218 603 2229 606
rect 2202 523 2205 546
rect 2218 516 2221 603
rect 2234 523 2237 643
rect 2250 623 2253 636
rect 2242 533 2245 606
rect 2258 543 2261 556
rect 2218 513 2237 516
rect 2210 393 2213 406
rect 2194 323 2197 386
rect 2218 346 2221 436
rect 2234 403 2237 513
rect 2266 386 2269 626
rect 2274 553 2277 816
rect 2282 796 2285 816
rect 2290 813 2293 823
rect 2282 793 2289 796
rect 2286 666 2289 793
rect 2282 663 2289 666
rect 2282 613 2285 663
rect 2290 613 2293 646
rect 2282 586 2285 606
rect 2282 583 2293 586
rect 2290 506 2293 583
rect 2298 576 2301 926
rect 2306 903 2309 926
rect 2314 923 2317 956
rect 2322 916 2325 1023
rect 2314 913 2325 916
rect 2306 803 2309 816
rect 2314 803 2317 913
rect 2330 896 2333 1016
rect 2354 956 2357 1036
rect 2370 963 2373 996
rect 2326 893 2333 896
rect 2338 953 2357 956
rect 2326 806 2329 893
rect 2322 803 2329 806
rect 2306 733 2309 746
rect 2306 673 2309 726
rect 2306 623 2309 636
rect 2314 613 2317 626
rect 2322 613 2325 803
rect 2338 786 2341 953
rect 2334 783 2341 786
rect 2334 676 2337 783
rect 2346 716 2349 816
rect 2354 726 2357 936
rect 2362 813 2365 826
rect 2378 806 2381 1016
rect 2386 1013 2389 1126
rect 2410 1113 2413 1233
rect 2418 1213 2421 1286
rect 2426 1263 2429 1323
rect 2442 1236 2445 1326
rect 2474 1316 2477 1336
rect 2482 1323 2485 1456
rect 2522 1346 2525 1416
rect 2538 1366 2541 1406
rect 2538 1363 2565 1366
rect 2490 1333 2493 1346
rect 2522 1343 2549 1346
rect 2514 1323 2525 1326
rect 2530 1316 2533 1326
rect 2474 1313 2533 1316
rect 2538 1313 2541 1336
rect 2546 1323 2549 1343
rect 2562 1316 2565 1363
rect 2554 1313 2565 1316
rect 2554 1263 2557 1313
rect 2434 1233 2445 1236
rect 2434 1186 2437 1233
rect 2434 1183 2445 1186
rect 2442 1146 2445 1183
rect 2458 1153 2461 1206
rect 2442 1143 2453 1146
rect 2442 1123 2445 1136
rect 2450 1076 2453 1143
rect 2434 1073 2453 1076
rect 2434 966 2437 1073
rect 2434 963 2453 966
rect 2386 923 2389 936
rect 2434 923 2437 946
rect 2442 883 2445 936
rect 2450 843 2453 963
rect 2458 856 2461 1116
rect 2466 1106 2469 1146
rect 2490 1126 2493 1146
rect 2498 1133 2501 1216
rect 2538 1213 2541 1236
rect 2506 1126 2509 1146
rect 2490 1123 2509 1126
rect 2538 1106 2541 1126
rect 2466 1103 2485 1106
rect 2482 1016 2485 1103
rect 2530 1103 2541 1106
rect 2530 1046 2533 1103
rect 2530 1043 2541 1046
rect 2466 1013 2485 1016
rect 2514 1023 2533 1026
rect 2514 1013 2517 1023
rect 2466 993 2469 1013
rect 2522 1006 2525 1016
rect 2530 1013 2533 1023
rect 2538 1006 2541 1043
rect 2554 1016 2557 1206
rect 2578 1126 2581 1446
rect 2586 1376 2589 1416
rect 2626 1413 2629 1526
rect 2642 1513 2645 1536
rect 2650 1523 2653 1546
rect 2666 1523 2669 1613
rect 2682 1603 2685 1636
rect 2714 1623 2717 1636
rect 2690 1593 2693 1606
rect 2674 1513 2677 1536
rect 2698 1523 2701 1616
rect 2714 1546 2717 1606
rect 2722 1603 2725 1616
rect 2706 1543 2717 1546
rect 2602 1403 2629 1406
rect 2602 1376 2605 1403
rect 2634 1396 2637 1446
rect 2626 1393 2637 1396
rect 2642 1393 2645 1416
rect 2658 1376 2661 1486
rect 2706 1413 2709 1543
rect 2722 1523 2725 1596
rect 2738 1543 2741 1616
rect 2754 1393 2757 1416
rect 2586 1373 2605 1376
rect 2654 1373 2661 1376
rect 2610 1256 2613 1336
rect 2610 1253 2621 1256
rect 2586 1133 2589 1216
rect 2618 1153 2621 1253
rect 2626 1213 2637 1216
rect 2594 1126 2597 1146
rect 2642 1133 2645 1326
rect 2654 1286 2657 1373
rect 2674 1323 2693 1326
rect 2654 1283 2661 1286
rect 2658 1236 2661 1283
rect 2654 1233 2661 1236
rect 2654 1176 2657 1233
rect 2654 1173 2661 1176
rect 2658 1156 2661 1173
rect 2658 1153 2669 1156
rect 2674 1153 2677 1206
rect 2650 1133 2653 1146
rect 2578 1123 2597 1126
rect 2466 923 2469 986
rect 2514 943 2517 1006
rect 2522 1003 2541 1006
rect 2550 1013 2557 1016
rect 2602 1013 2605 1126
rect 2642 1123 2653 1126
rect 2522 983 2525 1003
rect 2550 966 2553 1013
rect 2562 986 2565 1006
rect 2562 983 2569 986
rect 2534 963 2553 966
rect 2474 933 2485 936
rect 2474 913 2485 916
rect 2498 903 2501 936
rect 2522 923 2525 936
rect 2534 916 2537 963
rect 2530 913 2537 916
rect 2458 853 2485 856
rect 2386 813 2405 816
rect 2378 803 2397 806
rect 2362 793 2373 796
rect 2362 743 2365 793
rect 2354 723 2365 726
rect 2370 723 2389 726
rect 2346 713 2357 716
rect 2346 683 2349 713
rect 2362 706 2365 723
rect 2354 703 2365 706
rect 2334 673 2341 676
rect 2306 593 2309 606
rect 2338 603 2341 673
rect 2354 576 2357 703
rect 2394 626 2397 803
rect 2410 726 2413 836
rect 2418 813 2421 826
rect 2434 803 2437 816
rect 2426 733 2429 746
rect 2450 736 2453 816
rect 2474 813 2477 846
rect 2434 733 2453 736
rect 2466 736 2469 806
rect 2482 746 2485 853
rect 2530 826 2533 913
rect 2546 886 2549 956
rect 2566 916 2569 983
rect 2578 923 2581 946
rect 2566 913 2589 916
rect 2594 913 2597 1006
rect 2618 943 2621 956
rect 2602 933 2621 936
rect 2546 883 2565 886
rect 2506 823 2533 826
rect 2506 806 2509 823
rect 2538 813 2541 826
rect 2482 743 2489 746
rect 2466 733 2477 736
rect 2410 723 2421 726
rect 2418 656 2421 723
rect 2418 653 2425 656
rect 2394 623 2401 626
rect 2378 596 2381 606
rect 2374 593 2381 596
rect 2386 593 2389 616
rect 2298 573 2305 576
rect 2354 573 2365 576
rect 2282 503 2293 506
rect 2282 426 2285 503
rect 2302 496 2305 573
rect 2330 563 2357 566
rect 2330 556 2333 563
rect 2314 553 2333 556
rect 2314 533 2317 553
rect 2298 493 2305 496
rect 2282 423 2293 426
rect 2282 393 2285 406
rect 2266 383 2285 386
rect 2202 343 2221 346
rect 2242 343 2269 346
rect 2106 213 2109 226
rect 2034 123 2037 176
rect 2050 143 2053 206
rect 2114 203 2117 216
rect 2138 203 2141 246
rect 2202 213 2205 343
rect 2250 333 2261 336
rect 2210 313 2213 326
rect 2250 306 2253 326
rect 2242 303 2253 306
rect 2242 216 2245 303
rect 2258 216 2261 333
rect 2266 306 2269 343
rect 2282 313 2285 383
rect 2290 376 2293 423
rect 2298 413 2301 493
rect 2330 486 2333 536
rect 2354 523 2357 563
rect 2362 486 2365 573
rect 2330 483 2365 486
rect 2374 476 2377 593
rect 2398 486 2401 623
rect 2422 606 2425 653
rect 2434 643 2437 726
rect 2434 613 2437 626
rect 2442 613 2445 656
rect 2450 613 2453 726
rect 2458 723 2469 726
rect 2458 713 2469 716
rect 2466 693 2469 713
rect 2466 623 2469 646
rect 2474 623 2477 733
rect 2486 696 2489 743
rect 2498 733 2501 806
rect 2506 803 2517 806
rect 2546 803 2549 816
rect 2514 746 2517 803
rect 2506 743 2517 746
rect 2482 693 2489 696
rect 2482 606 2485 693
rect 2490 673 2501 676
rect 2498 623 2501 673
rect 2422 603 2445 606
rect 2418 533 2421 546
rect 2410 506 2413 526
rect 2410 503 2421 506
rect 2370 473 2377 476
rect 2394 483 2401 486
rect 2306 403 2309 426
rect 2314 403 2317 416
rect 2298 393 2349 396
rect 2290 373 2301 376
rect 2266 303 2285 306
rect 2242 213 2253 216
rect 2258 213 2269 216
rect 2274 213 2277 226
rect 2218 193 2221 206
rect 2138 163 2181 166
rect 2138 133 2141 163
rect 2138 113 2141 126
rect 2154 123 2157 136
rect 2178 123 2181 163
rect 2250 143 2253 213
rect 2258 193 2261 206
rect 2266 196 2269 213
rect 2282 203 2285 303
rect 2298 226 2301 373
rect 2290 223 2301 226
rect 2290 203 2293 223
rect 2266 193 2285 196
rect 2282 183 2285 193
rect 2266 133 2269 176
rect 2322 173 2325 376
rect 2346 323 2349 393
rect 2362 363 2365 396
rect 2370 346 2373 473
rect 2394 393 2397 483
rect 2418 446 2421 503
rect 2410 443 2421 446
rect 2410 423 2413 443
rect 2426 413 2429 426
rect 2434 383 2437 406
rect 2362 343 2373 346
rect 2362 286 2365 343
rect 2362 283 2373 286
rect 2370 243 2373 283
rect 2338 193 2341 216
rect 1578 83 1605 86
rect 2250 86 2253 126
rect 2290 86 2293 126
rect 2346 123 2349 146
rect 2354 143 2357 186
rect 2386 123 2389 146
rect 2402 133 2405 326
rect 2426 316 2429 326
rect 2426 313 2437 316
rect 2442 306 2445 603
rect 2474 533 2477 606
rect 2482 603 2493 606
rect 2490 526 2493 603
rect 2482 523 2493 526
rect 2458 373 2461 406
rect 2482 316 2485 523
rect 2506 456 2509 743
rect 2538 733 2541 746
rect 2530 713 2533 726
rect 2546 676 2549 726
rect 2538 673 2549 676
rect 2554 626 2557 806
rect 2562 723 2565 883
rect 2570 716 2573 886
rect 2566 713 2573 716
rect 2566 636 2569 713
rect 2522 623 2557 626
rect 2562 633 2569 636
rect 2530 613 2533 623
rect 2554 573 2557 606
rect 2502 453 2509 456
rect 2490 383 2493 416
rect 2502 396 2505 453
rect 2538 413 2541 546
rect 2554 506 2557 526
rect 2562 523 2565 633
rect 2570 516 2573 616
rect 2578 603 2581 906
rect 2586 896 2589 913
rect 2602 903 2605 933
rect 2626 903 2629 926
rect 2586 893 2593 896
rect 2634 893 2637 926
rect 2590 826 2593 893
rect 2586 823 2593 826
rect 2586 716 2589 823
rect 2602 813 2605 836
rect 2610 823 2621 826
rect 2626 813 2629 826
rect 2642 813 2645 1123
rect 2666 976 2669 1153
rect 2714 1133 2717 1216
rect 2754 1213 2757 1256
rect 2650 973 2669 976
rect 2706 976 2709 1126
rect 2706 973 2717 976
rect 2650 886 2653 973
rect 2658 963 2701 966
rect 2658 933 2661 963
rect 2658 903 2661 916
rect 2650 883 2657 886
rect 2594 733 2597 806
rect 2618 793 2621 806
rect 2626 733 2629 746
rect 2586 713 2597 716
rect 2594 646 2597 713
rect 2610 696 2613 726
rect 2618 723 2629 726
rect 2618 713 2621 723
rect 2626 703 2629 716
rect 2642 696 2645 806
rect 2654 706 2657 883
rect 2674 803 2677 936
rect 2698 923 2701 963
rect 2714 916 2717 973
rect 2706 913 2717 916
rect 2754 913 2757 926
rect 2698 793 2701 816
rect 2706 803 2709 913
rect 2754 813 2757 826
rect 2654 703 2669 706
rect 2610 693 2645 696
rect 2586 643 2597 646
rect 2586 613 2589 643
rect 2602 593 2605 606
rect 2634 533 2637 616
rect 2666 576 2669 703
rect 2674 603 2677 776
rect 2698 723 2701 746
rect 2754 713 2757 726
rect 2682 613 2685 626
rect 2722 623 2741 626
rect 2722 613 2725 623
rect 2690 593 2693 606
rect 2722 593 2725 606
rect 2730 603 2733 616
rect 2738 596 2741 623
rect 2730 593 2741 596
rect 2754 593 2757 606
rect 2666 573 2709 576
rect 2570 513 2581 516
rect 2554 503 2597 506
rect 2546 413 2549 426
rect 2502 393 2509 396
rect 2546 393 2549 406
rect 2570 403 2573 416
rect 2594 413 2597 503
rect 2650 393 2653 416
rect 2666 403 2669 573
rect 2682 536 2685 546
rect 2682 533 2701 536
rect 2698 426 2701 526
rect 2706 523 2709 573
rect 2730 523 2733 593
rect 2754 533 2757 546
rect 2698 423 2709 426
rect 2506 373 2509 393
rect 2690 376 2693 416
rect 2658 373 2693 376
rect 2570 343 2597 346
rect 2514 333 2525 336
rect 2490 323 2517 326
rect 2434 293 2437 306
rect 2442 303 2453 306
rect 2458 226 2461 316
rect 2466 293 2469 306
rect 2450 223 2461 226
rect 2450 213 2453 223
rect 2458 206 2461 216
rect 2466 213 2469 226
rect 2458 203 2469 206
rect 2474 133 2477 316
rect 2482 313 2509 316
rect 2530 306 2533 326
rect 2498 303 2533 306
rect 2498 226 2501 303
rect 2494 223 2501 226
rect 2482 133 2485 186
rect 2494 166 2497 223
rect 2490 163 2497 166
rect 2410 113 2413 126
rect 2482 116 2485 126
rect 2490 123 2493 163
rect 2498 116 2501 136
rect 2506 126 2509 206
rect 2514 133 2517 226
rect 2522 133 2525 303
rect 2530 213 2533 236
rect 2538 213 2541 336
rect 2546 223 2549 246
rect 2554 203 2557 256
rect 2570 183 2573 343
rect 2578 313 2581 326
rect 2586 316 2589 336
rect 2594 333 2597 343
rect 2626 326 2629 346
rect 2626 323 2637 326
rect 2658 323 2661 373
rect 2586 313 2621 316
rect 2634 276 2637 323
rect 2578 223 2581 236
rect 2538 133 2541 146
rect 2506 123 2525 126
rect 2482 113 2501 116
rect 2594 113 2597 156
rect 2602 143 2605 206
rect 2618 203 2621 276
rect 2626 273 2637 276
rect 2674 273 2677 366
rect 2706 296 2709 423
rect 2730 413 2749 416
rect 2730 376 2733 413
rect 2722 373 2733 376
rect 2722 323 2725 373
rect 2754 323 2757 336
rect 2698 293 2709 296
rect 2626 253 2629 273
rect 2698 236 2701 293
rect 2694 233 2701 236
rect 2658 143 2661 216
rect 2694 176 2697 233
rect 2706 213 2709 226
rect 2674 173 2697 176
rect 2602 123 2621 126
rect 2250 83 2293 86
rect 2658 86 2661 136
rect 2674 123 2677 173
rect 2698 86 2701 126
rect 2754 123 2757 146
rect 2658 83 2701 86
rect 2774 37 2794 2603
rect 2798 13 2818 2627
<< metal3 >>
rect 1201 2602 1630 2607
rect 945 2592 1110 2597
rect 417 2582 902 2587
rect 417 2567 422 2582
rect 897 2567 902 2582
rect 945 2567 950 2592
rect 1105 2587 1110 2592
rect 1201 2587 1206 2602
rect 1625 2597 1630 2602
rect 1625 2592 1718 2597
rect 1713 2587 1718 2592
rect 1105 2582 1206 2587
rect 1225 2582 1590 2587
rect 1713 2582 1742 2587
rect 1225 2577 1230 2582
rect 1193 2572 1230 2577
rect 1585 2577 1590 2582
rect 1585 2572 1614 2577
rect 1249 2567 1358 2572
rect 393 2562 422 2567
rect 569 2562 742 2567
rect 897 2562 950 2567
rect 1153 2562 1254 2567
rect 1353 2562 1758 2567
rect 569 2557 574 2562
rect 401 2552 486 2557
rect 545 2552 574 2557
rect 737 2557 742 2562
rect 1153 2557 1158 2562
rect 737 2552 1158 2557
rect 1169 2552 1238 2557
rect 1281 2552 1510 2557
rect 1585 2552 1630 2557
rect 1649 2552 1774 2557
rect 2105 2552 2190 2557
rect 2209 2552 2406 2557
rect 1169 2547 1174 2552
rect 2105 2547 2110 2552
rect 457 2542 662 2547
rect 689 2542 734 2547
rect 945 2542 1014 2547
rect 1113 2542 1174 2547
rect 1185 2542 1278 2547
rect 1545 2542 1710 2547
rect 1993 2542 2110 2547
rect 2185 2547 2190 2552
rect 2185 2542 2294 2547
rect 657 2537 662 2542
rect 945 2537 950 2542
rect 1009 2537 1118 2542
rect 1185 2537 1190 2542
rect 1297 2537 1526 2542
rect 473 2532 574 2537
rect 657 2532 718 2537
rect 865 2532 950 2537
rect 961 2532 982 2537
rect 1137 2532 1190 2537
rect 1265 2532 1302 2537
rect 1521 2532 1622 2537
rect 1793 2532 1910 2537
rect 1985 2532 2174 2537
rect 961 2527 966 2532
rect 1681 2527 1798 2532
rect 329 2522 526 2527
rect 521 2517 526 2522
rect 585 2522 678 2527
rect 809 2522 966 2527
rect 985 2522 1054 2527
rect 1113 2522 1510 2527
rect 1633 2522 1686 2527
rect 585 2517 590 2522
rect 521 2512 590 2517
rect 673 2512 678 2522
rect 1505 2517 1638 2522
rect 1905 2517 1910 2532
rect 2169 2527 2174 2532
rect 2305 2532 2390 2537
rect 2449 2532 2518 2537
rect 2577 2532 2678 2537
rect 2305 2527 2310 2532
rect 2169 2522 2310 2527
rect 689 2512 1198 2517
rect 1249 2512 1398 2517
rect 1457 2512 1486 2517
rect 1697 2512 1750 2517
rect 1817 2512 1894 2517
rect 1905 2512 1998 2517
rect 689 2507 694 2512
rect 641 2502 694 2507
rect 713 2502 1222 2507
rect 1305 2502 1374 2507
rect 1433 2502 1670 2507
rect 1705 2502 1814 2507
rect 1825 2502 1854 2507
rect 1865 2502 1926 2507
rect 2097 2502 2486 2507
rect 2521 2502 2590 2507
rect 2601 2502 2702 2507
rect 1825 2497 1830 2502
rect 577 2492 806 2497
rect 817 2492 998 2497
rect 1201 2492 1582 2497
rect 1825 2492 1934 2497
rect 817 2487 822 2492
rect 1017 2487 1182 2492
rect 1689 2487 1806 2492
rect 489 2482 566 2487
rect 649 2482 822 2487
rect 881 2482 1022 2487
rect 1177 2482 1550 2487
rect 1665 2482 1694 2487
rect 1801 2482 1846 2487
rect 1857 2482 1982 2487
rect 2281 2482 2558 2487
rect 561 2477 654 2482
rect 1857 2477 1862 2482
rect 2553 2477 2558 2482
rect 2633 2482 2662 2487
rect 2633 2477 2638 2482
rect 769 2472 1262 2477
rect 1281 2472 1502 2477
rect 1601 2472 1862 2477
rect 1873 2472 1998 2477
rect 2017 2472 2094 2477
rect 2553 2472 2638 2477
rect 1281 2467 1286 2472
rect 2017 2467 2022 2472
rect 345 2462 470 2467
rect 345 2457 350 2462
rect 321 2452 350 2457
rect 465 2457 470 2462
rect 505 2462 750 2467
rect 801 2462 910 2467
rect 1025 2462 1286 2467
rect 1329 2462 1910 2467
rect 1993 2462 2022 2467
rect 2089 2467 2094 2472
rect 2089 2462 2270 2467
rect 505 2457 510 2462
rect 465 2452 510 2457
rect 745 2457 750 2462
rect 905 2457 1030 2462
rect 1905 2457 1998 2462
rect 745 2452 886 2457
rect 1049 2452 1294 2457
rect 1329 2452 1414 2457
rect 1521 2452 1886 2457
rect 2265 2447 2270 2462
rect 2425 2462 2454 2467
rect 2425 2447 2430 2462
rect 521 2442 1694 2447
rect 1849 2442 2078 2447
rect 2265 2442 2430 2447
rect 281 2437 422 2442
rect 1713 2437 1822 2442
rect 193 2432 286 2437
rect 417 2432 470 2437
rect 513 2432 558 2437
rect 745 2432 838 2437
rect 1025 2432 1310 2437
rect 1385 2432 1486 2437
rect 1553 2432 1718 2437
rect 1817 2432 1846 2437
rect 1889 2432 1974 2437
rect 2537 2432 2670 2437
rect 297 2422 550 2427
rect 577 2422 710 2427
rect 729 2422 766 2427
rect 785 2422 1014 2427
rect 1129 2422 1158 2427
rect 1169 2422 1198 2427
rect 1321 2422 1902 2427
rect 1929 2422 2038 2427
rect 2649 2422 2742 2427
rect 577 2417 582 2422
rect 265 2412 294 2417
rect 289 2407 294 2412
rect 465 2412 494 2417
rect 505 2412 582 2417
rect 705 2417 710 2422
rect 785 2417 790 2422
rect 1009 2417 1134 2422
rect 1193 2417 1326 2422
rect 705 2412 790 2417
rect 1369 2412 2102 2417
rect 465 2407 470 2412
rect 169 2402 230 2407
rect 289 2402 470 2407
rect 529 2402 534 2412
rect 809 2407 982 2412
rect 585 2402 814 2407
rect 977 2402 1358 2407
rect 1425 2402 1454 2407
rect 1913 2402 2086 2407
rect 1353 2397 1430 2402
rect 1561 2397 1694 2402
rect 1753 2397 1862 2402
rect 129 2392 190 2397
rect 513 2392 614 2397
rect 665 2392 966 2397
rect 1081 2392 1110 2397
rect 1537 2392 1566 2397
rect 1689 2392 1758 2397
rect 1857 2392 1886 2397
rect 1969 2392 2070 2397
rect 2081 2392 2086 2402
rect 2657 2402 2734 2407
rect 2657 2397 2662 2402
rect 2497 2392 2550 2397
rect 2625 2392 2662 2397
rect 2729 2397 2734 2402
rect 2729 2392 2758 2397
rect 961 2387 1086 2392
rect 1185 2387 1278 2392
rect 1969 2387 1974 2392
rect 161 2382 246 2387
rect 257 2382 414 2387
rect 721 2382 822 2387
rect 841 2382 942 2387
rect 1161 2382 1190 2387
rect 1273 2382 1678 2387
rect 1769 2382 1974 2387
rect 2673 2382 2726 2387
rect 505 2377 694 2382
rect 817 2377 822 2382
rect 385 2372 510 2377
rect 689 2372 742 2377
rect 817 2372 934 2377
rect 961 2372 1134 2377
rect 1153 2372 1262 2377
rect 1449 2372 1574 2377
rect 1705 2372 2038 2377
rect 737 2367 742 2372
rect 961 2367 966 2372
rect 521 2362 694 2367
rect 737 2362 966 2367
rect 1129 2367 1134 2372
rect 1129 2362 1158 2367
rect 1217 2362 1414 2367
rect 1593 2362 1686 2367
rect 2113 2362 2190 2367
rect 2409 2362 2526 2367
rect 689 2357 694 2362
rect 1217 2357 1222 2362
rect 1593 2357 1598 2362
rect 305 2352 374 2357
rect 369 2347 374 2352
rect 433 2352 670 2357
rect 689 2352 982 2357
rect 993 2352 1222 2357
rect 1393 2352 1598 2357
rect 1681 2357 1686 2362
rect 1737 2357 1958 2362
rect 1681 2352 1742 2357
rect 1953 2352 2046 2357
rect 2633 2352 2710 2357
rect 433 2347 438 2352
rect 2481 2347 2590 2352
rect 369 2342 438 2347
rect 457 2342 750 2347
rect 969 2342 1054 2347
rect 1281 2342 1350 2347
rect 1369 2342 1478 2347
rect 1585 2342 1670 2347
rect 1753 2342 1846 2347
rect 1857 2342 1942 2347
rect 2201 2342 2294 2347
rect 2369 2342 2486 2347
rect 2585 2342 2702 2347
rect 769 2337 950 2342
rect 1665 2337 1758 2342
rect 1841 2337 1846 2342
rect 465 2332 582 2337
rect 617 2332 774 2337
rect 945 2332 1094 2337
rect 1337 2332 1454 2337
rect 1841 2332 1950 2337
rect 2025 2332 2142 2337
rect 2169 2332 2358 2337
rect 2505 2332 2582 2337
rect 577 2327 582 2332
rect 1473 2327 1622 2332
rect 561 2317 566 2327
rect 577 2322 1086 2327
rect 1113 2322 1214 2327
rect 1233 2322 1478 2327
rect 1617 2322 1942 2327
rect 2001 2322 2102 2327
rect 2121 2322 2502 2327
rect 2593 2322 2622 2327
rect 1113 2317 1118 2322
rect 337 2312 510 2317
rect 529 2312 1118 2317
rect 1209 2317 1214 2322
rect 2097 2317 2102 2322
rect 2497 2317 2502 2322
rect 2617 2317 2622 2322
rect 2681 2322 2710 2327
rect 2681 2317 2686 2322
rect 1209 2312 1606 2317
rect 1825 2312 1862 2317
rect 2097 2312 2126 2317
rect 2241 2312 2350 2317
rect 529 2307 534 2312
rect 377 2302 534 2307
rect 545 2302 934 2307
rect 1033 2302 1374 2307
rect 1425 2302 1494 2307
rect 1521 2302 1590 2307
rect 1609 2302 1678 2307
rect 1825 2302 1830 2312
rect 2121 2307 2230 2312
rect 2345 2307 2350 2312
rect 2433 2312 2462 2317
rect 2497 2312 2542 2317
rect 2617 2312 2686 2317
rect 2433 2307 2438 2312
rect 2225 2302 2326 2307
rect 2345 2302 2438 2307
rect 929 2297 1038 2302
rect 1521 2297 1526 2302
rect 457 2292 574 2297
rect 665 2292 726 2297
rect 841 2292 910 2297
rect 1057 2292 1358 2297
rect 1377 2292 1422 2297
rect 1441 2292 1526 2297
rect 1705 2292 1806 2297
rect 2105 2292 2222 2297
rect 393 2282 414 2287
rect 705 2282 862 2287
rect 1001 2282 1054 2287
rect 1129 2282 1334 2287
rect 1449 2282 1726 2287
rect 1849 2282 1918 2287
rect 1849 2277 1854 2282
rect 417 2272 1230 2277
rect 1305 2272 1550 2277
rect 1729 2272 1854 2277
rect 1913 2277 1918 2282
rect 1913 2272 1990 2277
rect 2017 2272 2134 2277
rect 2129 2267 2134 2272
rect 2233 2272 2566 2277
rect 2233 2267 2238 2272
rect 1057 2262 1790 2267
rect 1817 2262 2110 2267
rect 2129 2262 2238 2267
rect 473 2257 558 2262
rect 849 2257 1014 2262
rect 1057 2257 1062 2262
rect 449 2252 478 2257
rect 553 2252 854 2257
rect 1009 2252 1062 2257
rect 1081 2252 1510 2257
rect 1665 2252 1990 2257
rect 417 2242 542 2247
rect 865 2242 1606 2247
rect 1641 2242 1670 2247
rect 1809 2242 1854 2247
rect 2001 2242 2030 2247
rect 1689 2237 1758 2242
rect 1849 2237 2006 2242
rect 409 2232 502 2237
rect 529 2232 574 2237
rect 593 2232 742 2237
rect 761 2232 886 2237
rect 985 2232 1694 2237
rect 1753 2232 1830 2237
rect 497 2227 502 2232
rect 593 2227 598 2232
rect 145 2222 182 2227
rect 385 2222 414 2227
rect 425 2222 478 2227
rect 497 2222 598 2227
rect 737 2227 742 2232
rect 737 2222 822 2227
rect 833 2222 862 2227
rect 897 2222 1174 2227
rect 1225 2222 1510 2227
rect 1633 2222 1742 2227
rect 1833 2222 1886 2227
rect 1913 2222 1998 2227
rect 2057 2222 2126 2227
rect 2601 2222 2654 2227
rect 817 2217 822 2222
rect 161 2212 214 2217
rect 369 2212 510 2217
rect 609 2212 790 2217
rect 817 2212 990 2217
rect 1097 2212 1142 2217
rect 505 2207 614 2212
rect 1169 2207 1174 2222
rect 1185 2212 1630 2217
rect 1649 2212 1830 2217
rect 2049 2212 2134 2217
rect 2473 2212 2686 2217
rect 1825 2207 2054 2212
rect 2473 2207 2478 2212
rect 313 2202 358 2207
rect 465 2202 486 2207
rect 673 2202 734 2207
rect 897 2202 1158 2207
rect 1169 2202 1190 2207
rect 1209 2202 1334 2207
rect 1529 2202 1566 2207
rect 2073 2202 2174 2207
rect 2313 2202 2398 2207
rect 2417 2202 2478 2207
rect 1185 2197 1190 2202
rect 1345 2197 1534 2202
rect 1721 2197 1806 2202
rect 2313 2197 2318 2202
rect 273 2192 414 2197
rect 473 2192 542 2197
rect 601 2192 774 2197
rect 1185 2192 1350 2197
rect 1553 2192 1726 2197
rect 1801 2192 1830 2197
rect 1945 2192 2086 2197
rect 2289 2192 2318 2197
rect 2393 2197 2398 2202
rect 2393 2192 2598 2197
rect 2641 2192 2678 2197
rect 969 2187 1166 2192
rect 185 2182 310 2187
rect 609 2182 710 2187
rect 841 2182 894 2187
rect 945 2182 974 2187
rect 1161 2182 1222 2187
rect 1233 2182 1590 2187
rect 1737 2182 1774 2187
rect 1969 2182 2022 2187
rect 2321 2182 2478 2187
rect 2545 2182 2574 2187
rect 2657 2182 2726 2187
rect 729 2177 822 2182
rect 1233 2177 1238 2182
rect 1585 2177 1590 2182
rect 2041 2177 2142 2182
rect 217 2172 334 2177
rect 505 2172 598 2177
rect 593 2167 598 2172
rect 681 2172 734 2177
rect 817 2172 1238 2177
rect 1529 2172 1574 2177
rect 1585 2172 1734 2177
rect 1745 2172 2046 2177
rect 2137 2172 2166 2177
rect 681 2167 686 2172
rect 1257 2167 1510 2172
rect 369 2162 438 2167
rect 593 2162 686 2167
rect 705 2162 806 2167
rect 857 2162 1022 2167
rect 1105 2162 1262 2167
rect 1505 2162 1646 2167
rect 1961 2162 2134 2167
rect 2153 2162 2230 2167
rect 1017 2157 1110 2162
rect 241 2152 542 2157
rect 897 2152 942 2157
rect 977 2152 998 2157
rect 1129 2152 1294 2157
rect 1313 2152 1334 2157
rect 1369 2152 1582 2157
rect 1945 2152 2070 2157
rect 121 2142 174 2147
rect 217 2142 246 2147
rect 337 2142 366 2147
rect 441 2142 534 2147
rect 601 2142 654 2147
rect 681 2142 718 2147
rect 241 2137 342 2142
rect 897 2137 902 2152
rect 945 2142 982 2147
rect 641 2132 670 2137
rect 729 2132 902 2137
rect 665 2127 734 2132
rect 993 2127 998 2152
rect 1313 2147 1318 2152
rect 1017 2142 1142 2147
rect 1137 2137 1142 2142
rect 1217 2142 1438 2147
rect 1449 2142 1574 2147
rect 1665 2142 1798 2147
rect 1985 2142 2038 2147
rect 2049 2142 2126 2147
rect 2433 2142 2518 2147
rect 2593 2142 2622 2147
rect 1217 2137 1222 2142
rect 1665 2137 1670 2142
rect 1137 2132 1222 2137
rect 1297 2132 1670 2137
rect 1793 2137 1798 2142
rect 2033 2137 2038 2142
rect 2513 2137 2518 2142
rect 2641 2137 2646 2147
rect 2665 2142 2734 2147
rect 1793 2132 1822 2137
rect 1913 2132 1982 2137
rect 2033 2132 2118 2137
rect 2513 2132 2646 2137
rect 289 2122 342 2127
rect 577 2122 630 2127
rect 865 2122 934 2127
rect 977 2122 998 2127
rect 1073 2122 1118 2127
rect 1481 2122 1574 2127
rect 1793 2122 1846 2127
rect 1361 2117 1430 2122
rect 641 2112 854 2117
rect 993 2112 1366 2117
rect 1425 2112 2262 2117
rect 2281 2112 2454 2117
rect 2553 2112 2646 2117
rect 473 2107 646 2112
rect 849 2107 998 2112
rect 385 2102 478 2107
rect 1017 2102 1046 2107
rect 1105 2102 1182 2107
rect 1377 2102 1670 2107
rect 1713 2102 1790 2107
rect 1817 2102 2070 2107
rect 2105 2102 2174 2107
rect 1201 2097 1358 2102
rect 513 2092 654 2097
rect 825 2092 910 2097
rect 1081 2092 1206 2097
rect 1353 2092 1446 2097
rect 1721 2092 1902 2097
rect 1937 2092 1966 2097
rect 825 2087 830 2092
rect 537 2082 622 2087
rect 689 2082 830 2087
rect 905 2087 910 2092
rect 1441 2087 1702 2092
rect 905 2082 934 2087
rect 1009 2082 1302 2087
rect 1313 2082 1422 2087
rect 1697 2082 2030 2087
rect 841 2072 1646 2077
rect 1681 2072 1958 2077
rect 2041 2072 2134 2077
rect 1953 2067 2046 2072
rect 1145 2062 1262 2067
rect 1609 2062 1934 2067
rect 2577 2062 2670 2067
rect 857 2057 1054 2062
rect 1281 2057 1414 2062
rect 833 2052 862 2057
rect 1049 2052 1286 2057
rect 1409 2052 1438 2057
rect 1457 2052 1894 2057
rect 1929 2052 1998 2057
rect 2529 2052 2582 2057
rect 1457 2047 1462 2052
rect 785 2042 1038 2047
rect 1153 2042 1462 2047
rect 1585 2042 1782 2047
rect 1849 2042 1870 2047
rect 1881 2042 2014 2047
rect 1033 2037 1158 2042
rect 361 2032 422 2037
rect 673 2032 1014 2037
rect 1177 2032 1838 2037
rect 1977 2032 2022 2037
rect 1833 2027 1982 2032
rect 393 2022 438 2027
rect 481 2022 806 2027
rect 865 2022 1006 2027
rect 1065 2017 1070 2027
rect 1153 2022 1342 2027
rect 1353 2022 1430 2027
rect 1553 2022 1806 2027
rect 2017 2022 2022 2032
rect 2569 2022 2630 2027
rect 2625 2017 2630 2022
rect 273 2012 438 2017
rect 433 2007 438 2012
rect 521 2012 550 2017
rect 657 2012 886 2017
rect 1065 2012 1318 2017
rect 1441 2012 1614 2017
rect 1625 2012 1702 2017
rect 1897 2012 1982 2017
rect 2409 2012 2478 2017
rect 2601 2012 2630 2017
rect 521 2007 526 2012
rect 905 2007 982 2012
rect 225 2002 310 2007
rect 321 2002 382 2007
rect 433 2002 526 2007
rect 745 2002 790 2007
rect 809 2002 910 2007
rect 977 2002 1054 2007
rect 1113 2002 1718 2007
rect 1729 2002 1838 2007
rect 1049 1997 1118 2002
rect 1937 1997 1942 2012
rect 1985 2002 2070 2007
rect 2345 2002 2454 2007
rect 2657 1997 2662 2027
rect 217 1992 254 1997
rect 329 1992 414 1997
rect 601 1992 670 1997
rect 897 1992 966 1997
rect 1137 1992 1278 1997
rect 1361 1992 1430 1997
rect 1505 1992 1542 1997
rect 1937 1992 1966 1997
rect 2057 1992 2134 1997
rect 2225 1992 2286 1997
rect 2433 1992 2478 1997
rect 2601 1992 2742 1997
rect 601 1987 606 1992
rect 297 1982 390 1987
rect 433 1982 606 1987
rect 665 1987 670 1992
rect 1561 1987 1654 1992
rect 665 1982 694 1987
rect 817 1982 1030 1987
rect 1073 1982 1566 1987
rect 1649 1982 1678 1987
rect 2649 1982 2686 1987
rect 337 1972 478 1977
rect 617 1972 766 1977
rect 809 1972 854 1977
rect 937 1972 1086 1977
rect 1193 1972 1262 1977
rect 1353 1972 1422 1977
rect 1433 1972 1550 1977
rect 1593 1972 1630 1977
rect 1625 1967 1630 1972
rect 1689 1972 1830 1977
rect 1689 1967 1694 1972
rect 257 1962 558 1967
rect 577 1962 886 1967
rect 913 1962 958 1967
rect 993 1962 1254 1967
rect 1297 1962 1518 1967
rect 1625 1962 1694 1967
rect 297 1952 510 1957
rect 625 1952 1166 1957
rect 1417 1952 1606 1957
rect 1785 1952 1870 1957
rect 1889 1952 2054 1957
rect 1161 1947 1422 1952
rect 1889 1947 1894 1952
rect 2657 1947 2662 1957
rect 185 1942 214 1947
rect 265 1942 534 1947
rect 641 1942 822 1947
rect 1001 1942 1142 1947
rect 1441 1942 1518 1947
rect 1617 1942 1718 1947
rect 1729 1942 1894 1947
rect 2017 1942 2046 1947
rect 2129 1942 2214 1947
rect 2233 1942 2302 1947
rect 2369 1942 2454 1947
rect 2633 1942 2662 1947
rect 2673 1942 2726 1947
rect 841 1937 982 1942
rect 1617 1937 1622 1942
rect 177 1932 262 1937
rect 417 1932 438 1937
rect 609 1932 846 1937
rect 977 1932 1622 1937
rect 1713 1937 1718 1942
rect 2233 1937 2238 1942
rect 1713 1932 2006 1937
rect 2177 1932 2238 1937
rect 2297 1937 2302 1942
rect 2297 1932 2326 1937
rect 2601 1932 2734 1937
rect 225 1912 230 1932
rect 433 1927 438 1932
rect 249 1922 318 1927
rect 417 1922 438 1927
rect 481 1922 630 1927
rect 745 1922 790 1927
rect 825 1922 958 1927
rect 985 1922 1022 1927
rect 1041 1922 1078 1927
rect 1089 1922 1350 1927
rect 1969 1922 2118 1927
rect 2145 1922 2206 1927
rect 2281 1922 2398 1927
rect 2537 1922 2590 1927
rect 417 1912 422 1922
rect 1041 1917 1046 1922
rect 1761 1917 1894 1922
rect 521 1912 1046 1917
rect 1289 1912 1766 1917
rect 1889 1912 1950 1917
rect 2225 1912 2254 1917
rect 2569 1912 2598 1917
rect 1057 1907 1294 1912
rect 2065 1907 2230 1912
rect 2593 1907 2598 1912
rect 2665 1912 2710 1917
rect 2665 1907 2670 1912
rect 209 1902 302 1907
rect 337 1902 478 1907
rect 489 1902 542 1907
rect 625 1902 1062 1907
rect 1313 1902 1342 1907
rect 1777 1902 1878 1907
rect 625 1897 630 1902
rect 1361 1897 1710 1902
rect 2065 1897 2070 1907
rect 2593 1902 2670 1907
rect 2689 1902 2734 1907
rect 185 1892 214 1897
rect 209 1877 214 1892
rect 473 1892 630 1897
rect 665 1892 846 1897
rect 1081 1892 1206 1897
rect 473 1877 478 1892
rect 865 1887 1086 1892
rect 1201 1887 1206 1892
rect 1297 1892 1366 1897
rect 1705 1892 1766 1897
rect 1889 1892 2070 1897
rect 2081 1892 2214 1897
rect 2313 1892 2534 1897
rect 497 1882 614 1887
rect 689 1882 870 1887
rect 1201 1882 1230 1887
rect 1297 1877 1302 1892
rect 1761 1887 1894 1892
rect 1321 1882 1550 1887
rect 1577 1882 1694 1887
rect 209 1872 478 1877
rect 729 1872 862 1877
rect 873 1872 1302 1877
rect 1337 1872 1382 1877
rect 1393 1872 1438 1877
rect 1697 1872 1742 1877
rect 1809 1872 1878 1877
rect 873 1867 878 1872
rect 1809 1867 1814 1872
rect 569 1862 878 1867
rect 945 1862 1446 1867
rect 1537 1862 1814 1867
rect 1873 1867 1878 1872
rect 1873 1862 1902 1867
rect 2001 1862 2174 1867
rect 1537 1857 1542 1862
rect 761 1852 1166 1857
rect 1249 1852 1542 1857
rect 1681 1852 1790 1857
rect 1881 1852 1926 1857
rect 2529 1852 2662 1857
rect 1785 1847 1886 1852
rect 1945 1847 2118 1852
rect 665 1842 1766 1847
rect 1905 1842 1950 1847
rect 2113 1842 2238 1847
rect 2281 1842 2398 1847
rect 2577 1842 2734 1847
rect 1761 1837 1766 1842
rect 193 1832 222 1837
rect 633 1832 734 1837
rect 857 1832 1638 1837
rect 1689 1832 1750 1837
rect 1761 1832 2086 1837
rect 2273 1832 2302 1837
rect 729 1827 862 1832
rect 185 1822 262 1827
rect 393 1822 486 1827
rect 601 1822 710 1827
rect 1001 1822 1022 1827
rect 1049 1822 1166 1827
rect 1201 1822 1382 1827
rect 1497 1822 1550 1827
rect 1633 1822 1638 1832
rect 2121 1827 2254 1832
rect 1937 1822 1990 1827
rect 705 1817 710 1822
rect 881 1817 982 1822
rect 1377 1817 1502 1822
rect 1633 1817 1718 1822
rect 1985 1817 1990 1822
rect 2097 1822 2126 1827
rect 2249 1822 2366 1827
rect 2377 1822 2518 1827
rect 2545 1822 2622 1827
rect 2097 1817 2102 1822
rect 161 1812 198 1817
rect 233 1812 278 1817
rect 513 1812 590 1817
rect 585 1807 590 1812
rect 649 1812 686 1817
rect 705 1812 798 1817
rect 857 1812 886 1817
rect 977 1812 1358 1817
rect 1521 1812 1542 1817
rect 1553 1812 1614 1817
rect 1713 1812 1950 1817
rect 1985 1812 2102 1817
rect 2121 1812 2166 1817
rect 2177 1812 2230 1817
rect 2265 1812 2310 1817
rect 2537 1812 2638 1817
rect 649 1807 654 1812
rect 289 1802 334 1807
rect 585 1802 654 1807
rect 913 1802 1174 1807
rect 1233 1802 1966 1807
rect 2249 1802 2286 1807
rect 2569 1802 2710 1807
rect 673 1797 918 1802
rect 177 1792 278 1797
rect 385 1792 446 1797
rect 673 1777 678 1797
rect 937 1792 1150 1797
rect 1169 1792 1174 1802
rect 1289 1792 1366 1797
rect 1489 1792 1518 1797
rect 1625 1792 1670 1797
rect 1713 1792 1782 1797
rect 1793 1792 1886 1797
rect 1969 1792 2014 1797
rect 2081 1792 2150 1797
rect 745 1782 830 1787
rect 857 1782 1054 1787
rect 1089 1782 1158 1787
rect 1281 1782 1678 1787
rect 2049 1782 2078 1787
rect 745 1777 750 1782
rect 137 1772 214 1777
rect 417 1772 502 1777
rect 569 1772 678 1777
rect 689 1772 750 1777
rect 825 1777 830 1782
rect 1953 1777 2054 1782
rect 825 1772 950 1777
rect 1081 1772 1478 1777
rect 1649 1772 1958 1777
rect 689 1767 694 1772
rect 1473 1767 1590 1772
rect 1649 1767 1654 1772
rect 401 1762 694 1767
rect 761 1762 814 1767
rect 945 1762 1046 1767
rect 1121 1762 1206 1767
rect 1217 1762 1334 1767
rect 1425 1762 1454 1767
rect 1585 1762 1654 1767
rect 1745 1762 1766 1767
rect 1897 1762 1990 1767
rect 2001 1762 2126 1767
rect 2217 1762 2318 1767
rect 401 1757 406 1762
rect 1121 1757 1126 1762
rect 1329 1757 1430 1762
rect 345 1752 406 1757
rect 425 1752 1126 1757
rect 1145 1752 1310 1757
rect 1537 1752 1566 1757
rect 1921 1752 2062 1757
rect 2217 1752 2390 1757
rect 289 1742 486 1747
rect 545 1742 734 1747
rect 1025 1742 1118 1747
rect 1161 1742 1422 1747
rect 1545 1742 1942 1747
rect 1969 1742 2086 1747
rect 2113 1742 2134 1747
rect 2225 1742 2334 1747
rect 841 1737 966 1742
rect 2353 1737 2430 1742
rect 225 1732 414 1737
rect 537 1732 790 1737
rect 817 1732 846 1737
rect 961 1732 990 1737
rect 1177 1732 1262 1737
rect 1313 1732 1390 1737
rect 1873 1732 1982 1737
rect 2049 1732 2358 1737
rect 2425 1732 2558 1737
rect 2609 1732 2694 1737
rect 1009 1727 1142 1732
rect 593 1722 1014 1727
rect 1137 1722 1230 1727
rect 1409 1722 1566 1727
rect 1585 1722 1670 1727
rect 1801 1722 1902 1727
rect 2081 1722 2110 1727
rect 2209 1722 2246 1727
rect 2281 1722 2414 1727
rect 313 1717 430 1722
rect 1257 1717 1414 1722
rect 1561 1717 1566 1722
rect 1921 1717 2062 1722
rect 289 1712 318 1717
rect 425 1712 494 1717
rect 601 1712 702 1717
rect 793 1712 902 1717
rect 969 1712 1126 1717
rect 1233 1712 1262 1717
rect 1561 1712 1766 1717
rect 1785 1712 1926 1717
rect 2057 1712 2390 1717
rect 2665 1712 2742 1717
rect 1145 1707 1238 1712
rect 1761 1707 1766 1712
rect 2385 1707 2390 1712
rect 305 1702 334 1707
rect 377 1702 414 1707
rect 713 1702 1150 1707
rect 1257 1702 1726 1707
rect 1761 1702 1790 1707
rect 1889 1702 2094 1707
rect 2249 1702 2366 1707
rect 2385 1702 2422 1707
rect 1785 1697 1894 1702
rect 2129 1697 2230 1702
rect 449 1692 694 1697
rect 873 1692 1286 1697
rect 1617 1692 1662 1697
rect 2105 1692 2134 1697
rect 2225 1692 2294 1697
rect 713 1687 854 1692
rect 1305 1687 1598 1692
rect 441 1682 470 1687
rect 649 1682 718 1687
rect 849 1682 878 1687
rect 985 1682 1142 1687
rect 1225 1682 1310 1687
rect 1593 1682 1614 1687
rect 1673 1682 2278 1687
rect 465 1677 654 1682
rect 1609 1677 1678 1682
rect 185 1672 430 1677
rect 425 1667 430 1672
rect 673 1672 1182 1677
rect 1209 1672 1494 1677
rect 1553 1672 1582 1677
rect 673 1667 678 1672
rect 425 1662 678 1667
rect 697 1662 1086 1667
rect 1265 1662 1798 1667
rect 1873 1662 1958 1667
rect 1105 1657 1198 1662
rect 1265 1657 1270 1662
rect 1873 1657 1878 1662
rect 817 1652 1110 1657
rect 1193 1652 1270 1657
rect 1281 1652 1406 1657
rect 1473 1652 1614 1657
rect 1849 1652 1878 1657
rect 1953 1657 1958 1662
rect 2001 1662 2174 1667
rect 2001 1657 2006 1662
rect 1953 1652 2006 1657
rect 2169 1657 2174 1662
rect 2169 1652 2198 1657
rect 2217 1652 2350 1657
rect 1689 1647 1798 1652
rect 2217 1647 2222 1652
rect 377 1642 486 1647
rect 593 1642 654 1647
rect 665 1642 1694 1647
rect 1793 1642 2222 1647
rect 361 1632 606 1637
rect 849 1632 1238 1637
rect 1265 1632 1358 1637
rect 1369 1632 1510 1637
rect 1705 1632 1782 1637
rect 1897 1632 2014 1637
rect 2121 1632 2286 1637
rect 2681 1632 2718 1637
rect 641 1627 830 1632
rect 1617 1627 1686 1632
rect 2009 1627 2126 1632
rect 233 1622 550 1627
rect 585 1622 646 1627
rect 825 1622 1382 1627
rect 1505 1622 1622 1627
rect 1681 1622 1886 1627
rect 1401 1617 1510 1622
rect 1881 1617 1886 1622
rect 1961 1622 1990 1627
rect 2145 1622 2230 1627
rect 2305 1622 2382 1627
rect 2401 1622 2446 1627
rect 2497 1622 2550 1627
rect 1961 1617 1966 1622
rect 353 1612 422 1617
rect 657 1612 1406 1617
rect 1633 1612 1726 1617
rect 1825 1612 1846 1617
rect 1881 1612 1966 1617
rect 2041 1612 2262 1617
rect 2513 1612 2598 1617
rect 2609 1612 2726 1617
rect 521 1607 638 1612
rect 497 1602 526 1607
rect 633 1602 766 1607
rect 969 1602 998 1607
rect 1041 1602 1094 1607
rect 1161 1602 1214 1607
rect 1273 1602 1342 1607
rect 1377 1602 1494 1607
rect 1513 1602 1574 1607
rect 1601 1602 1622 1607
rect 1657 1602 1718 1607
rect 1761 1602 1822 1607
rect 369 1597 454 1602
rect 785 1597 886 1602
rect 1841 1597 1846 1612
rect 2113 1602 2214 1607
rect 2521 1602 2558 1607
rect 2113 1597 2118 1602
rect 2593 1597 2598 1612
rect 345 1592 374 1597
rect 449 1592 790 1597
rect 881 1592 1318 1597
rect 1441 1592 1790 1597
rect 1825 1592 1846 1597
rect 1905 1592 1942 1597
rect 1961 1592 2038 1597
rect 2089 1592 2118 1597
rect 2161 1592 2182 1597
rect 2257 1592 2550 1597
rect 2593 1592 2694 1597
rect 1313 1587 1446 1592
rect 2161 1587 2166 1592
rect 177 1582 334 1587
rect 329 1577 334 1582
rect 401 1582 438 1587
rect 641 1582 870 1587
rect 1025 1582 1078 1587
rect 1225 1582 1294 1587
rect 1465 1582 1630 1587
rect 1713 1582 1854 1587
rect 2025 1582 2062 1587
rect 2089 1582 2166 1587
rect 2177 1582 2222 1587
rect 2265 1582 2326 1587
rect 401 1577 406 1582
rect 497 1577 622 1582
rect 329 1572 406 1577
rect 473 1572 502 1577
rect 617 1572 694 1577
rect 689 1567 694 1572
rect 777 1572 1686 1577
rect 1697 1572 1742 1577
rect 777 1567 782 1572
rect 1681 1567 1686 1572
rect 2321 1567 2326 1582
rect 2489 1582 2518 1587
rect 2537 1582 2630 1587
rect 2489 1567 2494 1582
rect 425 1562 470 1567
rect 505 1562 638 1567
rect 689 1562 782 1567
rect 849 1562 1006 1567
rect 1233 1562 1278 1567
rect 1417 1562 1462 1567
rect 1473 1562 1494 1567
rect 1553 1562 1582 1567
rect 1681 1562 2030 1567
rect 2321 1562 2494 1567
rect 2513 1567 2518 1582
rect 2593 1572 2622 1577
rect 2593 1567 2598 1572
rect 2513 1562 2598 1567
rect 1025 1557 1142 1562
rect 1297 1557 1422 1562
rect 1457 1557 1462 1562
rect 353 1552 414 1557
rect 409 1547 414 1552
rect 473 1552 502 1557
rect 521 1552 662 1557
rect 801 1552 830 1557
rect 929 1552 1030 1557
rect 1137 1552 1166 1557
rect 1185 1552 1302 1557
rect 1457 1552 1662 1557
rect 1697 1552 1790 1557
rect 2073 1552 2110 1557
rect 2129 1552 2214 1557
rect 473 1547 478 1552
rect 825 1547 934 1552
rect 1697 1547 1702 1552
rect 2129 1547 2134 1552
rect 409 1542 478 1547
rect 593 1542 670 1547
rect 953 1542 1110 1547
rect 1121 1542 1174 1547
rect 1185 1542 1206 1547
rect 1321 1542 1430 1547
rect 1449 1542 1542 1547
rect 1625 1542 1702 1547
rect 1713 1542 1838 1547
rect 1849 1542 1878 1547
rect 2033 1542 2134 1547
rect 2209 1547 2214 1552
rect 2209 1542 2262 1547
rect 2561 1542 2742 1547
rect 593 1537 598 1542
rect 1225 1537 1326 1542
rect 1425 1537 1430 1542
rect 545 1532 598 1537
rect 609 1532 710 1537
rect 769 1532 862 1537
rect 1001 1532 1230 1537
rect 1425 1532 1494 1537
rect 1745 1532 1998 1537
rect 2145 1532 2198 1537
rect 1617 1527 1726 1532
rect 2145 1527 2150 1532
rect 689 1522 790 1527
rect 897 1522 1622 1527
rect 1721 1522 1814 1527
rect 2081 1522 2150 1527
rect 1953 1517 2062 1522
rect 273 1512 422 1517
rect 569 1512 1302 1517
rect 1521 1512 1958 1517
rect 2057 1512 2198 1517
rect 2625 1512 2678 1517
rect 1297 1507 1494 1512
rect 537 1502 574 1507
rect 649 1502 710 1507
rect 729 1502 814 1507
rect 889 1502 982 1507
rect 1001 1502 1038 1507
rect 1081 1502 1126 1507
rect 1169 1502 1206 1507
rect 1241 1502 1278 1507
rect 1489 1497 1494 1507
rect 1513 1502 1806 1507
rect 1969 1502 2014 1507
rect 2041 1502 2078 1507
rect 2121 1502 2190 1507
rect 425 1492 526 1497
rect 537 1492 878 1497
rect 1201 1492 1270 1497
rect 1345 1492 1470 1497
rect 1489 1492 1542 1497
rect 1657 1492 1774 1497
rect 1849 1492 1958 1497
rect 1953 1487 1958 1492
rect 2017 1492 2046 1497
rect 2017 1487 2022 1492
rect 657 1482 798 1487
rect 1065 1482 1230 1487
rect 1425 1482 1838 1487
rect 1953 1482 2022 1487
rect 2137 1482 2214 1487
rect 2481 1482 2662 1487
rect 1281 1477 1430 1482
rect 425 1472 534 1477
rect 1009 1472 1150 1477
rect 1225 1472 1286 1477
rect 1449 1472 1534 1477
rect 1641 1472 1766 1477
rect 241 1462 326 1467
rect 241 1457 246 1462
rect 217 1452 246 1457
rect 321 1457 326 1462
rect 425 1457 430 1472
rect 321 1452 430 1457
rect 529 1457 534 1472
rect 553 1462 694 1467
rect 801 1462 854 1467
rect 929 1462 1126 1467
rect 1297 1462 1654 1467
rect 1665 1462 1702 1467
rect 1809 1462 1854 1467
rect 1969 1462 2118 1467
rect 2273 1462 2326 1467
rect 2345 1462 2462 1467
rect 689 1457 782 1462
rect 1145 1457 1254 1462
rect 1297 1457 1302 1462
rect 1649 1457 1654 1462
rect 2345 1457 2350 1462
rect 529 1452 670 1457
rect 777 1452 822 1457
rect 993 1452 1150 1457
rect 1249 1452 1302 1457
rect 1433 1452 1526 1457
rect 1649 1452 1742 1457
rect 1849 1452 1942 1457
rect 2097 1452 2262 1457
rect 841 1447 942 1452
rect 2257 1447 2262 1452
rect 2329 1452 2350 1457
rect 2457 1457 2462 1462
rect 2457 1452 2486 1457
rect 2329 1447 2334 1452
rect 129 1442 310 1447
rect 441 1442 470 1447
rect 553 1442 582 1447
rect 745 1442 846 1447
rect 937 1442 1230 1447
rect 1329 1442 1598 1447
rect 1649 1442 1758 1447
rect 1841 1442 1918 1447
rect 2257 1442 2334 1447
rect 2361 1442 2390 1447
rect 465 1437 558 1442
rect 2385 1437 2390 1442
rect 2497 1442 2638 1447
rect 2497 1437 2502 1442
rect 185 1432 214 1437
rect 609 1432 998 1437
rect 1113 1432 1414 1437
rect 2057 1432 2110 1437
rect 2385 1432 2502 1437
rect 609 1427 614 1432
rect 1481 1427 1646 1432
rect 313 1422 614 1427
rect 705 1422 790 1427
rect 897 1422 958 1427
rect 985 1422 1190 1427
rect 1297 1422 1374 1427
rect 1385 1422 1486 1427
rect 1641 1422 1750 1427
rect 1833 1422 1982 1427
rect 2161 1422 2278 1427
rect 2161 1417 2166 1422
rect 569 1412 694 1417
rect 801 1412 878 1417
rect 1001 1412 1062 1417
rect 1121 1412 1630 1417
rect 1769 1412 1798 1417
rect 1985 1412 2166 1417
rect 2273 1417 2278 1422
rect 2273 1412 2302 1417
rect 689 1407 806 1412
rect 1793 1407 1990 1412
rect 353 1402 390 1407
rect 825 1402 1030 1407
rect 1065 1402 1470 1407
rect 1537 1402 1574 1407
rect 2177 1402 2222 1407
rect 1025 1397 1030 1402
rect 265 1392 318 1397
rect 457 1392 566 1397
rect 665 1392 702 1397
rect 873 1392 1014 1397
rect 1025 1392 1302 1397
rect 1393 1392 1590 1397
rect 1609 1392 1870 1397
rect 1897 1392 1998 1397
rect 2233 1392 2470 1397
rect 2641 1392 2758 1397
rect 929 1382 950 1387
rect 1129 1382 1214 1387
rect 1313 1382 1342 1387
rect 1457 1382 1566 1387
rect 1585 1382 1662 1387
rect 1977 1382 2078 1387
rect 361 1377 614 1382
rect 969 1377 1062 1382
rect 1209 1377 1302 1382
rect 1585 1377 1590 1382
rect 2225 1377 2334 1382
rect 185 1372 214 1377
rect 337 1372 366 1377
rect 609 1372 710 1377
rect 729 1372 854 1377
rect 905 1372 974 1377
rect 1057 1372 1086 1377
rect 1297 1372 1366 1377
rect 1377 1372 1590 1377
rect 1601 1372 1726 1377
rect 1753 1372 1878 1377
rect 2201 1372 2230 1377
rect 2329 1372 2358 1377
rect 729 1367 734 1372
rect 137 1362 326 1367
rect 321 1357 326 1362
rect 393 1362 422 1367
rect 473 1362 526 1367
rect 569 1362 734 1367
rect 849 1367 854 1372
rect 849 1362 1030 1367
rect 1049 1362 1078 1367
rect 1121 1362 1230 1367
rect 1449 1362 1630 1367
rect 1793 1362 1822 1367
rect 393 1357 398 1362
rect 1817 1357 1822 1362
rect 1889 1362 2006 1367
rect 2225 1362 2446 1367
rect 1889 1357 1894 1362
rect 2225 1357 2230 1362
rect 321 1352 398 1357
rect 497 1352 582 1357
rect 601 1352 774 1357
rect 793 1352 1158 1357
rect 1153 1347 1158 1352
rect 1241 1352 1374 1357
rect 1417 1352 1486 1357
rect 1601 1352 1694 1357
rect 1817 1352 1894 1357
rect 2105 1352 2230 1357
rect 1241 1347 1246 1352
rect 1481 1347 1606 1352
rect 185 1342 238 1347
rect 465 1342 510 1347
rect 617 1342 646 1347
rect 825 1342 854 1347
rect 505 1337 622 1342
rect 849 1337 854 1342
rect 953 1342 1134 1347
rect 1153 1342 1246 1347
rect 1425 1342 1462 1347
rect 1625 1342 1718 1347
rect 2361 1342 2494 1347
rect 953 1337 958 1342
rect 193 1332 334 1337
rect 481 1327 486 1337
rect 849 1332 958 1337
rect 977 1332 1046 1337
rect 1305 1332 1438 1337
rect 1545 1332 1942 1337
rect 1961 1332 2222 1337
rect 2337 1332 2406 1337
rect 481 1322 830 1327
rect 1153 1322 1286 1327
rect 1505 1322 1750 1327
rect 2521 1322 2678 1327
rect 1153 1317 1158 1322
rect 225 1312 270 1317
rect 353 1312 390 1317
rect 489 1312 518 1317
rect 225 1302 294 1307
rect 513 1297 518 1312
rect 801 1312 950 1317
rect 993 1312 1030 1317
rect 1073 1312 1158 1317
rect 1281 1317 1286 1322
rect 1281 1312 1358 1317
rect 1377 1312 1814 1317
rect 1849 1312 1918 1317
rect 1929 1312 2342 1317
rect 2409 1312 2542 1317
rect 801 1297 806 1312
rect 1137 1302 1214 1307
rect 1425 1302 1646 1307
rect 1881 1302 1998 1307
rect 1641 1297 1886 1302
rect 201 1292 246 1297
rect 513 1292 806 1297
rect 1009 1292 1046 1297
rect 1169 1292 1278 1297
rect 1297 1292 1390 1297
rect 1409 1292 1438 1297
rect 1521 1292 1622 1297
rect 1297 1287 1302 1292
rect 825 1282 998 1287
rect 1057 1282 1158 1287
rect 1169 1282 1302 1287
rect 1385 1287 1390 1292
rect 1385 1282 1470 1287
rect 1641 1282 1750 1287
rect 993 1277 1062 1282
rect 1153 1277 1158 1282
rect 1641 1277 1646 1282
rect 145 1272 286 1277
rect 329 1272 414 1277
rect 1153 1272 1646 1277
rect 1745 1277 1750 1282
rect 1825 1282 2254 1287
rect 2329 1282 2422 1287
rect 1825 1277 1830 1282
rect 1745 1272 1830 1277
rect 2249 1277 2254 1282
rect 2249 1272 2278 1277
rect 2449 1272 2534 1277
rect 329 1267 334 1272
rect 305 1262 334 1267
rect 409 1267 414 1272
rect 1929 1267 1998 1272
rect 2449 1267 2454 1272
rect 409 1262 806 1267
rect 1041 1262 1374 1267
rect 1473 1262 1734 1267
rect 801 1247 806 1262
rect 1729 1257 1734 1262
rect 1841 1262 1934 1267
rect 1993 1262 2270 1267
rect 1841 1257 1846 1262
rect 2265 1257 2270 1262
rect 2361 1262 2454 1267
rect 2529 1267 2534 1272
rect 2529 1262 2558 1267
rect 2361 1257 2366 1262
rect 945 1252 1030 1257
rect 1361 1252 1590 1257
rect 1025 1247 1366 1252
rect 1585 1247 1590 1252
rect 1657 1252 1710 1257
rect 1729 1252 1846 1257
rect 1945 1252 2038 1257
rect 2265 1252 2366 1257
rect 2385 1252 2758 1257
rect 1657 1247 1662 1252
rect 121 1242 398 1247
rect 801 1242 878 1247
rect 1385 1242 1518 1247
rect 1585 1242 1662 1247
rect 873 1237 878 1242
rect 1705 1237 1710 1252
rect 1945 1247 1950 1252
rect 1865 1242 1950 1247
rect 1865 1237 1870 1242
rect 2001 1237 2078 1242
rect 753 1232 790 1237
rect 873 1232 1374 1237
rect 1449 1232 1478 1237
rect 1705 1232 1870 1237
rect 1977 1232 2006 1237
rect 2073 1232 2246 1237
rect 2385 1232 2542 1237
rect 1369 1227 1454 1232
rect 481 1222 518 1227
rect 705 1222 806 1227
rect 1201 1217 1206 1227
rect 1489 1222 1598 1227
rect 1969 1222 2062 1227
rect 2081 1217 2214 1222
rect 233 1212 318 1217
rect 537 1212 686 1217
rect 825 1212 862 1217
rect 913 1212 1030 1217
rect 1057 1212 1102 1217
rect 1201 1212 1398 1217
rect 1889 1212 2086 1217
rect 2209 1212 2286 1217
rect 2321 1212 2430 1217
rect 441 1207 542 1212
rect 681 1207 806 1212
rect 913 1207 918 1212
rect 417 1202 446 1207
rect 801 1202 870 1207
rect 889 1202 918 1207
rect 1025 1207 1030 1212
rect 2425 1207 2430 1212
rect 2553 1212 2630 1217
rect 2553 1207 2558 1212
rect 1025 1202 1054 1207
rect 1169 1202 1190 1207
rect 1697 1202 1870 1207
rect 865 1197 870 1202
rect 1697 1197 1702 1202
rect 377 1192 598 1197
rect 657 1192 854 1197
rect 865 1192 1702 1197
rect 1865 1197 1870 1202
rect 2001 1202 2206 1207
rect 2425 1202 2558 1207
rect 2001 1197 2006 1202
rect 1865 1192 2006 1197
rect 2017 1192 2086 1197
rect 2265 1192 2406 1197
rect 849 1187 854 1192
rect 2105 1187 2230 1192
rect 313 1182 486 1187
rect 529 1182 574 1187
rect 849 1182 1126 1187
rect 1145 1182 1198 1187
rect 1809 1182 2070 1187
rect 2081 1182 2110 1187
rect 2225 1182 2286 1187
rect 1249 1177 1398 1182
rect 2065 1177 2070 1182
rect 641 1172 1254 1177
rect 1393 1172 1534 1177
rect 1713 1172 2022 1177
rect 2065 1172 2214 1177
rect 321 1162 422 1167
rect 473 1162 550 1167
rect 1137 1162 1382 1167
rect 1553 1162 1694 1167
rect 1777 1162 1918 1167
rect 2009 1162 2310 1167
rect 569 1157 1118 1162
rect 1409 1157 1558 1162
rect 1689 1157 1694 1162
rect 241 1152 574 1157
rect 1113 1152 1254 1157
rect 1393 1152 1414 1157
rect 1689 1152 1942 1157
rect 2017 1152 2046 1157
rect 2121 1152 2678 1157
rect 1249 1147 1398 1152
rect 2017 1147 2022 1152
rect 81 1142 142 1147
rect 305 1142 382 1147
rect 409 1142 470 1147
rect 545 1142 606 1147
rect 617 1142 1230 1147
rect 1417 1142 1526 1147
rect 1769 1142 2022 1147
rect 2033 1142 2350 1147
rect 185 1132 222 1137
rect 265 1132 302 1137
rect 801 1132 830 1137
rect 825 1127 830 1132
rect 953 1132 1006 1137
rect 953 1127 958 1132
rect 481 1122 678 1127
rect 825 1122 958 1127
rect 1001 1117 1006 1132
rect 1137 1132 1190 1137
rect 1137 1117 1142 1132
rect 1001 1112 1142 1117
rect 1185 1117 1190 1132
rect 1329 1132 1382 1137
rect 1329 1117 1334 1132
rect 1185 1112 1334 1117
rect 1377 1117 1382 1132
rect 1585 1132 1638 1137
rect 1585 1117 1590 1132
rect 1377 1112 1590 1117
rect 1633 1117 1638 1132
rect 1801 1132 1886 1137
rect 2185 1132 2230 1137
rect 2361 1132 2446 1137
rect 2593 1132 2654 1137
rect 1801 1117 1806 1132
rect 2225 1127 2366 1132
rect 1937 1122 2206 1127
rect 1633 1112 1806 1117
rect 1825 1112 1934 1117
rect 1961 1112 1990 1117
rect 1985 1097 1990 1112
rect 2313 1112 2462 1117
rect 2313 1107 2318 1112
rect 2217 1102 2318 1107
rect 2217 1097 2222 1102
rect 273 1092 310 1097
rect 1457 1092 1518 1097
rect 1985 1092 2222 1097
rect 889 1052 950 1057
rect 457 1032 518 1037
rect 1553 1032 2006 1037
rect 2297 1032 2358 1037
rect 1553 1027 1558 1032
rect 441 1022 550 1027
rect 1529 1022 1558 1027
rect 2001 1027 2006 1032
rect 2001 1022 2030 1027
rect 2065 1022 2126 1027
rect 2145 1017 2150 1027
rect 89 1012 190 1017
rect 337 1012 454 1017
rect 617 1012 758 1017
rect 1153 1012 1430 1017
rect 1577 1012 1966 1017
rect 2145 1012 2214 1017
rect 433 1002 574 1007
rect 617 997 622 1012
rect 753 997 758 1012
rect 1577 1007 1582 1012
rect 1489 1002 1582 1007
rect 1961 1007 1966 1012
rect 1961 1002 1990 1007
rect 265 992 310 997
rect 449 992 622 997
rect 665 992 734 997
rect 753 992 782 997
rect 921 992 1062 997
rect 1097 992 1278 997
rect 665 987 670 992
rect 633 982 670 987
rect 729 987 734 992
rect 1097 987 1102 992
rect 729 982 1102 987
rect 1273 987 1278 992
rect 1489 987 1494 1002
rect 1505 992 1710 997
rect 1729 992 1966 997
rect 1273 982 1494 987
rect 1657 982 1726 987
rect 2465 982 2526 987
rect 681 972 830 977
rect 1113 972 1262 977
rect 1681 972 1782 977
rect 825 967 1014 972
rect 1113 967 1118 972
rect 241 962 294 967
rect 473 962 502 967
rect 537 962 806 967
rect 1009 962 1118 967
rect 1625 962 1814 967
rect 1849 962 1974 967
rect 2001 962 2374 967
rect 369 952 758 957
rect 897 952 990 957
rect 1137 952 1166 957
rect 1249 952 1286 957
rect 1489 952 1734 957
rect 1753 952 1862 957
rect 2281 952 2318 957
rect 2545 952 2622 957
rect 753 947 758 952
rect 121 942 230 947
rect 441 942 734 947
rect 753 942 790 947
rect 881 942 910 947
rect 905 937 910 942
rect 969 942 1094 947
rect 1137 942 1206 947
rect 1433 942 1470 947
rect 969 937 974 942
rect 465 927 470 937
rect 481 932 566 937
rect 593 932 622 937
rect 785 932 814 937
rect 905 932 974 937
rect 1089 937 1094 942
rect 1089 932 1206 937
rect 617 927 622 932
rect 681 927 790 932
rect 1201 927 1206 932
rect 1297 932 1422 937
rect 1297 927 1302 932
rect 337 922 446 927
rect 465 922 486 927
rect 617 922 686 927
rect 1201 922 1302 927
rect 1417 927 1422 932
rect 1489 927 1494 952
rect 1569 942 1678 947
rect 1713 942 1806 947
rect 1945 942 2046 947
rect 2233 942 2262 947
rect 2305 942 2438 947
rect 2513 942 2582 947
rect 1833 937 1918 942
rect 1809 932 1838 937
rect 1913 932 1982 937
rect 1689 927 1766 932
rect 2257 927 2262 942
rect 2289 932 2390 937
rect 2473 932 2526 937
rect 1417 922 1494 927
rect 1561 922 1694 927
rect 1761 922 1902 927
rect 2257 922 2302 927
rect 2561 922 2678 927
rect 2321 917 2454 922
rect 113 912 198 917
rect 433 912 550 917
rect 705 912 846 917
rect 1145 912 1174 917
rect 1705 912 1734 917
rect 1841 912 1870 917
rect 2137 912 2326 917
rect 2449 912 2478 917
rect 1729 907 1846 912
rect 2561 907 2566 922
rect 2593 912 2758 917
rect 369 902 398 907
rect 1049 902 1182 907
rect 2265 902 2310 907
rect 2353 902 2566 907
rect 2577 902 2606 907
rect 2625 902 2662 907
rect 465 892 630 897
rect 729 892 926 897
rect 1657 892 1694 897
rect 1689 887 1694 892
rect 1801 892 1830 897
rect 2089 892 2134 897
rect 1801 887 1806 892
rect 673 882 726 887
rect 1225 882 1334 887
rect 1353 882 1486 887
rect 1689 882 1806 887
rect 2129 887 2134 892
rect 2249 892 2294 897
rect 2313 892 2638 897
rect 2249 887 2254 892
rect 2129 882 2254 887
rect 1225 877 1230 882
rect 1201 872 1230 877
rect 1329 877 1334 882
rect 2289 877 2294 892
rect 2417 882 2470 887
rect 2417 877 2422 882
rect 1329 872 1390 877
rect 2289 872 2422 877
rect 2465 877 2470 882
rect 2545 882 2574 887
rect 2545 877 2550 882
rect 2465 872 2550 877
rect 809 862 918 867
rect 1097 862 1262 867
rect 1913 862 2110 867
rect 809 857 814 862
rect 609 852 814 857
rect 913 857 918 862
rect 1281 857 1390 862
rect 913 852 942 857
rect 1073 852 1286 857
rect 1385 852 1446 857
rect 1913 847 1918 862
rect 2105 847 2110 862
rect 2129 852 2174 857
rect 2193 852 2430 857
rect 2193 847 2198 852
rect 1121 842 1374 847
rect 1889 842 1918 847
rect 2001 842 2086 847
rect 2105 842 2198 847
rect 2425 847 2430 852
rect 2425 842 2478 847
rect 993 837 1086 842
rect 2001 837 2006 842
rect 281 832 334 837
rect 825 832 998 837
rect 1081 832 1318 837
rect 1513 832 2006 837
rect 2081 837 2086 842
rect 2081 832 2414 837
rect 2601 832 2646 837
rect 393 822 510 827
rect 1009 822 1070 827
rect 1209 822 1582 827
rect 2017 822 2190 827
rect 1089 817 1190 822
rect 2417 817 2422 827
rect 2537 822 2614 827
rect 2625 822 2758 827
rect 465 812 542 817
rect 721 812 782 817
rect 1041 812 1094 817
rect 1185 812 1358 817
rect 1497 812 1526 817
rect 2049 812 2286 817
rect 2345 812 2422 817
rect 2433 812 2550 817
rect 1041 807 1046 812
rect 1353 807 1502 812
rect 129 802 254 807
rect 361 802 390 807
rect 553 802 838 807
rect 945 802 1046 807
rect 1057 802 1334 807
rect 1521 802 1566 807
rect 2057 802 2134 807
rect 2273 802 2310 807
rect 2641 802 2710 807
rect 385 797 390 802
rect 473 797 558 802
rect 1057 797 1062 802
rect 1521 797 1526 802
rect 385 792 478 797
rect 689 792 750 797
rect 745 787 750 792
rect 849 792 902 797
rect 913 792 1062 797
rect 1145 792 1214 797
rect 1337 792 1526 797
rect 1665 792 1734 797
rect 1753 792 1894 797
rect 2001 792 2118 797
rect 2161 792 2206 797
rect 2449 792 2502 797
rect 2617 792 2702 797
rect 849 787 854 792
rect 1753 787 1758 792
rect 497 782 558 787
rect 681 782 726 787
rect 745 782 854 787
rect 1137 782 1198 787
rect 1545 782 1758 787
rect 1889 787 1894 792
rect 1889 782 1918 787
rect 2121 782 2214 787
rect 2233 782 2382 787
rect 2233 777 2238 782
rect 1009 772 1254 777
rect 1273 772 1630 777
rect 1705 772 1846 777
rect 2009 772 2238 777
rect 2377 777 2382 782
rect 2377 772 2678 777
rect 593 762 870 767
rect 881 762 1078 767
rect 1337 762 1454 767
rect 1529 762 1694 767
rect 1857 762 1998 767
rect 2113 762 2366 767
rect 1689 757 1862 762
rect 1993 757 2118 762
rect 289 752 406 757
rect 1081 752 1318 757
rect 1481 752 1654 757
rect 2137 752 2182 757
rect 193 742 302 747
rect 321 742 430 747
rect 521 742 814 747
rect 889 742 966 747
rect 1001 742 1142 747
rect 1177 742 1422 747
rect 1569 742 1598 747
rect 1641 742 1758 747
rect 1793 742 1942 747
rect 2049 742 2134 747
rect 2257 742 2310 747
rect 2425 742 2542 747
rect 2625 742 2702 747
rect 273 737 278 742
rect 1793 737 1798 742
rect 273 732 342 737
rect 857 732 990 737
rect 1257 732 1622 737
rect 1633 732 1798 737
rect 1809 732 1862 737
rect 2001 732 2246 737
rect 721 727 838 732
rect 1793 727 1798 732
rect 577 722 654 727
rect 697 722 726 727
rect 833 722 950 727
rect 1009 722 1094 727
rect 1385 722 1646 727
rect 1793 722 1822 727
rect 1921 722 1990 727
rect 2257 722 2462 727
rect 1009 717 1014 722
rect 305 712 342 717
rect 473 712 550 717
rect 569 712 1014 717
rect 1089 717 1094 722
rect 1241 717 1350 722
rect 1985 717 2262 722
rect 1089 712 1118 717
rect 1217 712 1246 717
rect 1345 712 1374 717
rect 1433 712 1462 717
rect 1545 712 1910 717
rect 2529 712 2582 717
rect 2617 712 2758 717
rect 473 707 478 712
rect 449 702 478 707
rect 545 707 550 712
rect 2577 707 2582 712
rect 545 702 590 707
rect 633 702 726 707
rect 777 702 982 707
rect 993 702 1078 707
rect 1281 702 1350 707
rect 1361 702 1478 707
rect 1553 702 1630 707
rect 1657 702 1830 707
rect 1881 702 2086 707
rect 2201 702 2366 707
rect 2577 702 2630 707
rect 1097 697 1238 702
rect 1553 697 1558 702
rect 2201 697 2206 702
rect 209 692 478 697
rect 665 692 822 697
rect 833 692 1102 697
rect 1233 692 1558 697
rect 1577 692 1758 697
rect 817 687 822 692
rect 1753 687 1758 692
rect 1849 692 1926 697
rect 1937 692 2206 697
rect 2361 697 2366 702
rect 2361 692 2470 697
rect 1849 687 1854 692
rect 377 682 406 687
rect 401 677 406 682
rect 505 682 598 687
rect 705 682 750 687
rect 817 682 1222 687
rect 1289 682 1550 687
rect 1641 682 1670 687
rect 1753 682 1854 687
rect 1921 687 1926 692
rect 1921 682 2350 687
rect 505 677 510 682
rect 1545 677 1646 682
rect 401 672 510 677
rect 825 672 1382 677
rect 1425 672 1526 677
rect 1873 672 1902 677
rect 2225 672 2542 677
rect 1897 667 2230 672
rect 737 662 814 667
rect 1113 662 1486 667
rect 1585 662 1782 667
rect 809 657 1118 662
rect 1585 657 1590 662
rect 529 652 710 657
rect 1137 652 1166 657
rect 1297 652 1430 657
rect 1505 652 1590 657
rect 1777 657 1782 662
rect 2249 657 2342 662
rect 1777 652 2254 657
rect 2337 652 2446 657
rect 1161 647 1302 652
rect 409 642 510 647
rect 409 637 414 642
rect 385 632 414 637
rect 505 637 510 642
rect 729 642 878 647
rect 729 637 734 642
rect 505 632 678 637
rect 697 632 734 637
rect 873 637 878 642
rect 921 642 1014 647
rect 1033 642 1126 647
rect 1321 642 1414 647
rect 921 637 926 642
rect 873 632 926 637
rect 1009 637 1014 642
rect 1009 632 1286 637
rect 1361 632 1494 637
rect 673 627 678 632
rect 129 622 182 627
rect 265 622 318 627
rect 673 622 806 627
rect 817 622 894 627
rect 913 622 1006 627
rect 1233 622 1302 627
rect 1393 622 1470 627
rect 801 617 806 622
rect 1025 617 1214 622
rect 1505 617 1510 652
rect 1601 642 1766 647
rect 2097 642 2174 647
rect 2097 637 2102 642
rect 1609 632 1678 637
rect 1961 632 2102 637
rect 1529 622 1838 627
rect 2033 622 2134 627
rect 2225 622 2230 652
rect 2289 642 2326 647
rect 2433 642 2470 647
rect 2249 632 2310 637
rect 2313 622 2438 627
rect 2449 622 2526 627
rect 2585 622 2686 627
rect 345 612 414 617
rect 465 612 614 617
rect 681 612 782 617
rect 801 612 1030 617
rect 1209 612 1510 617
rect 1841 612 1870 617
rect 2081 612 2142 617
rect 1697 607 1822 612
rect 617 602 678 607
rect 673 597 678 602
rect 777 602 1158 607
rect 1217 602 1246 607
rect 1441 602 1630 607
rect 1673 602 1702 607
rect 1817 602 1990 607
rect 2121 602 2198 607
rect 2337 602 2382 607
rect 2673 602 2734 607
rect 777 597 782 602
rect 81 592 238 597
rect 393 592 510 597
rect 625 592 654 597
rect 673 592 782 597
rect 817 592 854 597
rect 977 592 1006 597
rect 649 577 654 592
rect 817 577 822 592
rect 1001 587 1006 592
rect 1073 592 1102 597
rect 1161 592 1190 597
rect 1073 587 1078 592
rect 841 582 910 587
rect 1001 582 1078 587
rect 1217 582 1222 602
rect 1241 597 1446 602
rect 1985 597 1990 602
rect 1465 592 1502 597
rect 1545 592 1862 597
rect 1889 592 1974 597
rect 1985 592 2062 597
rect 2137 592 2174 597
rect 2305 592 2390 597
rect 2465 592 2694 597
rect 2721 592 2758 597
rect 2465 587 2470 592
rect 1329 582 1574 587
rect 1665 582 1742 587
rect 1809 582 1910 587
rect 2353 582 2470 587
rect 1569 577 1670 582
rect 169 572 390 577
rect 649 572 822 577
rect 1177 572 1366 577
rect 1441 572 1550 577
rect 1705 572 1806 577
rect 1889 572 2158 577
rect 2233 572 2342 577
rect 2337 567 2342 572
rect 2481 572 2558 577
rect 2481 567 2486 572
rect 369 562 462 567
rect 1457 562 1718 567
rect 1729 562 1926 567
rect 2337 562 2486 567
rect 1713 557 1718 562
rect 2153 557 2238 562
rect 1409 552 1582 557
rect 1713 552 1750 557
rect 2097 552 2158 557
rect 2233 552 2278 557
rect 129 542 238 547
rect 1145 542 1398 547
rect 1393 537 1398 542
rect 1465 542 1542 547
rect 1729 542 1918 547
rect 1945 542 2014 547
rect 2169 542 2206 547
rect 2241 542 2542 547
rect 2681 542 2758 547
rect 1465 537 1470 542
rect 1729 537 1734 542
rect 1945 537 1950 542
rect 969 532 1030 537
rect 1393 532 1470 537
rect 1489 532 1734 537
rect 1753 532 1950 537
rect 2009 537 2014 542
rect 2009 532 2110 537
rect 361 522 430 527
rect 513 522 742 527
rect 761 522 982 527
rect 1873 522 1998 527
rect 737 517 742 522
rect 1633 517 1750 522
rect 737 512 822 517
rect 817 507 822 512
rect 921 512 974 517
rect 921 507 926 512
rect 817 502 926 507
rect 969 507 974 512
rect 1041 512 1358 517
rect 1537 512 1638 517
rect 1745 512 1774 517
rect 1817 512 1966 517
rect 1041 507 1046 512
rect 1961 507 1966 512
rect 2121 512 2190 517
rect 2121 507 2126 512
rect 969 502 1046 507
rect 1649 502 1718 507
rect 1961 502 2126 507
rect 1713 497 1718 502
rect 1561 492 1694 497
rect 1713 492 1910 497
rect 665 482 798 487
rect 753 472 854 477
rect 1177 472 1646 477
rect 1657 472 1782 477
rect 81 462 350 467
rect 1521 462 1550 467
rect 1705 462 1734 467
rect 1793 462 1878 467
rect 1545 457 1654 462
rect 1729 457 1798 462
rect 1649 452 1710 457
rect 1313 442 1446 447
rect 1465 442 1838 447
rect 2025 442 2126 447
rect 185 432 222 437
rect 969 432 1046 437
rect 1313 427 1318 442
rect 393 422 446 427
rect 681 422 774 427
rect 849 422 894 427
rect 969 422 1070 427
rect 1193 422 1270 427
rect 1289 422 1318 427
rect 1441 427 1446 442
rect 1713 432 1742 437
rect 1873 432 1902 437
rect 1977 432 2006 437
rect 2137 432 2222 437
rect 1737 427 1878 432
rect 2001 427 2142 432
rect 1441 422 1542 427
rect 1561 422 1694 427
rect 2305 422 2414 427
rect 2425 422 2550 427
rect 1193 417 1198 422
rect 241 412 686 417
rect 921 412 1198 417
rect 1265 417 1270 422
rect 1561 417 1566 422
rect 1265 412 1326 417
rect 1337 412 1430 417
rect 1425 407 1430 412
rect 1497 412 1566 417
rect 1689 417 1694 422
rect 1689 412 1774 417
rect 1793 412 1926 417
rect 1945 412 2118 417
rect 2569 412 2670 417
rect 1497 407 1502 412
rect 1793 407 1798 412
rect 1033 402 1166 407
rect 1425 402 1502 407
rect 1521 402 1798 407
rect 1921 407 1926 412
rect 1921 402 1990 407
rect 2281 402 2318 407
rect 801 392 902 397
rect 1209 392 1382 397
rect 1713 392 2214 397
rect 2545 392 2654 397
rect 1049 382 1070 387
rect 1153 382 1206 387
rect 1473 382 1574 387
rect 1593 382 1846 387
rect 1865 382 1982 387
rect 2169 382 2198 387
rect 2433 382 2494 387
rect 1473 377 1478 382
rect 409 372 478 377
rect 409 367 414 372
rect 385 362 414 367
rect 473 367 478 372
rect 921 372 1030 377
rect 921 367 926 372
rect 473 362 926 367
rect 1025 367 1030 372
rect 1225 372 1318 377
rect 1449 372 1478 377
rect 1569 377 1574 382
rect 1977 377 2174 382
rect 1569 372 1718 377
rect 1761 372 1862 377
rect 2321 372 2582 377
rect 1225 367 1230 372
rect 1025 362 1230 367
rect 1313 367 1318 372
rect 2577 367 2582 372
rect 1313 362 1582 367
rect 1777 362 2142 367
rect 1577 357 1782 362
rect 2137 357 2142 362
rect 2209 362 2366 367
rect 2577 362 2678 367
rect 2209 357 2214 362
rect 409 352 446 357
rect 1241 352 1302 357
rect 441 347 446 352
rect 1145 347 1246 352
rect 1297 347 1302 352
rect 1425 352 1454 357
rect 1497 352 1558 357
rect 1801 352 1830 357
rect 1425 347 1430 352
rect 1825 347 1830 352
rect 1913 352 1942 357
rect 2137 352 2214 357
rect 1913 347 1918 352
rect 297 342 422 347
rect 441 342 1150 347
rect 1297 342 1430 347
rect 1537 342 1638 347
rect 1737 342 1806 347
rect 1825 342 1918 347
rect 2033 342 2118 347
rect 1193 332 1278 337
rect 1193 327 1198 332
rect 689 322 918 327
rect 1169 322 1198 327
rect 1273 327 1278 332
rect 1489 332 1526 337
rect 1681 332 1758 337
rect 1977 332 2022 337
rect 2521 332 2758 337
rect 1489 327 1494 332
rect 1273 322 1494 327
rect 1505 322 1614 327
rect 1921 322 2038 327
rect 689 317 694 322
rect 2033 317 2038 322
rect 369 312 694 317
rect 857 312 1342 317
rect 1913 312 2014 317
rect 2033 312 2214 317
rect 2425 312 2582 317
rect 1153 292 1262 297
rect 2433 292 2470 297
rect 2617 272 2678 277
rect 2185 252 2294 257
rect 2185 247 2190 252
rect 2137 242 2190 247
rect 2289 247 2294 252
rect 2449 252 2526 257
rect 2553 252 2630 257
rect 2449 247 2454 252
rect 2289 242 2454 247
rect 2521 247 2526 252
rect 2521 242 2550 247
rect 2009 232 2086 237
rect 2529 232 2582 237
rect 2009 227 2014 232
rect 209 222 446 227
rect 1585 222 1694 227
rect 1985 222 2014 227
rect 2081 227 2086 232
rect 2081 222 2110 227
rect 2201 222 2278 227
rect 2465 222 2518 227
rect 1193 212 1310 217
rect 1193 207 1198 212
rect 585 202 1046 207
rect 1081 202 1198 207
rect 1305 207 1310 212
rect 1433 212 1542 217
rect 1433 207 1438 212
rect 1305 202 1438 207
rect 1537 207 1542 212
rect 1585 207 1590 222
rect 1537 202 1590 207
rect 1689 207 1694 222
rect 2705 217 2710 227
rect 1737 212 1830 217
rect 2281 212 2710 217
rect 1737 207 1742 212
rect 1689 202 1742 207
rect 1825 207 1830 212
rect 1825 202 2118 207
rect 2241 202 2294 207
rect 705 192 710 202
rect 1041 197 1046 202
rect 2241 197 2246 202
rect 1041 192 1142 197
rect 1137 187 1142 192
rect 1217 192 1302 197
rect 1217 187 1222 192
rect 905 182 934 187
rect 929 177 934 182
rect 1001 182 1030 187
rect 1137 182 1222 187
rect 1297 187 1302 192
rect 1409 192 1646 197
rect 2129 192 2246 197
rect 2257 192 2342 197
rect 1409 187 1414 192
rect 1297 182 1414 187
rect 1641 187 1646 192
rect 1905 187 2062 192
rect 2129 187 2134 192
rect 1641 182 1910 187
rect 2057 182 2134 187
rect 2281 182 2574 187
rect 1001 177 1006 182
rect 313 172 366 177
rect 529 172 598 177
rect 929 172 1006 177
rect 1929 172 2038 177
rect 2265 172 2326 177
rect 193 162 246 167
rect 625 162 718 167
rect 1257 162 1350 167
rect 1409 162 1478 167
rect 1521 162 1622 167
rect 433 152 486 157
rect 1649 152 1822 157
rect 2521 152 2598 157
rect 145 142 182 147
rect 177 137 182 142
rect 241 142 422 147
rect 241 137 246 142
rect 177 132 246 137
rect 417 137 422 142
rect 489 142 662 147
rect 489 137 494 142
rect 417 132 494 137
rect 657 137 662 142
rect 721 142 1142 147
rect 1153 142 1542 147
rect 1593 142 1678 147
rect 1913 142 2182 147
rect 2249 142 2494 147
rect 2513 142 2542 147
rect 2657 142 2758 147
rect 721 137 726 142
rect 657 132 726 137
rect 1137 137 1142 142
rect 1913 137 1918 142
rect 1137 132 1166 137
rect 1513 132 1590 137
rect 1161 127 1262 132
rect 1257 117 1262 127
rect 1513 117 1518 132
rect 1585 127 1590 132
rect 1689 132 1918 137
rect 2177 137 2182 142
rect 2177 132 2238 137
rect 1689 127 1694 132
rect 2233 127 2238 132
rect 2361 127 2502 132
rect 1537 122 1566 127
rect 1585 122 1694 127
rect 1929 122 2054 127
rect 745 112 862 117
rect 1097 112 1126 117
rect 1121 107 1126 112
rect 1209 112 1238 117
rect 1257 112 1518 117
rect 1209 107 1214 112
rect 1121 102 1214 107
rect 1561 107 1566 122
rect 1929 107 1934 122
rect 2049 117 2054 122
rect 2113 122 2158 127
rect 2233 122 2366 127
rect 2497 122 2678 127
rect 2113 117 2118 122
rect 2049 112 2118 117
rect 2137 112 2166 117
rect 1561 102 1934 107
rect 2161 107 2166 112
rect 2385 112 2414 117
rect 2385 107 2390 112
rect 2161 102 2390 107
use AND2X2  AND2X2_0
timestamp 1711307567
transform 1 0 2256 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1711307567
transform 1 0 1672 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1711307567
transform 1 0 1448 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1711307567
transform 1 0 936 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1711307567
transform 1 0 936 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1711307567
transform 1 0 480 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1711307567
transform 1 0 1544 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1711307567
transform 1 0 968 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1711307567
transform 1 0 2640 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1711307567
transform 1 0 1840 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1711307567
transform 1 0 1368 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1711307567
transform 1 0 1680 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1711307567
transform 1 0 696 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1711307567
transform 1 0 2160 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1711307567
transform 1 0 768 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1711307567
transform 1 0 520 0 1 2370
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1711307567
transform 1 0 1544 0 1 2370
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1711307567
transform 1 0 1472 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1711307567
transform 1 0 1768 0 1 2370
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1711307567
transform 1 0 648 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_20
timestamp 1711307567
transform 1 0 1224 0 1 2370
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1711307567
transform 1 0 1400 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1711307567
transform 1 0 2296 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_23
timestamp 1711307567
transform 1 0 1328 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1711307567
transform 1 0 480 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_25
timestamp 1711307567
transform 1 0 1720 0 -1 2370
box -8 -3 40 105
use AND2X2  AND2X2_26
timestamp 1711307567
transform 1 0 1824 0 -1 2370
box -8 -3 40 105
use AND2X2  AND2X2_27
timestamp 1711307567
transform 1 0 1976 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_28
timestamp 1711307567
transform 1 0 2520 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_29
timestamp 1711307567
transform 1 0 2464 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_30
timestamp 1711307567
transform 1 0 2456 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_31
timestamp 1711307567
transform 1 0 2264 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_32
timestamp 1711307567
transform 1 0 768 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_33
timestamp 1711307567
transform 1 0 1040 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_34
timestamp 1711307567
transform 1 0 1880 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_35
timestamp 1711307567
transform 1 0 1320 0 1 2370
box -8 -3 40 105
use AND2X2  AND2X2_36
timestamp 1711307567
transform 1 0 296 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_37
timestamp 1711307567
transform 1 0 456 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_38
timestamp 1711307567
transform 1 0 504 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_39
timestamp 1711307567
transform 1 0 416 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_40
timestamp 1711307567
transform 1 0 1040 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_41
timestamp 1711307567
transform 1 0 872 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_42
timestamp 1711307567
transform 1 0 1568 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_43
timestamp 1711307567
transform 1 0 1632 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_44
timestamp 1711307567
transform 1 0 2272 0 -1 2170
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1711307567
transform 1 0 2552 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1711307567
transform 1 0 1696 0 1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1711307567
transform 1 0 808 0 1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1711307567
transform 1 0 528 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1711307567
transform 1 0 880 0 1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1711307567
transform 1 0 784 0 -1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1711307567
transform 1 0 384 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1711307567
transform 1 0 272 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1711307567
transform 1 0 240 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1711307567
transform 1 0 368 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1711307567
transform 1 0 464 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1711307567
transform 1 0 400 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1711307567
transform 1 0 600 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1711307567
transform 1 0 368 0 -1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1711307567
transform 1 0 440 0 1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1711307567
transform 1 0 448 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1711307567
transform 1 0 688 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1711307567
transform 1 0 832 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1711307567
transform 1 0 768 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1711307567
transform 1 0 816 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1711307567
transform 1 0 1016 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1711307567
transform 1 0 1016 0 -1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1711307567
transform 1 0 896 0 -1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1711307567
transform 1 0 1104 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1711307567
transform 1 0 1200 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1711307567
transform 1 0 1240 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1711307567
transform 1 0 1160 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_27
timestamp 1711307567
transform 1 0 1168 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_28
timestamp 1711307567
transform 1 0 1256 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_29
timestamp 1711307567
transform 1 0 1520 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_30
timestamp 1711307567
transform 1 0 1512 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_31
timestamp 1711307567
transform 1 0 1712 0 -1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_32
timestamp 1711307567
transform 1 0 1720 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_33
timestamp 1711307567
transform 1 0 1624 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_34
timestamp 1711307567
transform 1 0 1768 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_35
timestamp 1711307567
transform 1 0 1896 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_36
timestamp 1711307567
transform 1 0 2088 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_37
timestamp 1711307567
transform 1 0 1912 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_38
timestamp 1711307567
transform 1 0 1968 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_39
timestamp 1711307567
transform 1 0 2592 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_40
timestamp 1711307567
transform 1 0 1536 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_41
timestamp 1711307567
transform 1 0 1304 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_42
timestamp 1711307567
transform 1 0 2232 0 -1 570
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1711307567
transform 1 0 464 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1711307567
transform 1 0 1384 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1711307567
transform 1 0 1272 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1711307567
transform 1 0 552 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1711307567
transform 1 0 1392 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1711307567
transform 1 0 1024 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1711307567
transform 1 0 336 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1711307567
transform 1 0 1584 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1711307567
transform 1 0 1856 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1711307567
transform 1 0 1248 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1711307567
transform 1 0 832 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1711307567
transform 1 0 1200 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1711307567
transform 1 0 376 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1711307567
transform 1 0 1544 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1711307567
transform 1 0 1448 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1711307567
transform 1 0 1320 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1711307567
transform 1 0 568 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1711307567
transform 1 0 1320 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1711307567
transform 1 0 360 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1711307567
transform 1 0 1544 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1711307567
transform 1 0 2560 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1711307567
transform 1 0 2648 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1711307567
transform 1 0 2696 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1711307567
transform 1 0 2632 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1711307567
transform 1 0 2592 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1711307567
transform 1 0 2688 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1711307567
transform 1 0 2120 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1711307567
transform 1 0 2040 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1711307567
transform 1 0 2128 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1711307567
transform 1 0 1968 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1711307567
transform 1 0 2088 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1711307567
transform 1 0 1960 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1711307567
transform 1 0 2160 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1711307567
transform 1 0 1920 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1711307567
transform 1 0 2032 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1711307567
transform 1 0 1896 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1711307567
transform 1 0 1888 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1711307567
transform 1 0 1752 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1711307567
transform 1 0 1816 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1711307567
transform 1 0 1672 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1711307567
transform 1 0 1288 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1711307567
transform 1 0 1216 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1711307567
transform 1 0 1160 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1711307567
transform 1 0 1152 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1711307567
transform 1 0 896 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1711307567
transform 1 0 752 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1711307567
transform 1 0 840 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1711307567
transform 1 0 824 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1711307567
transform 1 0 688 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1711307567
transform 1 0 640 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1711307567
transform 1 0 568 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1711307567
transform 1 0 600 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1711307567
transform 1 0 432 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1711307567
transform 1 0 440 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1711307567
transform 1 0 528 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_55
timestamp 1711307567
transform 1 0 528 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1711307567
transform 1 0 2552 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_57
timestamp 1711307567
transform 1 0 2520 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_58
timestamp 1711307567
transform 1 0 2512 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_59
timestamp 1711307567
transform 1 0 2392 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_60
timestamp 1711307567
transform 1 0 1712 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_61
timestamp 1711307567
transform 1 0 1704 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_62
timestamp 1711307567
transform 1 0 1848 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_63
timestamp 1711307567
transform 1 0 2384 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_64
timestamp 1711307567
transform 1 0 2512 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_65
timestamp 1711307567
transform 1 0 2384 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_66
timestamp 1711307567
transform 1 0 1928 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_67
timestamp 1711307567
transform 1 0 288 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_68
timestamp 1711307567
transform 1 0 208 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_69
timestamp 1711307567
transform 1 0 2184 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_70
timestamp 1711307567
transform 1 0 128 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_71
timestamp 1711307567
transform 1 0 208 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1711307567
transform 1 0 304 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_73
timestamp 1711307567
transform 1 0 184 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_74
timestamp 1711307567
transform 1 0 376 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_75
timestamp 1711307567
transform 1 0 456 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_76
timestamp 1711307567
transform 1 0 672 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_77
timestamp 1711307567
transform 1 0 656 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_78
timestamp 1711307567
transform 1 0 584 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_79
timestamp 1711307567
transform 1 0 968 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_80
timestamp 1711307567
transform 1 0 2312 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_81
timestamp 1711307567
transform 1 0 856 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_82
timestamp 1711307567
transform 1 0 1040 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_83
timestamp 1711307567
transform 1 0 1128 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_84
timestamp 1711307567
transform 1 0 1232 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_85
timestamp 1711307567
transform 1 0 1424 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_86
timestamp 1711307567
transform 1 0 1240 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_87
timestamp 1711307567
transform 1 0 1368 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_88
timestamp 1711307567
transform 1 0 1600 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_89
timestamp 1711307567
transform 1 0 1584 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_90
timestamp 1711307567
transform 1 0 1760 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_91
timestamp 1711307567
transform 1 0 2080 0 -1 1170
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1711307567
transform 1 0 1496 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1711307567
transform 1 0 1472 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1711307567
transform 1 0 2736 0 1 570
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1711307567
transform 1 0 2728 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1711307567
transform 1 0 2032 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1711307567
transform 1 0 1544 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1711307567
transform 1 0 1456 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1711307567
transform 1 0 1552 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1711307567
transform 1 0 1416 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1711307567
transform 1 0 1456 0 1 1170
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1711307567
transform 1 0 1904 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1711307567
transform 1 0 2216 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1711307567
transform 1 0 1656 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1711307567
transform 1 0 1928 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1711307567
transform 1 0 1992 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1711307567
transform 1 0 2016 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1711307567
transform 1 0 1848 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1711307567
transform 1 0 1824 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1711307567
transform 1 0 1976 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1711307567
transform 1 0 2200 0 1 170
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1711307567
transform 1 0 2192 0 1 370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1711307567
transform 1 0 2648 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1711307567
transform 1 0 2472 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1711307567
transform 1 0 2464 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1711307567
transform 1 0 2392 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1711307567
transform 1 0 2352 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1711307567
transform 1 0 2448 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1711307567
transform 1 0 2232 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1711307567
transform 1 0 2472 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1711307567
transform 1 0 2200 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1711307567
transform 1 0 2296 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1711307567
transform 1 0 2360 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1711307567
transform 1 0 2424 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1711307567
transform 1 0 2440 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1711307567
transform 1 0 2192 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1711307567
transform 1 0 2280 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1711307567
transform 1 0 2360 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1711307567
transform 1 0 2312 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1711307567
transform 1 0 2464 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1711307567
transform 1 0 2528 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1711307567
transform 1 0 2408 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1711307567
transform 1 0 96 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1711307567
transform 1 0 80 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1711307567
transform 1 0 80 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1711307567
transform 1 0 208 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1711307567
transform 1 0 296 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1711307567
transform 1 0 120 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1711307567
transform 1 0 368 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1711307567
transform 1 0 472 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1711307567
transform 1 0 752 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1711307567
transform 1 0 664 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1711307567
transform 1 0 584 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1711307567
transform 1 0 928 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1711307567
transform 1 0 840 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1711307567
transform 1 0 1008 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1711307567
transform 1 0 1048 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1711307567
transform 1 0 1216 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1711307567
transform 1 0 1344 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1711307567
transform 1 0 1144 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1711307567
transform 1 0 1304 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1711307567
transform 1 0 1600 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1711307567
transform 1 0 1496 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1711307567
transform 1 0 1704 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1711307567
transform 1 0 1696 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1711307567
transform 1 0 1608 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1711307567
transform 1 0 1808 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1711307567
transform 1 0 2336 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1711307567
transform 1 0 2432 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1711307567
transform 1 0 2184 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1711307567
transform 1 0 1976 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1711307567
transform 1 0 2096 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1711307567
transform 1 0 2240 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1711307567
transform 1 0 2072 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1711307567
transform 1 0 1424 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1711307567
transform 1 0 336 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1711307567
transform 1 0 72 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1711307567
transform 1 0 80 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1711307567
transform 1 0 80 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1711307567
transform 1 0 256 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1711307567
transform 1 0 136 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1711307567
transform 1 0 504 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1711307567
transform 1 0 376 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1711307567
transform 1 0 800 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1711307567
transform 1 0 768 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1711307567
transform 1 0 624 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1711307567
transform 1 0 920 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1711307567
transform 1 0 920 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1711307567
transform 1 0 1144 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1711307567
transform 1 0 1280 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1711307567
transform 1 0 1256 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1711307567
transform 1 0 1464 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1711307567
transform 1 0 1360 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1711307567
transform 1 0 1528 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1711307567
transform 1 0 1624 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1711307567
transform 1 0 1944 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1711307567
transform 1 0 2104 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1711307567
transform 1 0 2016 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1711307567
transform 1 0 2016 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1711307567
transform 1 0 1968 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1711307567
transform 1 0 2664 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1711307567
transform 1 0 2664 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1711307567
transform 1 0 2488 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1711307567
transform 1 0 2344 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1711307567
transform 1 0 2592 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1711307567
transform 1 0 2664 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1711307567
transform 1 0 2344 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1711307567
transform 1 0 2320 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1711307567
transform 1 0 224 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1711307567
transform 1 0 72 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1711307567
transform 1 0 72 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1711307567
transform 1 0 128 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1711307567
transform 1 0 232 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1711307567
transform 1 0 128 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1711307567
transform 1 0 504 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1711307567
transform 1 0 432 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1711307567
transform 1 0 624 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1711307567
transform 1 0 672 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1711307567
transform 1 0 552 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1711307567
transform 1 0 936 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1711307567
transform 1 0 848 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1711307567
transform 1 0 1048 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1711307567
transform 1 0 1048 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1711307567
transform 1 0 1184 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1711307567
transform 1 0 1640 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1711307567
transform 1 0 1304 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1711307567
transform 1 0 1384 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1711307567
transform 1 0 1768 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1711307567
transform 1 0 1736 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1711307567
transform 1 0 1768 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1711307567
transform 1 0 1808 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1711307567
transform 1 0 1776 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1711307567
transform 1 0 1888 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1711307567
transform 1 0 2664 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1711307567
transform 1 0 2600 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1711307567
transform 1 0 2448 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1711307567
transform 1 0 2112 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1711307567
transform 1 0 2352 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1711307567
transform 1 0 2544 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1711307567
transform 1 0 2192 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1711307567
transform 1 0 2312 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1711307567
transform 1 0 2448 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1711307567
transform 1 0 2560 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1711307567
transform 1 0 2256 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1711307567
transform 1 0 2656 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1711307567
transform 1 0 2664 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1711307567
transform 1 0 2664 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1711307567
transform 1 0 2608 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1711307567
transform 1 0 2144 0 -1 170
box -8 -3 104 105
use FILL  FILL_0
timestamp 1711307567
transform 1 0 2752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1
timestamp 1711307567
transform 1 0 2664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_2
timestamp 1711307567
transform 1 0 2600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_3
timestamp 1711307567
transform 1 0 2552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4
timestamp 1711307567
transform 1 0 2544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5
timestamp 1711307567
transform 1 0 2488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_6
timestamp 1711307567
transform 1 0 2192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_7
timestamp 1711307567
transform 1 0 2096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1711307567
transform 1 0 2032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_9
timestamp 1711307567
transform 1 0 2000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_10
timestamp 1711307567
transform 1 0 1944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_11
timestamp 1711307567
transform 1 0 1936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_12
timestamp 1711307567
transform 1 0 1896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_13
timestamp 1711307567
transform 1 0 1888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_14
timestamp 1711307567
transform 1 0 1816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_15
timestamp 1711307567
transform 1 0 1808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_16
timestamp 1711307567
transform 1 0 1800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_17
timestamp 1711307567
transform 1 0 1744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_18
timestamp 1711307567
transform 1 0 1704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_19
timestamp 1711307567
transform 1 0 1696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_20
timestamp 1711307567
transform 1 0 1688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_21
timestamp 1711307567
transform 1 0 1640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_22
timestamp 1711307567
transform 1 0 1632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_23
timestamp 1711307567
transform 1 0 1576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_24
timestamp 1711307567
transform 1 0 1544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_25
timestamp 1711307567
transform 1 0 1536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_26
timestamp 1711307567
transform 1 0 1464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_27
timestamp 1711307567
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_28
timestamp 1711307567
transform 1 0 1392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_29
timestamp 1711307567
transform 1 0 1384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_30
timestamp 1711307567
transform 1 0 1376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_31
timestamp 1711307567
transform 1 0 1304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_32
timestamp 1711307567
transform 1 0 1296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_33
timestamp 1711307567
transform 1 0 1288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_34
timestamp 1711307567
transform 1 0 1240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_35
timestamp 1711307567
transform 1 0 1192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_36
timestamp 1711307567
transform 1 0 1184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_37
timestamp 1711307567
transform 1 0 1176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_38
timestamp 1711307567
transform 1 0 1168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_39
timestamp 1711307567
transform 1 0 1160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_40
timestamp 1711307567
transform 1 0 1088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_41
timestamp 1711307567
transform 1 0 1080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_42
timestamp 1711307567
transform 1 0 1072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_43
timestamp 1711307567
transform 1 0 1016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_44
timestamp 1711307567
transform 1 0 1008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_45
timestamp 1711307567
transform 1 0 1000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_46
timestamp 1711307567
transform 1 0 944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_47
timestamp 1711307567
transform 1 0 936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_48
timestamp 1711307567
transform 1 0 928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_49
timestamp 1711307567
transform 1 0 888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_50
timestamp 1711307567
transform 1 0 848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_51
timestamp 1711307567
transform 1 0 840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_52
timestamp 1711307567
transform 1 0 832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_53
timestamp 1711307567
transform 1 0 768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_54
timestamp 1711307567
transform 1 0 760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_55
timestamp 1711307567
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_56
timestamp 1711307567
transform 1 0 680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_57
timestamp 1711307567
transform 1 0 672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_58
timestamp 1711307567
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_59
timestamp 1711307567
transform 1 0 608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_60
timestamp 1711307567
transform 1 0 600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_61
timestamp 1711307567
transform 1 0 536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_62
timestamp 1711307567
transform 1 0 496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_63
timestamp 1711307567
transform 1 0 440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_64
timestamp 1711307567
transform 1 0 432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_65
timestamp 1711307567
transform 1 0 424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_66
timestamp 1711307567
transform 1 0 360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_67
timestamp 1711307567
transform 1 0 352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_68
timestamp 1711307567
transform 1 0 344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_69
timestamp 1711307567
transform 1 0 288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_70
timestamp 1711307567
transform 1 0 280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_71
timestamp 1711307567
transform 1 0 272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_72
timestamp 1711307567
transform 1 0 264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_73
timestamp 1711307567
transform 1 0 256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_74
timestamp 1711307567
transform 1 0 248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_75
timestamp 1711307567
transform 1 0 240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_76
timestamp 1711307567
transform 1 0 232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_77
timestamp 1711307567
transform 1 0 224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_78
timestamp 1711307567
transform 1 0 216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_79
timestamp 1711307567
transform 1 0 208 0 -1 2570
box -8 -3 16 105
use FILL  FILL_80
timestamp 1711307567
transform 1 0 200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_81
timestamp 1711307567
transform 1 0 192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_82
timestamp 1711307567
transform 1 0 184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_83
timestamp 1711307567
transform 1 0 176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_84
timestamp 1711307567
transform 1 0 168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_85
timestamp 1711307567
transform 1 0 160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_86
timestamp 1711307567
transform 1 0 152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_87
timestamp 1711307567
transform 1 0 144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_88
timestamp 1711307567
transform 1 0 136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_89
timestamp 1711307567
transform 1 0 128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_90
timestamp 1711307567
transform 1 0 120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_91
timestamp 1711307567
transform 1 0 112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_92
timestamp 1711307567
transform 1 0 104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_93
timestamp 1711307567
transform 1 0 96 0 -1 2570
box -8 -3 16 105
use FILL  FILL_94
timestamp 1711307567
transform 1 0 88 0 -1 2570
box -8 -3 16 105
use FILL  FILL_95
timestamp 1711307567
transform 1 0 80 0 -1 2570
box -8 -3 16 105
use FILL  FILL_96
timestamp 1711307567
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_97
timestamp 1711307567
transform 1 0 2696 0 1 2370
box -8 -3 16 105
use FILL  FILL_98
timestamp 1711307567
transform 1 0 2688 0 1 2370
box -8 -3 16 105
use FILL  FILL_99
timestamp 1711307567
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use FILL  FILL_100
timestamp 1711307567
transform 1 0 2632 0 1 2370
box -8 -3 16 105
use FILL  FILL_101
timestamp 1711307567
transform 1 0 2544 0 1 2370
box -8 -3 16 105
use FILL  FILL_102
timestamp 1711307567
transform 1 0 2536 0 1 2370
box -8 -3 16 105
use FILL  FILL_103
timestamp 1711307567
transform 1 0 2528 0 1 2370
box -8 -3 16 105
use FILL  FILL_104
timestamp 1711307567
transform 1 0 2472 0 1 2370
box -8 -3 16 105
use FILL  FILL_105
timestamp 1711307567
transform 1 0 2464 0 1 2370
box -8 -3 16 105
use FILL  FILL_106
timestamp 1711307567
transform 1 0 2456 0 1 2370
box -8 -3 16 105
use FILL  FILL_107
timestamp 1711307567
transform 1 0 2448 0 1 2370
box -8 -3 16 105
use FILL  FILL_108
timestamp 1711307567
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use FILL  FILL_109
timestamp 1711307567
transform 1 0 2336 0 1 2370
box -8 -3 16 105
use FILL  FILL_110
timestamp 1711307567
transform 1 0 2328 0 1 2370
box -8 -3 16 105
use FILL  FILL_111
timestamp 1711307567
transform 1 0 2320 0 1 2370
box -8 -3 16 105
use FILL  FILL_112
timestamp 1711307567
transform 1 0 2312 0 1 2370
box -8 -3 16 105
use FILL  FILL_113
timestamp 1711307567
transform 1 0 2304 0 1 2370
box -8 -3 16 105
use FILL  FILL_114
timestamp 1711307567
transform 1 0 2296 0 1 2370
box -8 -3 16 105
use FILL  FILL_115
timestamp 1711307567
transform 1 0 2288 0 1 2370
box -8 -3 16 105
use FILL  FILL_116
timestamp 1711307567
transform 1 0 2184 0 1 2370
box -8 -3 16 105
use FILL  FILL_117
timestamp 1711307567
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_118
timestamp 1711307567
transform 1 0 2112 0 1 2370
box -8 -3 16 105
use FILL  FILL_119
timestamp 1711307567
transform 1 0 2104 0 1 2370
box -8 -3 16 105
use FILL  FILL_120
timestamp 1711307567
transform 1 0 2096 0 1 2370
box -8 -3 16 105
use FILL  FILL_121
timestamp 1711307567
transform 1 0 2088 0 1 2370
box -8 -3 16 105
use FILL  FILL_122
timestamp 1711307567
transform 1 0 2080 0 1 2370
box -8 -3 16 105
use FILL  FILL_123
timestamp 1711307567
transform 1 0 2072 0 1 2370
box -8 -3 16 105
use FILL  FILL_124
timestamp 1711307567
transform 1 0 2016 0 1 2370
box -8 -3 16 105
use FILL  FILL_125
timestamp 1711307567
transform 1 0 2008 0 1 2370
box -8 -3 16 105
use FILL  FILL_126
timestamp 1711307567
transform 1 0 2000 0 1 2370
box -8 -3 16 105
use FILL  FILL_127
timestamp 1711307567
transform 1 0 1992 0 1 2370
box -8 -3 16 105
use FILL  FILL_128
timestamp 1711307567
transform 1 0 1952 0 1 2370
box -8 -3 16 105
use FILL  FILL_129
timestamp 1711307567
transform 1 0 1912 0 1 2370
box -8 -3 16 105
use FILL  FILL_130
timestamp 1711307567
transform 1 0 1904 0 1 2370
box -8 -3 16 105
use FILL  FILL_131
timestamp 1711307567
transform 1 0 1896 0 1 2370
box -8 -3 16 105
use FILL  FILL_132
timestamp 1711307567
transform 1 0 1888 0 1 2370
box -8 -3 16 105
use FILL  FILL_133
timestamp 1711307567
transform 1 0 1848 0 1 2370
box -8 -3 16 105
use FILL  FILL_134
timestamp 1711307567
transform 1 0 1808 0 1 2370
box -8 -3 16 105
use FILL  FILL_135
timestamp 1711307567
transform 1 0 1800 0 1 2370
box -8 -3 16 105
use FILL  FILL_136
timestamp 1711307567
transform 1 0 1760 0 1 2370
box -8 -3 16 105
use FILL  FILL_137
timestamp 1711307567
transform 1 0 1752 0 1 2370
box -8 -3 16 105
use FILL  FILL_138
timestamp 1711307567
transform 1 0 1744 0 1 2370
box -8 -3 16 105
use FILL  FILL_139
timestamp 1711307567
transform 1 0 1736 0 1 2370
box -8 -3 16 105
use FILL  FILL_140
timestamp 1711307567
transform 1 0 1704 0 1 2370
box -8 -3 16 105
use FILL  FILL_141
timestamp 1711307567
transform 1 0 1696 0 1 2370
box -8 -3 16 105
use FILL  FILL_142
timestamp 1711307567
transform 1 0 1664 0 1 2370
box -8 -3 16 105
use FILL  FILL_143
timestamp 1711307567
transform 1 0 1656 0 1 2370
box -8 -3 16 105
use FILL  FILL_144
timestamp 1711307567
transform 1 0 1648 0 1 2370
box -8 -3 16 105
use FILL  FILL_145
timestamp 1711307567
transform 1 0 1640 0 1 2370
box -8 -3 16 105
use FILL  FILL_146
timestamp 1711307567
transform 1 0 1632 0 1 2370
box -8 -3 16 105
use FILL  FILL_147
timestamp 1711307567
transform 1 0 1592 0 1 2370
box -8 -3 16 105
use FILL  FILL_148
timestamp 1711307567
transform 1 0 1584 0 1 2370
box -8 -3 16 105
use FILL  FILL_149
timestamp 1711307567
transform 1 0 1576 0 1 2370
box -8 -3 16 105
use FILL  FILL_150
timestamp 1711307567
transform 1 0 1536 0 1 2370
box -8 -3 16 105
use FILL  FILL_151
timestamp 1711307567
transform 1 0 1528 0 1 2370
box -8 -3 16 105
use FILL  FILL_152
timestamp 1711307567
transform 1 0 1496 0 1 2370
box -8 -3 16 105
use FILL  FILL_153
timestamp 1711307567
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_154
timestamp 1711307567
transform 1 0 1480 0 1 2370
box -8 -3 16 105
use FILL  FILL_155
timestamp 1711307567
transform 1 0 1472 0 1 2370
box -8 -3 16 105
use FILL  FILL_156
timestamp 1711307567
transform 1 0 1432 0 1 2370
box -8 -3 16 105
use FILL  FILL_157
timestamp 1711307567
transform 1 0 1424 0 1 2370
box -8 -3 16 105
use FILL  FILL_158
timestamp 1711307567
transform 1 0 1416 0 1 2370
box -8 -3 16 105
use FILL  FILL_159
timestamp 1711307567
transform 1 0 1408 0 1 2370
box -8 -3 16 105
use FILL  FILL_160
timestamp 1711307567
transform 1 0 1368 0 1 2370
box -8 -3 16 105
use FILL  FILL_161
timestamp 1711307567
transform 1 0 1360 0 1 2370
box -8 -3 16 105
use FILL  FILL_162
timestamp 1711307567
transform 1 0 1352 0 1 2370
box -8 -3 16 105
use FILL  FILL_163
timestamp 1711307567
transform 1 0 1312 0 1 2370
box -8 -3 16 105
use FILL  FILL_164
timestamp 1711307567
transform 1 0 1304 0 1 2370
box -8 -3 16 105
use FILL  FILL_165
timestamp 1711307567
transform 1 0 1272 0 1 2370
box -8 -3 16 105
use FILL  FILL_166
timestamp 1711307567
transform 1 0 1264 0 1 2370
box -8 -3 16 105
use FILL  FILL_167
timestamp 1711307567
transform 1 0 1256 0 1 2370
box -8 -3 16 105
use FILL  FILL_168
timestamp 1711307567
transform 1 0 1216 0 1 2370
box -8 -3 16 105
use FILL  FILL_169
timestamp 1711307567
transform 1 0 1208 0 1 2370
box -8 -3 16 105
use FILL  FILL_170
timestamp 1711307567
transform 1 0 1200 0 1 2370
box -8 -3 16 105
use FILL  FILL_171
timestamp 1711307567
transform 1 0 1192 0 1 2370
box -8 -3 16 105
use FILL  FILL_172
timestamp 1711307567
transform 1 0 1168 0 1 2370
box -8 -3 16 105
use FILL  FILL_173
timestamp 1711307567
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_174
timestamp 1711307567
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use FILL  FILL_175
timestamp 1711307567
transform 1 0 1120 0 1 2370
box -8 -3 16 105
use FILL  FILL_176
timestamp 1711307567
transform 1 0 1112 0 1 2370
box -8 -3 16 105
use FILL  FILL_177
timestamp 1711307567
transform 1 0 1104 0 1 2370
box -8 -3 16 105
use FILL  FILL_178
timestamp 1711307567
transform 1 0 1096 0 1 2370
box -8 -3 16 105
use FILL  FILL_179
timestamp 1711307567
transform 1 0 1064 0 1 2370
box -8 -3 16 105
use FILL  FILL_180
timestamp 1711307567
transform 1 0 1056 0 1 2370
box -8 -3 16 105
use FILL  FILL_181
timestamp 1711307567
transform 1 0 1048 0 1 2370
box -8 -3 16 105
use FILL  FILL_182
timestamp 1711307567
transform 1 0 1024 0 1 2370
box -8 -3 16 105
use FILL  FILL_183
timestamp 1711307567
transform 1 0 1016 0 1 2370
box -8 -3 16 105
use FILL  FILL_184
timestamp 1711307567
transform 1 0 1008 0 1 2370
box -8 -3 16 105
use FILL  FILL_185
timestamp 1711307567
transform 1 0 1000 0 1 2370
box -8 -3 16 105
use FILL  FILL_186
timestamp 1711307567
transform 1 0 992 0 1 2370
box -8 -3 16 105
use FILL  FILL_187
timestamp 1711307567
transform 1 0 984 0 1 2370
box -8 -3 16 105
use FILL  FILL_188
timestamp 1711307567
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_189
timestamp 1711307567
transform 1 0 936 0 1 2370
box -8 -3 16 105
use FILL  FILL_190
timestamp 1711307567
transform 1 0 928 0 1 2370
box -8 -3 16 105
use FILL  FILL_191
timestamp 1711307567
transform 1 0 920 0 1 2370
box -8 -3 16 105
use FILL  FILL_192
timestamp 1711307567
transform 1 0 912 0 1 2370
box -8 -3 16 105
use FILL  FILL_193
timestamp 1711307567
transform 1 0 904 0 1 2370
box -8 -3 16 105
use FILL  FILL_194
timestamp 1711307567
transform 1 0 896 0 1 2370
box -8 -3 16 105
use FILL  FILL_195
timestamp 1711307567
transform 1 0 888 0 1 2370
box -8 -3 16 105
use FILL  FILL_196
timestamp 1711307567
transform 1 0 880 0 1 2370
box -8 -3 16 105
use FILL  FILL_197
timestamp 1711307567
transform 1 0 872 0 1 2370
box -8 -3 16 105
use FILL  FILL_198
timestamp 1711307567
transform 1 0 832 0 1 2370
box -8 -3 16 105
use FILL  FILL_199
timestamp 1711307567
transform 1 0 824 0 1 2370
box -8 -3 16 105
use FILL  FILL_200
timestamp 1711307567
transform 1 0 816 0 1 2370
box -8 -3 16 105
use FILL  FILL_201
timestamp 1711307567
transform 1 0 808 0 1 2370
box -8 -3 16 105
use FILL  FILL_202
timestamp 1711307567
transform 1 0 800 0 1 2370
box -8 -3 16 105
use FILL  FILL_203
timestamp 1711307567
transform 1 0 792 0 1 2370
box -8 -3 16 105
use FILL  FILL_204
timestamp 1711307567
transform 1 0 784 0 1 2370
box -8 -3 16 105
use FILL  FILL_205
timestamp 1711307567
transform 1 0 736 0 1 2370
box -8 -3 16 105
use FILL  FILL_206
timestamp 1711307567
transform 1 0 728 0 1 2370
box -8 -3 16 105
use FILL  FILL_207
timestamp 1711307567
transform 1 0 720 0 1 2370
box -8 -3 16 105
use FILL  FILL_208
timestamp 1711307567
transform 1 0 712 0 1 2370
box -8 -3 16 105
use FILL  FILL_209
timestamp 1711307567
transform 1 0 688 0 1 2370
box -8 -3 16 105
use FILL  FILL_210
timestamp 1711307567
transform 1 0 680 0 1 2370
box -8 -3 16 105
use FILL  FILL_211
timestamp 1711307567
transform 1 0 672 0 1 2370
box -8 -3 16 105
use FILL  FILL_212
timestamp 1711307567
transform 1 0 632 0 1 2370
box -8 -3 16 105
use FILL  FILL_213
timestamp 1711307567
transform 1 0 624 0 1 2370
box -8 -3 16 105
use FILL  FILL_214
timestamp 1711307567
transform 1 0 616 0 1 2370
box -8 -3 16 105
use FILL  FILL_215
timestamp 1711307567
transform 1 0 608 0 1 2370
box -8 -3 16 105
use FILL  FILL_216
timestamp 1711307567
transform 1 0 568 0 1 2370
box -8 -3 16 105
use FILL  FILL_217
timestamp 1711307567
transform 1 0 560 0 1 2370
box -8 -3 16 105
use FILL  FILL_218
timestamp 1711307567
transform 1 0 552 0 1 2370
box -8 -3 16 105
use FILL  FILL_219
timestamp 1711307567
transform 1 0 512 0 1 2370
box -8 -3 16 105
use FILL  FILL_220
timestamp 1711307567
transform 1 0 504 0 1 2370
box -8 -3 16 105
use FILL  FILL_221
timestamp 1711307567
transform 1 0 472 0 1 2370
box -8 -3 16 105
use FILL  FILL_222
timestamp 1711307567
transform 1 0 448 0 1 2370
box -8 -3 16 105
use FILL  FILL_223
timestamp 1711307567
transform 1 0 440 0 1 2370
box -8 -3 16 105
use FILL  FILL_224
timestamp 1711307567
transform 1 0 432 0 1 2370
box -8 -3 16 105
use FILL  FILL_225
timestamp 1711307567
transform 1 0 424 0 1 2370
box -8 -3 16 105
use FILL  FILL_226
timestamp 1711307567
transform 1 0 376 0 1 2370
box -8 -3 16 105
use FILL  FILL_227
timestamp 1711307567
transform 1 0 368 0 1 2370
box -8 -3 16 105
use FILL  FILL_228
timestamp 1711307567
transform 1 0 360 0 1 2370
box -8 -3 16 105
use FILL  FILL_229
timestamp 1711307567
transform 1 0 352 0 1 2370
box -8 -3 16 105
use FILL  FILL_230
timestamp 1711307567
transform 1 0 320 0 1 2370
box -8 -3 16 105
use FILL  FILL_231
timestamp 1711307567
transform 1 0 288 0 1 2370
box -8 -3 16 105
use FILL  FILL_232
timestamp 1711307567
transform 1 0 280 0 1 2370
box -8 -3 16 105
use FILL  FILL_233
timestamp 1711307567
transform 1 0 248 0 1 2370
box -8 -3 16 105
use FILL  FILL_234
timestamp 1711307567
transform 1 0 240 0 1 2370
box -8 -3 16 105
use FILL  FILL_235
timestamp 1711307567
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_236
timestamp 1711307567
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_237
timestamp 1711307567
transform 1 0 152 0 1 2370
box -8 -3 16 105
use FILL  FILL_238
timestamp 1711307567
transform 1 0 144 0 1 2370
box -8 -3 16 105
use FILL  FILL_239
timestamp 1711307567
transform 1 0 120 0 1 2370
box -8 -3 16 105
use FILL  FILL_240
timestamp 1711307567
transform 1 0 112 0 1 2370
box -8 -3 16 105
use FILL  FILL_241
timestamp 1711307567
transform 1 0 104 0 1 2370
box -8 -3 16 105
use FILL  FILL_242
timestamp 1711307567
transform 1 0 96 0 1 2370
box -8 -3 16 105
use FILL  FILL_243
timestamp 1711307567
transform 1 0 88 0 1 2370
box -8 -3 16 105
use FILL  FILL_244
timestamp 1711307567
transform 1 0 80 0 1 2370
box -8 -3 16 105
use FILL  FILL_245
timestamp 1711307567
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_246
timestamp 1711307567
transform 1 0 2752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_247
timestamp 1711307567
transform 1 0 2744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_248
timestamp 1711307567
transform 1 0 2736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_249
timestamp 1711307567
transform 1 0 2688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_250
timestamp 1711307567
transform 1 0 2680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_251
timestamp 1711307567
transform 1 0 2672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_252
timestamp 1711307567
transform 1 0 2632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_253
timestamp 1711307567
transform 1 0 2624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_254
timestamp 1711307567
transform 1 0 2592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_255
timestamp 1711307567
transform 1 0 2552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_256
timestamp 1711307567
transform 1 0 2544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_257
timestamp 1711307567
transform 1 0 2440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_258
timestamp 1711307567
transform 1 0 2432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_259
timestamp 1711307567
transform 1 0 2424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_260
timestamp 1711307567
transform 1 0 2392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_261
timestamp 1711307567
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_262
timestamp 1711307567
transform 1 0 2376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_263
timestamp 1711307567
transform 1 0 2272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_264
timestamp 1711307567
transform 1 0 2264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_265
timestamp 1711307567
transform 1 0 2256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_266
timestamp 1711307567
transform 1 0 2248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_267
timestamp 1711307567
transform 1 0 2240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_268
timestamp 1711307567
transform 1 0 2232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_269
timestamp 1711307567
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_270
timestamp 1711307567
transform 1 0 2192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_271
timestamp 1711307567
transform 1 0 2160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_272
timestamp 1711307567
transform 1 0 2152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_273
timestamp 1711307567
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_274
timestamp 1711307567
transform 1 0 2136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_275
timestamp 1711307567
transform 1 0 2096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_276
timestamp 1711307567
transform 1 0 2088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_277
timestamp 1711307567
transform 1 0 2080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_278
timestamp 1711307567
transform 1 0 2056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_279
timestamp 1711307567
transform 1 0 2048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_280
timestamp 1711307567
transform 1 0 2040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_281
timestamp 1711307567
transform 1 0 2032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_282
timestamp 1711307567
transform 1 0 1992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_283
timestamp 1711307567
transform 1 0 1984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_284
timestamp 1711307567
transform 1 0 1976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_285
timestamp 1711307567
transform 1 0 1968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_286
timestamp 1711307567
transform 1 0 1960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_287
timestamp 1711307567
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_288
timestamp 1711307567
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_289
timestamp 1711307567
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_290
timestamp 1711307567
transform 1 0 1888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_291
timestamp 1711307567
transform 1 0 1880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_292
timestamp 1711307567
transform 1 0 1872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_293
timestamp 1711307567
transform 1 0 1816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_294
timestamp 1711307567
transform 1 0 1808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_295
timestamp 1711307567
transform 1 0 1800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_296
timestamp 1711307567
transform 1 0 1760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_297
timestamp 1711307567
transform 1 0 1752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_298
timestamp 1711307567
transform 1 0 1712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_299
timestamp 1711307567
transform 1 0 1704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_300
timestamp 1711307567
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_301
timestamp 1711307567
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_302
timestamp 1711307567
transform 1 0 1680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_303
timestamp 1711307567
transform 1 0 1632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_304
timestamp 1711307567
transform 1 0 1624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_305
timestamp 1711307567
transform 1 0 1616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_306
timestamp 1711307567
transform 1 0 1608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_307
timestamp 1711307567
transform 1 0 1584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_308
timestamp 1711307567
transform 1 0 1552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_309
timestamp 1711307567
transform 1 0 1544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_310
timestamp 1711307567
transform 1 0 1536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_311
timestamp 1711307567
transform 1 0 1528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_312
timestamp 1711307567
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_313
timestamp 1711307567
transform 1 0 1472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_314
timestamp 1711307567
transform 1 0 1464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_315
timestamp 1711307567
transform 1 0 1456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_316
timestamp 1711307567
transform 1 0 1448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_317
timestamp 1711307567
transform 1 0 1400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_318
timestamp 1711307567
transform 1 0 1392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_319
timestamp 1711307567
transform 1 0 1384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_320
timestamp 1711307567
transform 1 0 1376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_321
timestamp 1711307567
transform 1 0 1368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_322
timestamp 1711307567
transform 1 0 1320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_323
timestamp 1711307567
transform 1 0 1312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_324
timestamp 1711307567
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_325
timestamp 1711307567
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_326
timestamp 1711307567
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_327
timestamp 1711307567
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_328
timestamp 1711307567
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_329
timestamp 1711307567
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_330
timestamp 1711307567
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_331
timestamp 1711307567
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_332
timestamp 1711307567
transform 1 0 1168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_333
timestamp 1711307567
transform 1 0 1160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_334
timestamp 1711307567
transform 1 0 1152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_335
timestamp 1711307567
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_336
timestamp 1711307567
transform 1 0 1104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_337
timestamp 1711307567
transform 1 0 1096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_338
timestamp 1711307567
transform 1 0 1088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_339
timestamp 1711307567
transform 1 0 1080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_340
timestamp 1711307567
transform 1 0 1072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_341
timestamp 1711307567
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_342
timestamp 1711307567
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_343
timestamp 1711307567
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_344
timestamp 1711307567
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_345
timestamp 1711307567
transform 1 0 992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_346
timestamp 1711307567
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_347
timestamp 1711307567
transform 1 0 944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_348
timestamp 1711307567
transform 1 0 936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_349
timestamp 1711307567
transform 1 0 928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_350
timestamp 1711307567
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_351
timestamp 1711307567
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_352
timestamp 1711307567
transform 1 0 872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_353
timestamp 1711307567
transform 1 0 864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_354
timestamp 1711307567
transform 1 0 832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_355
timestamp 1711307567
transform 1 0 824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_356
timestamp 1711307567
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_357
timestamp 1711307567
transform 1 0 776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_358
timestamp 1711307567
transform 1 0 768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_359
timestamp 1711307567
transform 1 0 760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_360
timestamp 1711307567
transform 1 0 752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_361
timestamp 1711307567
transform 1 0 744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_362
timestamp 1711307567
transform 1 0 696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_363
timestamp 1711307567
transform 1 0 688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_364
timestamp 1711307567
transform 1 0 680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_365
timestamp 1711307567
transform 1 0 672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_366
timestamp 1711307567
transform 1 0 640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_367
timestamp 1711307567
transform 1 0 632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_368
timestamp 1711307567
transform 1 0 624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_369
timestamp 1711307567
transform 1 0 616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_370
timestamp 1711307567
transform 1 0 608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_371
timestamp 1711307567
transform 1 0 576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_372
timestamp 1711307567
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_373
timestamp 1711307567
transform 1 0 536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_374
timestamp 1711307567
transform 1 0 528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_375
timestamp 1711307567
transform 1 0 520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_376
timestamp 1711307567
transform 1 0 512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_377
timestamp 1711307567
transform 1 0 504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_378
timestamp 1711307567
transform 1 0 456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_379
timestamp 1711307567
transform 1 0 448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_380
timestamp 1711307567
transform 1 0 440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_381
timestamp 1711307567
transform 1 0 432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_382
timestamp 1711307567
transform 1 0 424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_383
timestamp 1711307567
transform 1 0 416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_384
timestamp 1711307567
transform 1 0 376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_385
timestamp 1711307567
transform 1 0 368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_386
timestamp 1711307567
transform 1 0 360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_387
timestamp 1711307567
transform 1 0 336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_388
timestamp 1711307567
transform 1 0 328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_389
timestamp 1711307567
transform 1 0 320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_390
timestamp 1711307567
transform 1 0 312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_391
timestamp 1711307567
transform 1 0 280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_392
timestamp 1711307567
transform 1 0 272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_393
timestamp 1711307567
transform 1 0 264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_394
timestamp 1711307567
transform 1 0 232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_395
timestamp 1711307567
transform 1 0 224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_396
timestamp 1711307567
transform 1 0 216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_397
timestamp 1711307567
transform 1 0 208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_398
timestamp 1711307567
transform 1 0 200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_399
timestamp 1711307567
transform 1 0 192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_400
timestamp 1711307567
transform 1 0 184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_401
timestamp 1711307567
transform 1 0 176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_402
timestamp 1711307567
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_403
timestamp 1711307567
transform 1 0 2672 0 1 2170
box -8 -3 16 105
use FILL  FILL_404
timestamp 1711307567
transform 1 0 2624 0 1 2170
box -8 -3 16 105
use FILL  FILL_405
timestamp 1711307567
transform 1 0 2616 0 1 2170
box -8 -3 16 105
use FILL  FILL_406
timestamp 1711307567
transform 1 0 2464 0 1 2170
box -8 -3 16 105
use FILL  FILL_407
timestamp 1711307567
transform 1 0 2456 0 1 2170
box -8 -3 16 105
use FILL  FILL_408
timestamp 1711307567
transform 1 0 2352 0 1 2170
box -8 -3 16 105
use FILL  FILL_409
timestamp 1711307567
transform 1 0 2344 0 1 2170
box -8 -3 16 105
use FILL  FILL_410
timestamp 1711307567
transform 1 0 2336 0 1 2170
box -8 -3 16 105
use FILL  FILL_411
timestamp 1711307567
transform 1 0 2328 0 1 2170
box -8 -3 16 105
use FILL  FILL_412
timestamp 1711307567
transform 1 0 2224 0 1 2170
box -8 -3 16 105
use FILL  FILL_413
timestamp 1711307567
transform 1 0 2216 0 1 2170
box -8 -3 16 105
use FILL  FILL_414
timestamp 1711307567
transform 1 0 2208 0 1 2170
box -8 -3 16 105
use FILL  FILL_415
timestamp 1711307567
transform 1 0 2200 0 1 2170
box -8 -3 16 105
use FILL  FILL_416
timestamp 1711307567
transform 1 0 2144 0 1 2170
box -8 -3 16 105
use FILL  FILL_417
timestamp 1711307567
transform 1 0 2136 0 1 2170
box -8 -3 16 105
use FILL  FILL_418
timestamp 1711307567
transform 1 0 2128 0 1 2170
box -8 -3 16 105
use FILL  FILL_419
timestamp 1711307567
transform 1 0 2096 0 1 2170
box -8 -3 16 105
use FILL  FILL_420
timestamp 1711307567
transform 1 0 2088 0 1 2170
box -8 -3 16 105
use FILL  FILL_421
timestamp 1711307567
transform 1 0 2040 0 1 2170
box -8 -3 16 105
use FILL  FILL_422
timestamp 1711307567
transform 1 0 2032 0 1 2170
box -8 -3 16 105
use FILL  FILL_423
timestamp 1711307567
transform 1 0 2024 0 1 2170
box -8 -3 16 105
use FILL  FILL_424
timestamp 1711307567
transform 1 0 2016 0 1 2170
box -8 -3 16 105
use FILL  FILL_425
timestamp 1711307567
transform 1 0 1960 0 1 2170
box -8 -3 16 105
use FILL  FILL_426
timestamp 1711307567
transform 1 0 1952 0 1 2170
box -8 -3 16 105
use FILL  FILL_427
timestamp 1711307567
transform 1 0 1944 0 1 2170
box -8 -3 16 105
use FILL  FILL_428
timestamp 1711307567
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use FILL  FILL_429
timestamp 1711307567
transform 1 0 1888 0 1 2170
box -8 -3 16 105
use FILL  FILL_430
timestamp 1711307567
transform 1 0 1880 0 1 2170
box -8 -3 16 105
use FILL  FILL_431
timestamp 1711307567
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_432
timestamp 1711307567
transform 1 0 1832 0 1 2170
box -8 -3 16 105
use FILL  FILL_433
timestamp 1711307567
transform 1 0 1792 0 1 2170
box -8 -3 16 105
use FILL  FILL_434
timestamp 1711307567
transform 1 0 1784 0 1 2170
box -8 -3 16 105
use FILL  FILL_435
timestamp 1711307567
transform 1 0 1776 0 1 2170
box -8 -3 16 105
use FILL  FILL_436
timestamp 1711307567
transform 1 0 1736 0 1 2170
box -8 -3 16 105
use FILL  FILL_437
timestamp 1711307567
transform 1 0 1728 0 1 2170
box -8 -3 16 105
use FILL  FILL_438
timestamp 1711307567
transform 1 0 1688 0 1 2170
box -8 -3 16 105
use FILL  FILL_439
timestamp 1711307567
transform 1 0 1680 0 1 2170
box -8 -3 16 105
use FILL  FILL_440
timestamp 1711307567
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use FILL  FILL_441
timestamp 1711307567
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use FILL  FILL_442
timestamp 1711307567
transform 1 0 1616 0 1 2170
box -8 -3 16 105
use FILL  FILL_443
timestamp 1711307567
transform 1 0 1608 0 1 2170
box -8 -3 16 105
use FILL  FILL_444
timestamp 1711307567
transform 1 0 1600 0 1 2170
box -8 -3 16 105
use FILL  FILL_445
timestamp 1711307567
transform 1 0 1592 0 1 2170
box -8 -3 16 105
use FILL  FILL_446
timestamp 1711307567
transform 1 0 1584 0 1 2170
box -8 -3 16 105
use FILL  FILL_447
timestamp 1711307567
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_448
timestamp 1711307567
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use FILL  FILL_449
timestamp 1711307567
transform 1 0 1520 0 1 2170
box -8 -3 16 105
use FILL  FILL_450
timestamp 1711307567
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_451
timestamp 1711307567
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_452
timestamp 1711307567
transform 1 0 1472 0 1 2170
box -8 -3 16 105
use FILL  FILL_453
timestamp 1711307567
transform 1 0 1432 0 1 2170
box -8 -3 16 105
use FILL  FILL_454
timestamp 1711307567
transform 1 0 1424 0 1 2170
box -8 -3 16 105
use FILL  FILL_455
timestamp 1711307567
transform 1 0 1416 0 1 2170
box -8 -3 16 105
use FILL  FILL_456
timestamp 1711307567
transform 1 0 1408 0 1 2170
box -8 -3 16 105
use FILL  FILL_457
timestamp 1711307567
transform 1 0 1360 0 1 2170
box -8 -3 16 105
use FILL  FILL_458
timestamp 1711307567
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_459
timestamp 1711307567
transform 1 0 1344 0 1 2170
box -8 -3 16 105
use FILL  FILL_460
timestamp 1711307567
transform 1 0 1336 0 1 2170
box -8 -3 16 105
use FILL  FILL_461
timestamp 1711307567
transform 1 0 1328 0 1 2170
box -8 -3 16 105
use FILL  FILL_462
timestamp 1711307567
transform 1 0 1280 0 1 2170
box -8 -3 16 105
use FILL  FILL_463
timestamp 1711307567
transform 1 0 1272 0 1 2170
box -8 -3 16 105
use FILL  FILL_464
timestamp 1711307567
transform 1 0 1264 0 1 2170
box -8 -3 16 105
use FILL  FILL_465
timestamp 1711307567
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use FILL  FILL_466
timestamp 1711307567
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use FILL  FILL_467
timestamp 1711307567
transform 1 0 1240 0 1 2170
box -8 -3 16 105
use FILL  FILL_468
timestamp 1711307567
transform 1 0 1192 0 1 2170
box -8 -3 16 105
use FILL  FILL_469
timestamp 1711307567
transform 1 0 1184 0 1 2170
box -8 -3 16 105
use FILL  FILL_470
timestamp 1711307567
transform 1 0 1176 0 1 2170
box -8 -3 16 105
use FILL  FILL_471
timestamp 1711307567
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_472
timestamp 1711307567
transform 1 0 1160 0 1 2170
box -8 -3 16 105
use FILL  FILL_473
timestamp 1711307567
transform 1 0 1128 0 1 2170
box -8 -3 16 105
use FILL  FILL_474
timestamp 1711307567
transform 1 0 1120 0 1 2170
box -8 -3 16 105
use FILL  FILL_475
timestamp 1711307567
transform 1 0 1112 0 1 2170
box -8 -3 16 105
use FILL  FILL_476
timestamp 1711307567
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_477
timestamp 1711307567
transform 1 0 1072 0 1 2170
box -8 -3 16 105
use FILL  FILL_478
timestamp 1711307567
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_479
timestamp 1711307567
transform 1 0 1056 0 1 2170
box -8 -3 16 105
use FILL  FILL_480
timestamp 1711307567
transform 1 0 1024 0 1 2170
box -8 -3 16 105
use FILL  FILL_481
timestamp 1711307567
transform 1 0 1016 0 1 2170
box -8 -3 16 105
use FILL  FILL_482
timestamp 1711307567
transform 1 0 1008 0 1 2170
box -8 -3 16 105
use FILL  FILL_483
timestamp 1711307567
transform 1 0 1000 0 1 2170
box -8 -3 16 105
use FILL  FILL_484
timestamp 1711307567
transform 1 0 992 0 1 2170
box -8 -3 16 105
use FILL  FILL_485
timestamp 1711307567
transform 1 0 944 0 1 2170
box -8 -3 16 105
use FILL  FILL_486
timestamp 1711307567
transform 1 0 936 0 1 2170
box -8 -3 16 105
use FILL  FILL_487
timestamp 1711307567
transform 1 0 928 0 1 2170
box -8 -3 16 105
use FILL  FILL_488
timestamp 1711307567
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_489
timestamp 1711307567
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_490
timestamp 1711307567
transform 1 0 872 0 1 2170
box -8 -3 16 105
use FILL  FILL_491
timestamp 1711307567
transform 1 0 864 0 1 2170
box -8 -3 16 105
use FILL  FILL_492
timestamp 1711307567
transform 1 0 856 0 1 2170
box -8 -3 16 105
use FILL  FILL_493
timestamp 1711307567
transform 1 0 848 0 1 2170
box -8 -3 16 105
use FILL  FILL_494
timestamp 1711307567
transform 1 0 840 0 1 2170
box -8 -3 16 105
use FILL  FILL_495
timestamp 1711307567
transform 1 0 800 0 1 2170
box -8 -3 16 105
use FILL  FILL_496
timestamp 1711307567
transform 1 0 792 0 1 2170
box -8 -3 16 105
use FILL  FILL_497
timestamp 1711307567
transform 1 0 784 0 1 2170
box -8 -3 16 105
use FILL  FILL_498
timestamp 1711307567
transform 1 0 744 0 1 2170
box -8 -3 16 105
use FILL  FILL_499
timestamp 1711307567
transform 1 0 736 0 1 2170
box -8 -3 16 105
use FILL  FILL_500
timestamp 1711307567
transform 1 0 728 0 1 2170
box -8 -3 16 105
use FILL  FILL_501
timestamp 1711307567
transform 1 0 680 0 1 2170
box -8 -3 16 105
use FILL  FILL_502
timestamp 1711307567
transform 1 0 672 0 1 2170
box -8 -3 16 105
use FILL  FILL_503
timestamp 1711307567
transform 1 0 664 0 1 2170
box -8 -3 16 105
use FILL  FILL_504
timestamp 1711307567
transform 1 0 656 0 1 2170
box -8 -3 16 105
use FILL  FILL_505
timestamp 1711307567
transform 1 0 600 0 1 2170
box -8 -3 16 105
use FILL  FILL_506
timestamp 1711307567
transform 1 0 592 0 1 2170
box -8 -3 16 105
use FILL  FILL_507
timestamp 1711307567
transform 1 0 584 0 1 2170
box -8 -3 16 105
use FILL  FILL_508
timestamp 1711307567
transform 1 0 576 0 1 2170
box -8 -3 16 105
use FILL  FILL_509
timestamp 1711307567
transform 1 0 520 0 1 2170
box -8 -3 16 105
use FILL  FILL_510
timestamp 1711307567
transform 1 0 512 0 1 2170
box -8 -3 16 105
use FILL  FILL_511
timestamp 1711307567
transform 1 0 504 0 1 2170
box -8 -3 16 105
use FILL  FILL_512
timestamp 1711307567
transform 1 0 496 0 1 2170
box -8 -3 16 105
use FILL  FILL_513
timestamp 1711307567
transform 1 0 488 0 1 2170
box -8 -3 16 105
use FILL  FILL_514
timestamp 1711307567
transform 1 0 432 0 1 2170
box -8 -3 16 105
use FILL  FILL_515
timestamp 1711307567
transform 1 0 424 0 1 2170
box -8 -3 16 105
use FILL  FILL_516
timestamp 1711307567
transform 1 0 416 0 1 2170
box -8 -3 16 105
use FILL  FILL_517
timestamp 1711307567
transform 1 0 368 0 1 2170
box -8 -3 16 105
use FILL  FILL_518
timestamp 1711307567
transform 1 0 360 0 1 2170
box -8 -3 16 105
use FILL  FILL_519
timestamp 1711307567
transform 1 0 320 0 1 2170
box -8 -3 16 105
use FILL  FILL_520
timestamp 1711307567
transform 1 0 312 0 1 2170
box -8 -3 16 105
use FILL  FILL_521
timestamp 1711307567
transform 1 0 304 0 1 2170
box -8 -3 16 105
use FILL  FILL_522
timestamp 1711307567
transform 1 0 272 0 1 2170
box -8 -3 16 105
use FILL  FILL_523
timestamp 1711307567
transform 1 0 232 0 1 2170
box -8 -3 16 105
use FILL  FILL_524
timestamp 1711307567
transform 1 0 224 0 1 2170
box -8 -3 16 105
use FILL  FILL_525
timestamp 1711307567
transform 1 0 216 0 1 2170
box -8 -3 16 105
use FILL  FILL_526
timestamp 1711307567
transform 1 0 176 0 1 2170
box -8 -3 16 105
use FILL  FILL_527
timestamp 1711307567
transform 1 0 136 0 1 2170
box -8 -3 16 105
use FILL  FILL_528
timestamp 1711307567
transform 1 0 128 0 1 2170
box -8 -3 16 105
use FILL  FILL_529
timestamp 1711307567
transform 1 0 120 0 1 2170
box -8 -3 16 105
use FILL  FILL_530
timestamp 1711307567
transform 1 0 112 0 1 2170
box -8 -3 16 105
use FILL  FILL_531
timestamp 1711307567
transform 1 0 104 0 1 2170
box -8 -3 16 105
use FILL  FILL_532
timestamp 1711307567
transform 1 0 96 0 1 2170
box -8 -3 16 105
use FILL  FILL_533
timestamp 1711307567
transform 1 0 88 0 1 2170
box -8 -3 16 105
use FILL  FILL_534
timestamp 1711307567
transform 1 0 80 0 1 2170
box -8 -3 16 105
use FILL  FILL_535
timestamp 1711307567
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_536
timestamp 1711307567
transform 1 0 2752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_537
timestamp 1711307567
transform 1 0 2744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_538
timestamp 1711307567
transform 1 0 2656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_539
timestamp 1711307567
transform 1 0 2648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_540
timestamp 1711307567
transform 1 0 2640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_541
timestamp 1711307567
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_542
timestamp 1711307567
transform 1 0 2584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_543
timestamp 1711307567
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_544
timestamp 1711307567
transform 1 0 2536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_545
timestamp 1711307567
transform 1 0 2528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_546
timestamp 1711307567
transform 1 0 2520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_547
timestamp 1711307567
transform 1 0 2512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_548
timestamp 1711307567
transform 1 0 2504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_549
timestamp 1711307567
transform 1 0 2496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_550
timestamp 1711307567
transform 1 0 2440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_551
timestamp 1711307567
transform 1 0 2432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_552
timestamp 1711307567
transform 1 0 2424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_553
timestamp 1711307567
transform 1 0 2416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_554
timestamp 1711307567
transform 1 0 2408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_555
timestamp 1711307567
transform 1 0 2304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_556
timestamp 1711307567
transform 1 0 2264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_557
timestamp 1711307567
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_558
timestamp 1711307567
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_559
timestamp 1711307567
transform 1 0 2208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_560
timestamp 1711307567
transform 1 0 2200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_561
timestamp 1711307567
transform 1 0 2160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_562
timestamp 1711307567
transform 1 0 2136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_563
timestamp 1711307567
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_564
timestamp 1711307567
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_565
timestamp 1711307567
transform 1 0 2072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_566
timestamp 1711307567
transform 1 0 2064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_567
timestamp 1711307567
transform 1 0 2040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_568
timestamp 1711307567
transform 1 0 2032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_569
timestamp 1711307567
transform 1 0 2024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_570
timestamp 1711307567
transform 1 0 1984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_571
timestamp 1711307567
transform 1 0 1976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_572
timestamp 1711307567
transform 1 0 1944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_573
timestamp 1711307567
transform 1 0 1936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_574
timestamp 1711307567
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_575
timestamp 1711307567
transform 1 0 1872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_576
timestamp 1711307567
transform 1 0 1864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_577
timestamp 1711307567
transform 1 0 1856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_578
timestamp 1711307567
transform 1 0 1848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_579
timestamp 1711307567
transform 1 0 1800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_580
timestamp 1711307567
transform 1 0 1792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_581
timestamp 1711307567
transform 1 0 1760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_582
timestamp 1711307567
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_583
timestamp 1711307567
transform 1 0 1712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_584
timestamp 1711307567
transform 1 0 1704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_585
timestamp 1711307567
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_586
timestamp 1711307567
transform 1 0 1672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_587
timestamp 1711307567
transform 1 0 1664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_588
timestamp 1711307567
transform 1 0 1616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_589
timestamp 1711307567
transform 1 0 1608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_590
timestamp 1711307567
transform 1 0 1600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_591
timestamp 1711307567
transform 1 0 1592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_592
timestamp 1711307567
transform 1 0 1584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_593
timestamp 1711307567
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_594
timestamp 1711307567
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_595
timestamp 1711307567
transform 1 0 1520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_596
timestamp 1711307567
transform 1 0 1488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_597
timestamp 1711307567
transform 1 0 1480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_598
timestamp 1711307567
transform 1 0 1472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_599
timestamp 1711307567
transform 1 0 1440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_600
timestamp 1711307567
transform 1 0 1432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_601
timestamp 1711307567
transform 1 0 1424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_602
timestamp 1711307567
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_603
timestamp 1711307567
transform 1 0 1360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_604
timestamp 1711307567
transform 1 0 1352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_605
timestamp 1711307567
transform 1 0 1344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_606
timestamp 1711307567
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_607
timestamp 1711307567
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_608
timestamp 1711307567
transform 1 0 1280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_609
timestamp 1711307567
transform 1 0 1272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_610
timestamp 1711307567
transform 1 0 1264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_611
timestamp 1711307567
transform 1 0 1256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_612
timestamp 1711307567
transform 1 0 1248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_613
timestamp 1711307567
transform 1 0 1240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_614
timestamp 1711307567
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_615
timestamp 1711307567
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_616
timestamp 1711307567
transform 1 0 1184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_617
timestamp 1711307567
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_618
timestamp 1711307567
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_619
timestamp 1711307567
transform 1 0 1136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_620
timestamp 1711307567
transform 1 0 1096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_621
timestamp 1711307567
transform 1 0 1088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_622
timestamp 1711307567
transform 1 0 1080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_623
timestamp 1711307567
transform 1 0 1072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_624
timestamp 1711307567
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_625
timestamp 1711307567
transform 1 0 1016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_626
timestamp 1711307567
transform 1 0 1008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_627
timestamp 1711307567
transform 1 0 1000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_628
timestamp 1711307567
transform 1 0 992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_629
timestamp 1711307567
transform 1 0 984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_630
timestamp 1711307567
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_631
timestamp 1711307567
transform 1 0 936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_632
timestamp 1711307567
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_633
timestamp 1711307567
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_634
timestamp 1711307567
transform 1 0 888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_635
timestamp 1711307567
transform 1 0 856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_636
timestamp 1711307567
transform 1 0 824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_637
timestamp 1711307567
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_638
timestamp 1711307567
transform 1 0 808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_639
timestamp 1711307567
transform 1 0 800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_640
timestamp 1711307567
transform 1 0 760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_641
timestamp 1711307567
transform 1 0 752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_642
timestamp 1711307567
transform 1 0 744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_643
timestamp 1711307567
transform 1 0 712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_644
timestamp 1711307567
transform 1 0 704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_645
timestamp 1711307567
transform 1 0 672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_646
timestamp 1711307567
transform 1 0 664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_647
timestamp 1711307567
transform 1 0 656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_648
timestamp 1711307567
transform 1 0 648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_649
timestamp 1711307567
transform 1 0 592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_650
timestamp 1711307567
transform 1 0 584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_651
timestamp 1711307567
transform 1 0 576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_652
timestamp 1711307567
transform 1 0 568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_653
timestamp 1711307567
transform 1 0 504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_654
timestamp 1711307567
transform 1 0 496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_655
timestamp 1711307567
transform 1 0 488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_656
timestamp 1711307567
transform 1 0 480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_657
timestamp 1711307567
transform 1 0 424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_658
timestamp 1711307567
transform 1 0 416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_659
timestamp 1711307567
transform 1 0 408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_660
timestamp 1711307567
transform 1 0 400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_661
timestamp 1711307567
transform 1 0 392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_662
timestamp 1711307567
transform 1 0 384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_663
timestamp 1711307567
transform 1 0 376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_664
timestamp 1711307567
transform 1 0 328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_665
timestamp 1711307567
transform 1 0 320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_666
timestamp 1711307567
transform 1 0 312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_667
timestamp 1711307567
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_668
timestamp 1711307567
transform 1 0 264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_669
timestamp 1711307567
transform 1 0 256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_670
timestamp 1711307567
transform 1 0 248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_671
timestamp 1711307567
transform 1 0 240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_672
timestamp 1711307567
transform 1 0 208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_673
timestamp 1711307567
transform 1 0 184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_674
timestamp 1711307567
transform 1 0 176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_675
timestamp 1711307567
transform 1 0 168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_676
timestamp 1711307567
transform 1 0 160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_677
timestamp 1711307567
transform 1 0 152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_678
timestamp 1711307567
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_679
timestamp 1711307567
transform 1 0 120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_680
timestamp 1711307567
transform 1 0 112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_681
timestamp 1711307567
transform 1 0 104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_682
timestamp 1711307567
transform 1 0 96 0 -1 2170
box -8 -3 16 105
use FILL  FILL_683
timestamp 1711307567
transform 1 0 88 0 -1 2170
box -8 -3 16 105
use FILL  FILL_684
timestamp 1711307567
transform 1 0 80 0 -1 2170
box -8 -3 16 105
use FILL  FILL_685
timestamp 1711307567
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_686
timestamp 1711307567
transform 1 0 2752 0 1 1970
box -8 -3 16 105
use FILL  FILL_687
timestamp 1711307567
transform 1 0 2720 0 1 1970
box -8 -3 16 105
use FILL  FILL_688
timestamp 1711307567
transform 1 0 2688 0 1 1970
box -8 -3 16 105
use FILL  FILL_689
timestamp 1711307567
transform 1 0 2680 0 1 1970
box -8 -3 16 105
use FILL  FILL_690
timestamp 1711307567
transform 1 0 2640 0 1 1970
box -8 -3 16 105
use FILL  FILL_691
timestamp 1711307567
transform 1 0 2632 0 1 1970
box -8 -3 16 105
use FILL  FILL_692
timestamp 1711307567
transform 1 0 2456 0 1 1970
box -8 -3 16 105
use FILL  FILL_693
timestamp 1711307567
transform 1 0 2352 0 1 1970
box -8 -3 16 105
use FILL  FILL_694
timestamp 1711307567
transform 1 0 2344 0 1 1970
box -8 -3 16 105
use FILL  FILL_695
timestamp 1711307567
transform 1 0 2336 0 1 1970
box -8 -3 16 105
use FILL  FILL_696
timestamp 1711307567
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use FILL  FILL_697
timestamp 1711307567
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use FILL  FILL_698
timestamp 1711307567
transform 1 0 2296 0 1 1970
box -8 -3 16 105
use FILL  FILL_699
timestamp 1711307567
transform 1 0 2288 0 1 1970
box -8 -3 16 105
use FILL  FILL_700
timestamp 1711307567
transform 1 0 2280 0 1 1970
box -8 -3 16 105
use FILL  FILL_701
timestamp 1711307567
transform 1 0 2272 0 1 1970
box -8 -3 16 105
use FILL  FILL_702
timestamp 1711307567
transform 1 0 2264 0 1 1970
box -8 -3 16 105
use FILL  FILL_703
timestamp 1711307567
transform 1 0 2208 0 1 1970
box -8 -3 16 105
use FILL  FILL_704
timestamp 1711307567
transform 1 0 2200 0 1 1970
box -8 -3 16 105
use FILL  FILL_705
timestamp 1711307567
transform 1 0 2192 0 1 1970
box -8 -3 16 105
use FILL  FILL_706
timestamp 1711307567
transform 1 0 2184 0 1 1970
box -8 -3 16 105
use FILL  FILL_707
timestamp 1711307567
transform 1 0 2176 0 1 1970
box -8 -3 16 105
use FILL  FILL_708
timestamp 1711307567
transform 1 0 2136 0 1 1970
box -8 -3 16 105
use FILL  FILL_709
timestamp 1711307567
transform 1 0 2128 0 1 1970
box -8 -3 16 105
use FILL  FILL_710
timestamp 1711307567
transform 1 0 2120 0 1 1970
box -8 -3 16 105
use FILL  FILL_711
timestamp 1711307567
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_712
timestamp 1711307567
transform 1 0 2072 0 1 1970
box -8 -3 16 105
use FILL  FILL_713
timestamp 1711307567
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use FILL  FILL_714
timestamp 1711307567
transform 1 0 2024 0 1 1970
box -8 -3 16 105
use FILL  FILL_715
timestamp 1711307567
transform 1 0 2016 0 1 1970
box -8 -3 16 105
use FILL  FILL_716
timestamp 1711307567
transform 1 0 2008 0 1 1970
box -8 -3 16 105
use FILL  FILL_717
timestamp 1711307567
transform 1 0 1968 0 1 1970
box -8 -3 16 105
use FILL  FILL_718
timestamp 1711307567
transform 1 0 1960 0 1 1970
box -8 -3 16 105
use FILL  FILL_719
timestamp 1711307567
transform 1 0 1920 0 1 1970
box -8 -3 16 105
use FILL  FILL_720
timestamp 1711307567
transform 1 0 1912 0 1 1970
box -8 -3 16 105
use FILL  FILL_721
timestamp 1711307567
transform 1 0 1904 0 1 1970
box -8 -3 16 105
use FILL  FILL_722
timestamp 1711307567
transform 1 0 1896 0 1 1970
box -8 -3 16 105
use FILL  FILL_723
timestamp 1711307567
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_724
timestamp 1711307567
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_725
timestamp 1711307567
transform 1 0 1832 0 1 1970
box -8 -3 16 105
use FILL  FILL_726
timestamp 1711307567
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_727
timestamp 1711307567
transform 1 0 1784 0 1 1970
box -8 -3 16 105
use FILL  FILL_728
timestamp 1711307567
transform 1 0 1752 0 1 1970
box -8 -3 16 105
use FILL  FILL_729
timestamp 1711307567
transform 1 0 1728 0 1 1970
box -8 -3 16 105
use FILL  FILL_730
timestamp 1711307567
transform 1 0 1720 0 1 1970
box -8 -3 16 105
use FILL  FILL_731
timestamp 1711307567
transform 1 0 1712 0 1 1970
box -8 -3 16 105
use FILL  FILL_732
timestamp 1711307567
transform 1 0 1704 0 1 1970
box -8 -3 16 105
use FILL  FILL_733
timestamp 1711307567
transform 1 0 1648 0 1 1970
box -8 -3 16 105
use FILL  FILL_734
timestamp 1711307567
transform 1 0 1640 0 1 1970
box -8 -3 16 105
use FILL  FILL_735
timestamp 1711307567
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use FILL  FILL_736
timestamp 1711307567
transform 1 0 1624 0 1 1970
box -8 -3 16 105
use FILL  FILL_737
timestamp 1711307567
transform 1 0 1576 0 1 1970
box -8 -3 16 105
use FILL  FILL_738
timestamp 1711307567
transform 1 0 1552 0 1 1970
box -8 -3 16 105
use FILL  FILL_739
timestamp 1711307567
transform 1 0 1544 0 1 1970
box -8 -3 16 105
use FILL  FILL_740
timestamp 1711307567
transform 1 0 1536 0 1 1970
box -8 -3 16 105
use FILL  FILL_741
timestamp 1711307567
transform 1 0 1528 0 1 1970
box -8 -3 16 105
use FILL  FILL_742
timestamp 1711307567
transform 1 0 1472 0 1 1970
box -8 -3 16 105
use FILL  FILL_743
timestamp 1711307567
transform 1 0 1464 0 1 1970
box -8 -3 16 105
use FILL  FILL_744
timestamp 1711307567
transform 1 0 1456 0 1 1970
box -8 -3 16 105
use FILL  FILL_745
timestamp 1711307567
transform 1 0 1448 0 1 1970
box -8 -3 16 105
use FILL  FILL_746
timestamp 1711307567
transform 1 0 1392 0 1 1970
box -8 -3 16 105
use FILL  FILL_747
timestamp 1711307567
transform 1 0 1384 0 1 1970
box -8 -3 16 105
use FILL  FILL_748
timestamp 1711307567
transform 1 0 1376 0 1 1970
box -8 -3 16 105
use FILL  FILL_749
timestamp 1711307567
transform 1 0 1368 0 1 1970
box -8 -3 16 105
use FILL  FILL_750
timestamp 1711307567
transform 1 0 1312 0 1 1970
box -8 -3 16 105
use FILL  FILL_751
timestamp 1711307567
transform 1 0 1304 0 1 1970
box -8 -3 16 105
use FILL  FILL_752
timestamp 1711307567
transform 1 0 1296 0 1 1970
box -8 -3 16 105
use FILL  FILL_753
timestamp 1711307567
transform 1 0 1288 0 1 1970
box -8 -3 16 105
use FILL  FILL_754
timestamp 1711307567
transform 1 0 1248 0 1 1970
box -8 -3 16 105
use FILL  FILL_755
timestamp 1711307567
transform 1 0 1240 0 1 1970
box -8 -3 16 105
use FILL  FILL_756
timestamp 1711307567
transform 1 0 1232 0 1 1970
box -8 -3 16 105
use FILL  FILL_757
timestamp 1711307567
transform 1 0 1192 0 1 1970
box -8 -3 16 105
use FILL  FILL_758
timestamp 1711307567
transform 1 0 1184 0 1 1970
box -8 -3 16 105
use FILL  FILL_759
timestamp 1711307567
transform 1 0 1176 0 1 1970
box -8 -3 16 105
use FILL  FILL_760
timestamp 1711307567
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_761
timestamp 1711307567
transform 1 0 1144 0 1 1970
box -8 -3 16 105
use FILL  FILL_762
timestamp 1711307567
transform 1 0 1112 0 1 1970
box -8 -3 16 105
use FILL  FILL_763
timestamp 1711307567
transform 1 0 1104 0 1 1970
box -8 -3 16 105
use FILL  FILL_764
timestamp 1711307567
transform 1 0 1096 0 1 1970
box -8 -3 16 105
use FILL  FILL_765
timestamp 1711307567
transform 1 0 1088 0 1 1970
box -8 -3 16 105
use FILL  FILL_766
timestamp 1711307567
transform 1 0 1080 0 1 1970
box -8 -3 16 105
use FILL  FILL_767
timestamp 1711307567
transform 1 0 1032 0 1 1970
box -8 -3 16 105
use FILL  FILL_768
timestamp 1711307567
transform 1 0 1024 0 1 1970
box -8 -3 16 105
use FILL  FILL_769
timestamp 1711307567
transform 1 0 1016 0 1 1970
box -8 -3 16 105
use FILL  FILL_770
timestamp 1711307567
transform 1 0 1008 0 1 1970
box -8 -3 16 105
use FILL  FILL_771
timestamp 1711307567
transform 1 0 1000 0 1 1970
box -8 -3 16 105
use FILL  FILL_772
timestamp 1711307567
transform 1 0 968 0 1 1970
box -8 -3 16 105
use FILL  FILL_773
timestamp 1711307567
transform 1 0 960 0 1 1970
box -8 -3 16 105
use FILL  FILL_774
timestamp 1711307567
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_775
timestamp 1711307567
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_776
timestamp 1711307567
transform 1 0 912 0 1 1970
box -8 -3 16 105
use FILL  FILL_777
timestamp 1711307567
transform 1 0 904 0 1 1970
box -8 -3 16 105
use FILL  FILL_778
timestamp 1711307567
transform 1 0 856 0 1 1970
box -8 -3 16 105
use FILL  FILL_779
timestamp 1711307567
transform 1 0 848 0 1 1970
box -8 -3 16 105
use FILL  FILL_780
timestamp 1711307567
transform 1 0 840 0 1 1970
box -8 -3 16 105
use FILL  FILL_781
timestamp 1711307567
transform 1 0 832 0 1 1970
box -8 -3 16 105
use FILL  FILL_782
timestamp 1711307567
transform 1 0 824 0 1 1970
box -8 -3 16 105
use FILL  FILL_783
timestamp 1711307567
transform 1 0 760 0 1 1970
box -8 -3 16 105
use FILL  FILL_784
timestamp 1711307567
transform 1 0 752 0 1 1970
box -8 -3 16 105
use FILL  FILL_785
timestamp 1711307567
transform 1 0 744 0 1 1970
box -8 -3 16 105
use FILL  FILL_786
timestamp 1711307567
transform 1 0 712 0 1 1970
box -8 -3 16 105
use FILL  FILL_787
timestamp 1711307567
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FILL  FILL_788
timestamp 1711307567
transform 1 0 656 0 1 1970
box -8 -3 16 105
use FILL  FILL_789
timestamp 1711307567
transform 1 0 648 0 1 1970
box -8 -3 16 105
use FILL  FILL_790
timestamp 1711307567
transform 1 0 640 0 1 1970
box -8 -3 16 105
use FILL  FILL_791
timestamp 1711307567
transform 1 0 632 0 1 1970
box -8 -3 16 105
use FILL  FILL_792
timestamp 1711307567
transform 1 0 624 0 1 1970
box -8 -3 16 105
use FILL  FILL_793
timestamp 1711307567
transform 1 0 584 0 1 1970
box -8 -3 16 105
use FILL  FILL_794
timestamp 1711307567
transform 1 0 576 0 1 1970
box -8 -3 16 105
use FILL  FILL_795
timestamp 1711307567
transform 1 0 568 0 1 1970
box -8 -3 16 105
use FILL  FILL_796
timestamp 1711307567
transform 1 0 560 0 1 1970
box -8 -3 16 105
use FILL  FILL_797
timestamp 1711307567
transform 1 0 520 0 1 1970
box -8 -3 16 105
use FILL  FILL_798
timestamp 1711307567
transform 1 0 512 0 1 1970
box -8 -3 16 105
use FILL  FILL_799
timestamp 1711307567
transform 1 0 504 0 1 1970
box -8 -3 16 105
use FILL  FILL_800
timestamp 1711307567
transform 1 0 496 0 1 1970
box -8 -3 16 105
use FILL  FILL_801
timestamp 1711307567
transform 1 0 472 0 1 1970
box -8 -3 16 105
use FILL  FILL_802
timestamp 1711307567
transform 1 0 440 0 1 1970
box -8 -3 16 105
use FILL  FILL_803
timestamp 1711307567
transform 1 0 432 0 1 1970
box -8 -3 16 105
use FILL  FILL_804
timestamp 1711307567
transform 1 0 408 0 1 1970
box -8 -3 16 105
use FILL  FILL_805
timestamp 1711307567
transform 1 0 400 0 1 1970
box -8 -3 16 105
use FILL  FILL_806
timestamp 1711307567
transform 1 0 352 0 1 1970
box -8 -3 16 105
use FILL  FILL_807
timestamp 1711307567
transform 1 0 344 0 1 1970
box -8 -3 16 105
use FILL  FILL_808
timestamp 1711307567
transform 1 0 336 0 1 1970
box -8 -3 16 105
use FILL  FILL_809
timestamp 1711307567
transform 1 0 328 0 1 1970
box -8 -3 16 105
use FILL  FILL_810
timestamp 1711307567
transform 1 0 288 0 1 1970
box -8 -3 16 105
use FILL  FILL_811
timestamp 1711307567
transform 1 0 280 0 1 1970
box -8 -3 16 105
use FILL  FILL_812
timestamp 1711307567
transform 1 0 248 0 1 1970
box -8 -3 16 105
use FILL  FILL_813
timestamp 1711307567
transform 1 0 240 0 1 1970
box -8 -3 16 105
use FILL  FILL_814
timestamp 1711307567
transform 1 0 232 0 1 1970
box -8 -3 16 105
use FILL  FILL_815
timestamp 1711307567
transform 1 0 208 0 1 1970
box -8 -3 16 105
use FILL  FILL_816
timestamp 1711307567
transform 1 0 200 0 1 1970
box -8 -3 16 105
use FILL  FILL_817
timestamp 1711307567
transform 1 0 192 0 1 1970
box -8 -3 16 105
use FILL  FILL_818
timestamp 1711307567
transform 1 0 184 0 1 1970
box -8 -3 16 105
use FILL  FILL_819
timestamp 1711307567
transform 1 0 176 0 1 1970
box -8 -3 16 105
use FILL  FILL_820
timestamp 1711307567
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_821
timestamp 1711307567
transform 1 0 2752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_822
timestamp 1711307567
transform 1 0 2744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_823
timestamp 1711307567
transform 1 0 2680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_824
timestamp 1711307567
transform 1 0 2672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_825
timestamp 1711307567
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_826
timestamp 1711307567
transform 1 0 2592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_827
timestamp 1711307567
transform 1 0 2584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_828
timestamp 1711307567
transform 1 0 2432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_829
timestamp 1711307567
transform 1 0 2424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_830
timestamp 1711307567
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_831
timestamp 1711307567
transform 1 0 2408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_832
timestamp 1711307567
transform 1 0 2400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_833
timestamp 1711307567
transform 1 0 2344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_834
timestamp 1711307567
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_835
timestamp 1711307567
transform 1 0 2328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_836
timestamp 1711307567
transform 1 0 2272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_837
timestamp 1711307567
transform 1 0 2264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_838
timestamp 1711307567
transform 1 0 2256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_839
timestamp 1711307567
transform 1 0 2248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_840
timestamp 1711307567
transform 1 0 2184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_841
timestamp 1711307567
transform 1 0 2176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_842
timestamp 1711307567
transform 1 0 2152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_843
timestamp 1711307567
transform 1 0 2144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_844
timestamp 1711307567
transform 1 0 2088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_845
timestamp 1711307567
transform 1 0 2080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_846
timestamp 1711307567
transform 1 0 2072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_847
timestamp 1711307567
transform 1 0 2040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_848
timestamp 1711307567
transform 1 0 2008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_849
timestamp 1711307567
transform 1 0 2000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_850
timestamp 1711307567
transform 1 0 1992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_851
timestamp 1711307567
transform 1 0 1968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_852
timestamp 1711307567
transform 1 0 1960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_853
timestamp 1711307567
transform 1 0 1928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_854
timestamp 1711307567
transform 1 0 1896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_855
timestamp 1711307567
transform 1 0 1888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_856
timestamp 1711307567
transform 1 0 1880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_857
timestamp 1711307567
transform 1 0 1824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_858
timestamp 1711307567
transform 1 0 1816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_859
timestamp 1711307567
transform 1 0 1808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_860
timestamp 1711307567
transform 1 0 1800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_861
timestamp 1711307567
transform 1 0 1792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_862
timestamp 1711307567
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_863
timestamp 1711307567
transform 1 0 1736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_864
timestamp 1711307567
transform 1 0 1728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_865
timestamp 1711307567
transform 1 0 1696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_866
timestamp 1711307567
transform 1 0 1688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_867
timestamp 1711307567
transform 1 0 1680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_868
timestamp 1711307567
transform 1 0 1648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_869
timestamp 1711307567
transform 1 0 1640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_870
timestamp 1711307567
transform 1 0 1632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_871
timestamp 1711307567
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_872
timestamp 1711307567
transform 1 0 1592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_873
timestamp 1711307567
transform 1 0 1584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_874
timestamp 1711307567
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_875
timestamp 1711307567
transform 1 0 1552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_876
timestamp 1711307567
transform 1 0 1544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_877
timestamp 1711307567
transform 1 0 1504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_878
timestamp 1711307567
transform 1 0 1496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_879
timestamp 1711307567
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_880
timestamp 1711307567
transform 1 0 1480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_881
timestamp 1711307567
transform 1 0 1448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_882
timestamp 1711307567
transform 1 0 1440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_883
timestamp 1711307567
transform 1 0 1400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_884
timestamp 1711307567
transform 1 0 1392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_885
timestamp 1711307567
transform 1 0 1384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_886
timestamp 1711307567
transform 1 0 1376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_887
timestamp 1711307567
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_888
timestamp 1711307567
transform 1 0 1360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_889
timestamp 1711307567
transform 1 0 1312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_890
timestamp 1711307567
transform 1 0 1304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_891
timestamp 1711307567
transform 1 0 1296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_892
timestamp 1711307567
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_893
timestamp 1711307567
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_894
timestamp 1711307567
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_895
timestamp 1711307567
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_896
timestamp 1711307567
transform 1 0 1224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_897
timestamp 1711307567
transform 1 0 1216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_898
timestamp 1711307567
transform 1 0 1208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_899
timestamp 1711307567
transform 1 0 1200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_900
timestamp 1711307567
transform 1 0 1192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_901
timestamp 1711307567
transform 1 0 1160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_902
timestamp 1711307567
transform 1 0 1152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_903
timestamp 1711307567
transform 1 0 1144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_904
timestamp 1711307567
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_905
timestamp 1711307567
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_906
timestamp 1711307567
transform 1 0 1096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_907
timestamp 1711307567
transform 1 0 1088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_908
timestamp 1711307567
transform 1 0 1080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_909
timestamp 1711307567
transform 1 0 1048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_910
timestamp 1711307567
transform 1 0 1040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_911
timestamp 1711307567
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_912
timestamp 1711307567
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_913
timestamp 1711307567
transform 1 0 984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_914
timestamp 1711307567
transform 1 0 976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_915
timestamp 1711307567
transform 1 0 968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_916
timestamp 1711307567
transform 1 0 960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_917
timestamp 1711307567
transform 1 0 952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_918
timestamp 1711307567
transform 1 0 912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_919
timestamp 1711307567
transform 1 0 904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_920
timestamp 1711307567
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_921
timestamp 1711307567
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_922
timestamp 1711307567
transform 1 0 880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_923
timestamp 1711307567
transform 1 0 872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_924
timestamp 1711307567
transform 1 0 824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_925
timestamp 1711307567
transform 1 0 816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_926
timestamp 1711307567
transform 1 0 808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_927
timestamp 1711307567
transform 1 0 800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_928
timestamp 1711307567
transform 1 0 792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_929
timestamp 1711307567
transform 1 0 752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_930
timestamp 1711307567
transform 1 0 744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_931
timestamp 1711307567
transform 1 0 736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_932
timestamp 1711307567
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_933
timestamp 1711307567
transform 1 0 688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_934
timestamp 1711307567
transform 1 0 680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_935
timestamp 1711307567
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_936
timestamp 1711307567
transform 1 0 632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_937
timestamp 1711307567
transform 1 0 624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_938
timestamp 1711307567
transform 1 0 568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_939
timestamp 1711307567
transform 1 0 560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_940
timestamp 1711307567
transform 1 0 552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_941
timestamp 1711307567
transform 1 0 544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_942
timestamp 1711307567
transform 1 0 512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_943
timestamp 1711307567
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_944
timestamp 1711307567
transform 1 0 464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_945
timestamp 1711307567
transform 1 0 456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_946
timestamp 1711307567
transform 1 0 448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_947
timestamp 1711307567
transform 1 0 392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_948
timestamp 1711307567
transform 1 0 384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_949
timestamp 1711307567
transform 1 0 376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_950
timestamp 1711307567
transform 1 0 368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_951
timestamp 1711307567
transform 1 0 360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_952
timestamp 1711307567
transform 1 0 312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_953
timestamp 1711307567
transform 1 0 304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_954
timestamp 1711307567
transform 1 0 264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_955
timestamp 1711307567
transform 1 0 256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_956
timestamp 1711307567
transform 1 0 248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_957
timestamp 1711307567
transform 1 0 240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_958
timestamp 1711307567
transform 1 0 168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_959
timestamp 1711307567
transform 1 0 160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_960
timestamp 1711307567
transform 1 0 152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_961
timestamp 1711307567
transform 1 0 144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_962
timestamp 1711307567
transform 1 0 136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_963
timestamp 1711307567
transform 1 0 128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_964
timestamp 1711307567
transform 1 0 120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_965
timestamp 1711307567
transform 1 0 112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_966
timestamp 1711307567
transform 1 0 104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_967
timestamp 1711307567
transform 1 0 96 0 -1 1970
box -8 -3 16 105
use FILL  FILL_968
timestamp 1711307567
transform 1 0 88 0 -1 1970
box -8 -3 16 105
use FILL  FILL_969
timestamp 1711307567
transform 1 0 80 0 -1 1970
box -8 -3 16 105
use FILL  FILL_970
timestamp 1711307567
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_971
timestamp 1711307567
transform 1 0 2752 0 1 1770
box -8 -3 16 105
use FILL  FILL_972
timestamp 1711307567
transform 1 0 2744 0 1 1770
box -8 -3 16 105
use FILL  FILL_973
timestamp 1711307567
transform 1 0 2696 0 1 1770
box -8 -3 16 105
use FILL  FILL_974
timestamp 1711307567
transform 1 0 2672 0 1 1770
box -8 -3 16 105
use FILL  FILL_975
timestamp 1711307567
transform 1 0 2664 0 1 1770
box -8 -3 16 105
use FILL  FILL_976
timestamp 1711307567
transform 1 0 2608 0 1 1770
box -8 -3 16 105
use FILL  FILL_977
timestamp 1711307567
transform 1 0 2600 0 1 1770
box -8 -3 16 105
use FILL  FILL_978
timestamp 1711307567
transform 1 0 2528 0 1 1770
box -8 -3 16 105
use FILL  FILL_979
timestamp 1711307567
transform 1 0 2520 0 1 1770
box -8 -3 16 105
use FILL  FILL_980
timestamp 1711307567
transform 1 0 2416 0 1 1770
box -8 -3 16 105
use FILL  FILL_981
timestamp 1711307567
transform 1 0 2408 0 1 1770
box -8 -3 16 105
use FILL  FILL_982
timestamp 1711307567
transform 1 0 2400 0 1 1770
box -8 -3 16 105
use FILL  FILL_983
timestamp 1711307567
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use FILL  FILL_984
timestamp 1711307567
transform 1 0 2336 0 1 1770
box -8 -3 16 105
use FILL  FILL_985
timestamp 1711307567
transform 1 0 2328 0 1 1770
box -8 -3 16 105
use FILL  FILL_986
timestamp 1711307567
transform 1 0 2320 0 1 1770
box -8 -3 16 105
use FILL  FILL_987
timestamp 1711307567
transform 1 0 2312 0 1 1770
box -8 -3 16 105
use FILL  FILL_988
timestamp 1711307567
transform 1 0 2256 0 1 1770
box -8 -3 16 105
use FILL  FILL_989
timestamp 1711307567
transform 1 0 2248 0 1 1770
box -8 -3 16 105
use FILL  FILL_990
timestamp 1711307567
transform 1 0 2240 0 1 1770
box -8 -3 16 105
use FILL  FILL_991
timestamp 1711307567
transform 1 0 2232 0 1 1770
box -8 -3 16 105
use FILL  FILL_992
timestamp 1711307567
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_993
timestamp 1711307567
transform 1 0 2152 0 1 1770
box -8 -3 16 105
use FILL  FILL_994
timestamp 1711307567
transform 1 0 2144 0 1 1770
box -8 -3 16 105
use FILL  FILL_995
timestamp 1711307567
transform 1 0 2136 0 1 1770
box -8 -3 16 105
use FILL  FILL_996
timestamp 1711307567
transform 1 0 2096 0 1 1770
box -8 -3 16 105
use FILL  FILL_997
timestamp 1711307567
transform 1 0 2088 0 1 1770
box -8 -3 16 105
use FILL  FILL_998
timestamp 1711307567
transform 1 0 2080 0 1 1770
box -8 -3 16 105
use FILL  FILL_999
timestamp 1711307567
transform 1 0 2032 0 1 1770
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1711307567
transform 1 0 2024 0 1 1770
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1711307567
transform 1 0 2016 0 1 1770
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1711307567
transform 1 0 2008 0 1 1770
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1711307567
transform 1 0 1944 0 1 1770
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1711307567
transform 1 0 1936 0 1 1770
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1711307567
transform 1 0 1928 0 1 1770
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1711307567
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1711307567
transform 1 0 1856 0 1 1770
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1711307567
transform 1 0 1848 0 1 1770
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1711307567
transform 1 0 1840 0 1 1770
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1711307567
transform 1 0 1832 0 1 1770
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1711307567
transform 1 0 1776 0 1 1770
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1711307567
transform 1 0 1736 0 1 1770
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1711307567
transform 1 0 1704 0 1 1770
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1711307567
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1711307567
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1711307567
transform 1 0 1664 0 1 1770
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1711307567
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1711307567
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1711307567
transform 1 0 1608 0 1 1770
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1711307567
transform 1 0 1600 0 1 1770
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1711307567
transform 1 0 1560 0 1 1770
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1711307567
transform 1 0 1528 0 1 1770
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1711307567
transform 1 0 1520 0 1 1770
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1711307567
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1711307567
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1711307567
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1711307567
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1711307567
transform 1 0 1424 0 1 1770
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1711307567
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1711307567
transform 1 0 1384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1711307567
transform 1 0 1344 0 1 1770
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1711307567
transform 1 0 1336 0 1 1770
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1711307567
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1711307567
transform 1 0 1320 0 1 1770
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1711307567
transform 1 0 1312 0 1 1770
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1711307567
transform 1 0 1264 0 1 1770
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1711307567
transform 1 0 1256 0 1 1770
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1711307567
transform 1 0 1248 0 1 1770
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1711307567
transform 1 0 1240 0 1 1770
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1711307567
transform 1 0 1232 0 1 1770
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1711307567
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1711307567
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1711307567
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1711307567
transform 1 0 1168 0 1 1770
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1711307567
transform 1 0 1160 0 1 1770
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1711307567
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1711307567
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1711307567
transform 1 0 1104 0 1 1770
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1711307567
transform 1 0 1080 0 1 1770
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1711307567
transform 1 0 1072 0 1 1770
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1711307567
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1711307567
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1711307567
transform 1 0 1032 0 1 1770
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1711307567
transform 1 0 1024 0 1 1770
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1711307567
transform 1 0 992 0 1 1770
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1711307567
transform 1 0 984 0 1 1770
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1711307567
transform 1 0 976 0 1 1770
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1711307567
transform 1 0 968 0 1 1770
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1711307567
transform 1 0 928 0 1 1770
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1711307567
transform 1 0 920 0 1 1770
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1711307567
transform 1 0 912 0 1 1770
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1711307567
transform 1 0 888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1711307567
transform 1 0 880 0 1 1770
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1711307567
transform 1 0 872 0 1 1770
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1711307567
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1711307567
transform 1 0 832 0 1 1770
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1711307567
transform 1 0 824 0 1 1770
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1711307567
transform 1 0 816 0 1 1770
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1711307567
transform 1 0 808 0 1 1770
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1711307567
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1711307567
transform 1 0 768 0 1 1770
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1711307567
transform 1 0 760 0 1 1770
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1711307567
transform 1 0 752 0 1 1770
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1711307567
transform 1 0 744 0 1 1770
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1711307567
transform 1 0 712 0 1 1770
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1711307567
transform 1 0 704 0 1 1770
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1711307567
transform 1 0 696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1711307567
transform 1 0 688 0 1 1770
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1711307567
transform 1 0 648 0 1 1770
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1711307567
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1711307567
transform 1 0 632 0 1 1770
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1711307567
transform 1 0 624 0 1 1770
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1711307567
transform 1 0 616 0 1 1770
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1711307567
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1711307567
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1711307567
transform 1 0 560 0 1 1770
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1711307567
transform 1 0 552 0 1 1770
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1711307567
transform 1 0 544 0 1 1770
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1711307567
transform 1 0 536 0 1 1770
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1711307567
transform 1 0 528 0 1 1770
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1711307567
transform 1 0 496 0 1 1770
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1711307567
transform 1 0 488 0 1 1770
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1711307567
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1711307567
transform 1 0 440 0 1 1770
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1711307567
transform 1 0 432 0 1 1770
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1711307567
transform 1 0 392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1711307567
transform 1 0 384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1711307567
transform 1 0 376 0 1 1770
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1711307567
transform 1 0 368 0 1 1770
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1711307567
transform 1 0 360 0 1 1770
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1711307567
transform 1 0 328 0 1 1770
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1711307567
transform 1 0 320 0 1 1770
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1711307567
transform 1 0 312 0 1 1770
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1711307567
transform 1 0 280 0 1 1770
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1711307567
transform 1 0 272 0 1 1770
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1711307567
transform 1 0 232 0 1 1770
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1711307567
transform 1 0 224 0 1 1770
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1711307567
transform 1 0 216 0 1 1770
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1711307567
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1711307567
transform 1 0 168 0 1 1770
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1711307567
transform 1 0 160 0 1 1770
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1711307567
transform 1 0 152 0 1 1770
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1711307567
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1711307567
transform 1 0 120 0 1 1770
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1711307567
transform 1 0 112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1711307567
transform 1 0 104 0 1 1770
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1711307567
transform 1 0 96 0 1 1770
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1711307567
transform 1 0 88 0 1 1770
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1711307567
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1711307567
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1711307567
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1711307567
transform 1 0 2744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1711307567
transform 1 0 2696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1711307567
transform 1 0 2688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1711307567
transform 1 0 2640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1711307567
transform 1 0 2632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1711307567
transform 1 0 2600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1711307567
transform 1 0 2592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1711307567
transform 1 0 2568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1711307567
transform 1 0 2560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1711307567
transform 1 0 2456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1711307567
transform 1 0 2448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1711307567
transform 1 0 2440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1711307567
transform 1 0 2432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1711307567
transform 1 0 2424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1711307567
transform 1 0 2368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1711307567
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1711307567
transform 1 0 2352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1711307567
transform 1 0 2312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1711307567
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1711307567
transform 1 0 2296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1711307567
transform 1 0 2256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1711307567
transform 1 0 2248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1711307567
transform 1 0 2208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1711307567
transform 1 0 2200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1711307567
transform 1 0 2192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1711307567
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1711307567
transform 1 0 2152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1711307567
transform 1 0 2144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1711307567
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1711307567
transform 1 0 2104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1711307567
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1711307567
transform 1 0 2056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1711307567
transform 1 0 2048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1711307567
transform 1 0 2040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1711307567
transform 1 0 2008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1711307567
transform 1 0 2000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1711307567
transform 1 0 1992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1711307567
transform 1 0 1984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1711307567
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1711307567
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1711307567
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1711307567
transform 1 0 1920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1711307567
transform 1 0 1872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1711307567
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1711307567
transform 1 0 1856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1711307567
transform 1 0 1824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1711307567
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1711307567
transform 1 0 1792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1711307567
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1711307567
transform 1 0 1744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1711307567
transform 1 0 1736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1711307567
transform 1 0 1728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1711307567
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1711307567
transform 1 0 1688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1711307567
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1711307567
transform 1 0 1656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1711307567
transform 1 0 1632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1711307567
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1711307567
transform 1 0 1600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1711307567
transform 1 0 1592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1711307567
transform 1 0 1584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1711307567
transform 1 0 1536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1711307567
transform 1 0 1528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1711307567
transform 1 0 1520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1711307567
transform 1 0 1512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1711307567
transform 1 0 1504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1711307567
transform 1 0 1464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1711307567
transform 1 0 1456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1711307567
transform 1 0 1448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1711307567
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1711307567
transform 1 0 1400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1711307567
transform 1 0 1360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1711307567
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1711307567
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1711307567
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1711307567
transform 1 0 1296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1711307567
transform 1 0 1288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1711307567
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1711307567
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1711307567
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1711307567
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1711307567
transform 1 0 1200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1711307567
transform 1 0 1192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1711307567
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1711307567
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1711307567
transform 1 0 1144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1711307567
transform 1 0 1136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1711307567
transform 1 0 1128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1711307567
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1711307567
transform 1 0 1080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1711307567
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1711307567
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1711307567
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1711307567
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1711307567
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1711307567
transform 1 0 1000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1711307567
transform 1 0 992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1711307567
transform 1 0 968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1711307567
transform 1 0 960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1711307567
transform 1 0 952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1711307567
transform 1 0 944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1711307567
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1711307567
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1711307567
transform 1 0 888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1711307567
transform 1 0 880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1711307567
transform 1 0 856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1711307567
transform 1 0 848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1711307567
transform 1 0 816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1711307567
transform 1 0 808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1711307567
transform 1 0 800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1711307567
transform 1 0 792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1711307567
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1711307567
transform 1 0 752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1711307567
transform 1 0 744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1711307567
transform 1 0 736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1711307567
transform 1 0 704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1711307567
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1711307567
transform 1 0 656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1711307567
transform 1 0 648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1711307567
transform 1 0 640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1711307567
transform 1 0 632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1711307567
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1711307567
transform 1 0 584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1711307567
transform 1 0 576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1711307567
transform 1 0 568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1711307567
transform 1 0 536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1711307567
transform 1 0 528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1711307567
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1711307567
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1711307567
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1711307567
transform 1 0 440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1711307567
transform 1 0 432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1711307567
transform 1 0 424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1711307567
transform 1 0 416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1711307567
transform 1 0 376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1711307567
transform 1 0 368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1711307567
transform 1 0 360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1711307567
transform 1 0 352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1711307567
transform 1 0 288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1711307567
transform 1 0 280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1711307567
transform 1 0 272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1711307567
transform 1 0 264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1711307567
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1711307567
transform 1 0 232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1711307567
transform 1 0 224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1711307567
transform 1 0 216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1711307567
transform 1 0 208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1711307567
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1711307567
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1711307567
transform 1 0 88 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1711307567
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1711307567
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1711307567
transform 1 0 2752 0 1 1570
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1711307567
transform 1 0 2744 0 1 1570
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1711307567
transform 1 0 2680 0 1 1570
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1711307567
transform 1 0 2672 0 1 1570
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1711307567
transform 1 0 2584 0 1 1570
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1711307567
transform 1 0 2576 0 1 1570
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1711307567
transform 1 0 2568 0 1 1570
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1711307567
transform 1 0 2504 0 1 1570
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1711307567
transform 1 0 2400 0 1 1570
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1711307567
transform 1 0 2392 0 1 1570
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1711307567
transform 1 0 2384 0 1 1570
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1711307567
transform 1 0 2336 0 1 1570
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1711307567
transform 1 0 2328 0 1 1570
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1711307567
transform 1 0 2288 0 1 1570
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1711307567
transform 1 0 2248 0 1 1570
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1711307567
transform 1 0 2240 0 1 1570
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1711307567
transform 1 0 2232 0 1 1570
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1711307567
transform 1 0 2200 0 1 1570
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1711307567
transform 1 0 2192 0 1 1570
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1711307567
transform 1 0 2152 0 1 1570
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1711307567
transform 1 0 2144 0 1 1570
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1711307567
transform 1 0 2112 0 1 1570
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1711307567
transform 1 0 2104 0 1 1570
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1711307567
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1711307567
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1711307567
transform 1 0 2064 0 1 1570
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1711307567
transform 1 0 2032 0 1 1570
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1711307567
transform 1 0 1992 0 1 1570
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1711307567
transform 1 0 1984 0 1 1570
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1711307567
transform 1 0 1976 0 1 1570
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1711307567
transform 1 0 1944 0 1 1570
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1711307567
transform 1 0 1936 0 1 1570
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1711307567
transform 1 0 1928 0 1 1570
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1711307567
transform 1 0 1920 0 1 1570
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1711307567
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1711307567
transform 1 0 1856 0 1 1570
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1711307567
transform 1 0 1848 0 1 1570
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1711307567
transform 1 0 1800 0 1 1570
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1711307567
transform 1 0 1792 0 1 1570
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1711307567
transform 1 0 1784 0 1 1570
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1711307567
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1711307567
transform 1 0 1728 0 1 1570
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1711307567
transform 1 0 1720 0 1 1570
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1711307567
transform 1 0 1712 0 1 1570
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1711307567
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1711307567
transform 1 0 1640 0 1 1570
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1711307567
transform 1 0 1632 0 1 1570
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1711307567
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1711307567
transform 1 0 1592 0 1 1570
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1711307567
transform 1 0 1584 0 1 1570
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1711307567
transform 1 0 1544 0 1 1570
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1711307567
transform 1 0 1536 0 1 1570
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1711307567
transform 1 0 1528 0 1 1570
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1711307567
transform 1 0 1520 0 1 1570
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1711307567
transform 1 0 1496 0 1 1570
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1711307567
transform 1 0 1456 0 1 1570
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1711307567
transform 1 0 1448 0 1 1570
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1711307567
transform 1 0 1440 0 1 1570
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1711307567
transform 1 0 1432 0 1 1570
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1711307567
transform 1 0 1400 0 1 1570
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1711307567
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1711307567
transform 1 0 1360 0 1 1570
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1711307567
transform 1 0 1352 0 1 1570
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1711307567
transform 1 0 1344 0 1 1570
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1711307567
transform 1 0 1336 0 1 1570
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1711307567
transform 1 0 1304 0 1 1570
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1711307567
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1711307567
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1711307567
transform 1 0 1256 0 1 1570
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1711307567
transform 1 0 1248 0 1 1570
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1711307567
transform 1 0 1216 0 1 1570
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1711307567
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1711307567
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1711307567
transform 1 0 1160 0 1 1570
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1711307567
transform 1 0 1152 0 1 1570
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1711307567
transform 1 0 1144 0 1 1570
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1711307567
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1711307567
transform 1 0 1104 0 1 1570
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1711307567
transform 1 0 1096 0 1 1570
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1711307567
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1711307567
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1711307567
transform 1 0 1024 0 1 1570
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1711307567
transform 1 0 1016 0 1 1570
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1711307567
transform 1 0 1008 0 1 1570
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1711307567
transform 1 0 1000 0 1 1570
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1711307567
transform 1 0 992 0 1 1570
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1711307567
transform 1 0 944 0 1 1570
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1711307567
transform 1 0 936 0 1 1570
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1711307567
transform 1 0 928 0 1 1570
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1711307567
transform 1 0 920 0 1 1570
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1711307567
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1711307567
transform 1 0 888 0 1 1570
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1711307567
transform 1 0 856 0 1 1570
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1711307567
transform 1 0 848 0 1 1570
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1711307567
transform 1 0 816 0 1 1570
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1711307567
transform 1 0 808 0 1 1570
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1711307567
transform 1 0 800 0 1 1570
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1711307567
transform 1 0 792 0 1 1570
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1711307567
transform 1 0 760 0 1 1570
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1711307567
transform 1 0 752 0 1 1570
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1711307567
transform 1 0 728 0 1 1570
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1711307567
transform 1 0 688 0 1 1570
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1711307567
transform 1 0 680 0 1 1570
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1711307567
transform 1 0 672 0 1 1570
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1711307567
transform 1 0 664 0 1 1570
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1711307567
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1711307567
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1711307567
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1711307567
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1711307567
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1711307567
transform 1 0 544 0 1 1570
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1711307567
transform 1 0 536 0 1 1570
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1711307567
transform 1 0 496 0 1 1570
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1711307567
transform 1 0 488 0 1 1570
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1711307567
transform 1 0 480 0 1 1570
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1711307567
transform 1 0 432 0 1 1570
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1711307567
transform 1 0 424 0 1 1570
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1711307567
transform 1 0 416 0 1 1570
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1711307567
transform 1 0 408 0 1 1570
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1711307567
transform 1 0 400 0 1 1570
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1711307567
transform 1 0 344 0 1 1570
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1711307567
transform 1 0 336 0 1 1570
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1711307567
transform 1 0 328 0 1 1570
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1711307567
transform 1 0 320 0 1 1570
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1711307567
transform 1 0 312 0 1 1570
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1711307567
transform 1 0 280 0 1 1570
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1711307567
transform 1 0 272 0 1 1570
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1711307567
transform 1 0 232 0 1 1570
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1711307567
transform 1 0 224 0 1 1570
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1711307567
transform 1 0 216 0 1 1570
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1711307567
transform 1 0 208 0 1 1570
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1711307567
transform 1 0 200 0 1 1570
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1711307567
transform 1 0 192 0 1 1570
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1711307567
transform 1 0 184 0 1 1570
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1711307567
transform 1 0 176 0 1 1570
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1711307567
transform 1 0 168 0 1 1570
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1711307567
transform 1 0 160 0 1 1570
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1711307567
transform 1 0 152 0 1 1570
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1711307567
transform 1 0 144 0 1 1570
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1711307567
transform 1 0 136 0 1 1570
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1711307567
transform 1 0 128 0 1 1570
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1711307567
transform 1 0 120 0 1 1570
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1711307567
transform 1 0 112 0 1 1570
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1711307567
transform 1 0 104 0 1 1570
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1711307567
transform 1 0 96 0 1 1570
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1711307567
transform 1 0 88 0 1 1570
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1711307567
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1711307567
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1711307567
transform 1 0 2752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1711307567
transform 1 0 2744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1711307567
transform 1 0 2736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1711307567
transform 1 0 2728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1711307567
transform 1 0 2704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1711307567
transform 1 0 2696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1711307567
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1711307567
transform 1 0 2680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1711307567
transform 1 0 2672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1711307567
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1711307567
transform 1 0 2600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1711307567
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1711307567
transform 1 0 2584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1711307567
transform 1 0 2576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1711307567
transform 1 0 2568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1711307567
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1711307567
transform 1 0 2456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1711307567
transform 1 0 2448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1711307567
transform 1 0 2440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1711307567
transform 1 0 2432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1711307567
transform 1 0 2424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1711307567
transform 1 0 2416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1711307567
transform 1 0 2408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1711307567
transform 1 0 2400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1711307567
transform 1 0 2392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1711307567
transform 1 0 2384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1711307567
transform 1 0 2376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1711307567
transform 1 0 2368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1711307567
transform 1 0 2360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1711307567
transform 1 0 2352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1711307567
transform 1 0 2344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1711307567
transform 1 0 2336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1711307567
transform 1 0 2312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1711307567
transform 1 0 2304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1711307567
transform 1 0 2296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1711307567
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1711307567
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1711307567
transform 1 0 2256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1711307567
transform 1 0 2232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1711307567
transform 1 0 2224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1711307567
transform 1 0 2216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1711307567
transform 1 0 2208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1711307567
transform 1 0 2168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1711307567
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1711307567
transform 1 0 2152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1711307567
transform 1 0 2120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1711307567
transform 1 0 2112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1711307567
transform 1 0 2104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1711307567
transform 1 0 2040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1711307567
transform 1 0 2032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1711307567
transform 1 0 2024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1711307567
transform 1 0 2016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1711307567
transform 1 0 1952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1711307567
transform 1 0 1944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1711307567
transform 1 0 1936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1711307567
transform 1 0 1896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1711307567
transform 1 0 1888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1711307567
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1711307567
transform 1 0 1824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1711307567
transform 1 0 1816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1711307567
transform 1 0 1808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1711307567
transform 1 0 1800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1711307567
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1711307567
transform 1 0 1736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1711307567
transform 1 0 1728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1711307567
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1711307567
transform 1 0 1664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1711307567
transform 1 0 1656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1711307567
transform 1 0 1648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1711307567
transform 1 0 1600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1711307567
transform 1 0 1592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1711307567
transform 1 0 1584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1711307567
transform 1 0 1544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1711307567
transform 1 0 1504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1711307567
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1711307567
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1711307567
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1711307567
transform 1 0 1408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1711307567
transform 1 0 1400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1711307567
transform 1 0 1392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1711307567
transform 1 0 1352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1711307567
transform 1 0 1312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1711307567
transform 1 0 1304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1711307567
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1711307567
transform 1 0 1232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1711307567
transform 1 0 1224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1711307567
transform 1 0 1216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1711307567
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1711307567
transform 1 0 1168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1711307567
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1711307567
transform 1 0 1120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1711307567
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1711307567
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1711307567
transform 1 0 1056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1711307567
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1711307567
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1711307567
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1711307567
transform 1 0 984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1711307567
transform 1 0 976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1711307567
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1711307567
transform 1 0 944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1711307567
transform 1 0 936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1711307567
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1711307567
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1711307567
transform 1 0 872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1711307567
transform 1 0 864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1711307567
transform 1 0 824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1711307567
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1711307567
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1711307567
transform 1 0 768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1711307567
transform 1 0 736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1711307567
transform 1 0 728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1711307567
transform 1 0 720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1711307567
transform 1 0 680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1711307567
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1711307567
transform 1 0 640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1711307567
transform 1 0 608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1711307567
transform 1 0 600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1711307567
transform 1 0 592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1711307567
transform 1 0 544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1711307567
transform 1 0 536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1711307567
transform 1 0 528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1711307567
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1711307567
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1711307567
transform 1 0 456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1711307567
transform 1 0 448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1711307567
transform 1 0 408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1711307567
transform 1 0 400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1711307567
transform 1 0 392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1711307567
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1711307567
transform 1 0 352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1711307567
transform 1 0 344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1711307567
transform 1 0 312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1711307567
transform 1 0 304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1711307567
transform 1 0 296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1711307567
transform 1 0 288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1711307567
transform 1 0 280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1711307567
transform 1 0 240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1711307567
transform 1 0 232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1711307567
transform 1 0 224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1711307567
transform 1 0 216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1711307567
transform 1 0 112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1711307567
transform 1 0 104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1711307567
transform 1 0 96 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1711307567
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1711307567
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1711307567
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1711307567
transform 1 0 2024 0 1 1370
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1711307567
transform 1 0 2016 0 1 1370
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1711307567
transform 1 0 1952 0 1 1370
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1711307567
transform 1 0 1944 0 1 1370
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1711307567
transform 1 0 1936 0 1 1370
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1711307567
transform 1 0 1928 0 1 1370
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1711307567
transform 1 0 1920 0 1 1370
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1711307567
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1711307567
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1711307567
transform 1 0 1824 0 1 1370
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1711307567
transform 1 0 1816 0 1 1370
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1711307567
transform 1 0 1784 0 1 1370
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1711307567
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1711307567
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1711307567
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1711307567
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1711307567
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1711307567
transform 1 0 1672 0 1 1370
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1711307567
transform 1 0 1664 0 1 1370
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1711307567
transform 1 0 1592 0 1 1370
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1711307567
transform 1 0 1584 0 1 1370
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1711307567
transform 1 0 1576 0 1 1370
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1711307567
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1711307567
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1711307567
transform 1 0 1472 0 1 1370
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1711307567
transform 1 0 1440 0 1 1370
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1711307567
transform 1 0 1432 0 1 1370
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1711307567
transform 1 0 1424 0 1 1370
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1711307567
transform 1 0 1376 0 1 1370
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1711307567
transform 1 0 1368 0 1 1370
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1711307567
transform 1 0 1360 0 1 1370
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1711307567
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1711307567
transform 1 0 1304 0 1 1370
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1711307567
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1711307567
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1711307567
transform 1 0 1240 0 1 1370
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1711307567
transform 1 0 1232 0 1 1370
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1711307567
transform 1 0 1224 0 1 1370
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1711307567
transform 1 0 1216 0 1 1370
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1711307567
transform 1 0 1192 0 1 1370
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1711307567
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1711307567
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1711307567
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1711307567
transform 1 0 1120 0 1 1370
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1711307567
transform 1 0 1112 0 1 1370
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1711307567
transform 1 0 1104 0 1 1370
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1711307567
transform 1 0 1096 0 1 1370
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1711307567
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1711307567
transform 1 0 1032 0 1 1370
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1711307567
transform 1 0 1024 0 1 1370
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1711307567
transform 1 0 1016 0 1 1370
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1711307567
transform 1 0 1008 0 1 1370
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1711307567
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1711307567
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1711307567
transform 1 0 944 0 1 1370
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1711307567
transform 1 0 936 0 1 1370
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1711307567
transform 1 0 904 0 1 1370
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1711307567
transform 1 0 864 0 1 1370
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1711307567
transform 1 0 856 0 1 1370
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1711307567
transform 1 0 824 0 1 1370
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1711307567
transform 1 0 816 0 1 1370
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1711307567
transform 1 0 792 0 1 1370
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1711307567
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1711307567
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1711307567
transform 1 0 728 0 1 1370
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1711307567
transform 1 0 720 0 1 1370
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1711307567
transform 1 0 712 0 1 1370
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1711307567
transform 1 0 704 0 1 1370
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1711307567
transform 1 0 696 0 1 1370
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1711307567
transform 1 0 640 0 1 1370
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1711307567
transform 1 0 632 0 1 1370
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1711307567
transform 1 0 624 0 1 1370
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1711307567
transform 1 0 616 0 1 1370
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1711307567
transform 1 0 608 0 1 1370
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1711307567
transform 1 0 576 0 1 1370
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1711307567
transform 1 0 568 0 1 1370
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1711307567
transform 1 0 528 0 1 1370
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1711307567
transform 1 0 520 0 1 1370
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1711307567
transform 1 0 512 0 1 1370
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1711307567
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1711307567
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1711307567
transform 1 0 456 0 1 1370
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1711307567
transform 1 0 416 0 1 1370
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1711307567
transform 1 0 408 0 1 1370
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1711307567
transform 1 0 400 0 1 1370
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1711307567
transform 1 0 360 0 1 1370
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1711307567
transform 1 0 352 0 1 1370
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1711307567
transform 1 0 344 0 1 1370
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1711307567
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1711307567
transform 1 0 304 0 1 1370
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1711307567
transform 1 0 200 0 1 1370
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1711307567
transform 1 0 192 0 1 1370
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1711307567
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1711307567
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1711307567
transform 1 0 168 0 1 1370
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1711307567
transform 1 0 160 0 1 1370
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1711307567
transform 1 0 152 0 1 1370
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1711307567
transform 1 0 144 0 1 1370
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1711307567
transform 1 0 136 0 1 1370
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1711307567
transform 1 0 128 0 1 1370
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1711307567
transform 1 0 120 0 1 1370
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1711307567
transform 1 0 112 0 1 1370
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1711307567
transform 1 0 104 0 1 1370
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1711307567
transform 1 0 96 0 1 1370
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1711307567
transform 1 0 88 0 1 1370
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1711307567
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1711307567
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1711307567
transform 1 0 2752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1711307567
transform 1 0 2744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1711307567
transform 1 0 2736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1711307567
transform 1 0 2728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1711307567
transform 1 0 2720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1711307567
transform 1 0 2712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1711307567
transform 1 0 2704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1711307567
transform 1 0 2696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1711307567
transform 1 0 2592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1711307567
transform 1 0 2584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1711307567
transform 1 0 2576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1711307567
transform 1 0 2568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1711307567
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1711307567
transform 1 0 2552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1711307567
transform 1 0 2504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1711307567
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1711307567
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1711307567
transform 1 0 2464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1711307567
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1711307567
transform 1 0 2448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1711307567
transform 1 0 2440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1711307567
transform 1 0 2432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1711307567
transform 1 0 2424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1711307567
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1711307567
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1711307567
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1711307567
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1711307567
transform 1 0 2344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1711307567
transform 1 0 2320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1711307567
transform 1 0 2312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1711307567
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1711307567
transform 1 0 2296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1711307567
transform 1 0 2288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1711307567
transform 1 0 2280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1711307567
transform 1 0 2176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1711307567
transform 1 0 2168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1711307567
transform 1 0 2160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1711307567
transform 1 0 2152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1711307567
transform 1 0 2144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1711307567
transform 1 0 2136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1711307567
transform 1 0 2128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1711307567
transform 1 0 2120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1711307567
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1711307567
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1711307567
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1711307567
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1711307567
transform 1 0 2064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1711307567
transform 1 0 2056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1711307567
transform 1 0 2048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1711307567
transform 1 0 2040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1711307567
transform 1 0 2016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1711307567
transform 1 0 2008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1711307567
transform 1 0 2000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1711307567
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1711307567
transform 1 0 1952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1711307567
transform 1 0 1944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1711307567
transform 1 0 1904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1711307567
transform 1 0 1896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1711307567
transform 1 0 1864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1711307567
transform 1 0 1856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1711307567
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1711307567
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1711307567
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1711307567
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1711307567
transform 1 0 1752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1711307567
transform 1 0 1744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1711307567
transform 1 0 1736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1711307567
transform 1 0 1728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1711307567
transform 1 0 1664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1711307567
transform 1 0 1656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1711307567
transform 1 0 1616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1711307567
transform 1 0 1576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1711307567
transform 1 0 1568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1711307567
transform 1 0 1560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1711307567
transform 1 0 1552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1711307567
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1711307567
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1711307567
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1711307567
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1711307567
transform 1 0 1432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1711307567
transform 1 0 1384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1711307567
transform 1 0 1376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1711307567
transform 1 0 1368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1711307567
transform 1 0 1360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1711307567
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1711307567
transform 1 0 1280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1711307567
transform 1 0 1272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1711307567
transform 1 0 1264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1711307567
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1711307567
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1711307567
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1711307567
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1711307567
transform 1 0 1160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1711307567
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1711307567
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1711307567
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1711307567
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1711307567
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1711307567
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1711307567
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1711307567
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1711307567
transform 1 0 1000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1711307567
transform 1 0 960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1711307567
transform 1 0 952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1711307567
transform 1 0 944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1711307567
transform 1 0 936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1711307567
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1711307567
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1711307567
transform 1 0 880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1711307567
transform 1 0 872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1711307567
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1711307567
transform 1 0 840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1711307567
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1711307567
transform 1 0 824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1711307567
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1711307567
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1711307567
transform 1 0 768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1711307567
transform 1 0 760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1711307567
transform 1 0 752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1711307567
transform 1 0 744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1711307567
transform 1 0 720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1711307567
transform 1 0 680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1711307567
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1711307567
transform 1 0 664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1711307567
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1711307567
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1711307567
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1711307567
transform 1 0 608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1711307567
transform 1 0 600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1711307567
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1711307567
transform 1 0 560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1711307567
transform 1 0 552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1711307567
transform 1 0 544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1711307567
transform 1 0 536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1711307567
transform 1 0 528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1711307567
transform 1 0 496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1711307567
transform 1 0 488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1711307567
transform 1 0 480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1711307567
transform 1 0 440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1711307567
transform 1 0 432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1711307567
transform 1 0 424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1711307567
transform 1 0 416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1711307567
transform 1 0 408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1711307567
transform 1 0 400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1711307567
transform 1 0 392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1711307567
transform 1 0 288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1711307567
transform 1 0 280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1711307567
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1711307567
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1711307567
transform 1 0 256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1711307567
transform 1 0 248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1711307567
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1711307567
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1711307567
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1711307567
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1711307567
transform 1 0 168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1711307567
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1711307567
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1711307567
transform 1 0 104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1711307567
transform 1 0 96 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1711307567
transform 1 0 88 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1711307567
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1711307567
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1711307567
transform 1 0 2656 0 1 1170
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1711307567
transform 1 0 2648 0 1 1170
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1711307567
transform 1 0 2640 0 1 1170
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1711307567
transform 1 0 2440 0 1 1170
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1711307567
transform 1 0 2432 0 1 1170
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1711307567
transform 1 0 2424 0 1 1170
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1711307567
transform 1 0 2376 0 1 1170
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1711307567
transform 1 0 2368 0 1 1170
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1711307567
transform 1 0 2360 0 1 1170
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1711307567
transform 1 0 2352 0 1 1170
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1711307567
transform 1 0 2304 0 1 1170
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1711307567
transform 1 0 2264 0 1 1170
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1711307567
transform 1 0 2256 0 1 1170
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1711307567
transform 1 0 2248 0 1 1170
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1711307567
transform 1 0 2240 0 1 1170
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1711307567
transform 1 0 2232 0 1 1170
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1711307567
transform 1 0 2224 0 1 1170
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1711307567
transform 1 0 2176 0 1 1170
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1711307567
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1711307567
transform 1 0 1968 0 1 1170
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1711307567
transform 1 0 1920 0 1 1170
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1711307567
transform 1 0 1912 0 1 1170
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1711307567
transform 1 0 1904 0 1 1170
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1711307567
transform 1 0 1800 0 1 1170
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1711307567
transform 1 0 1600 0 1 1170
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1711307567
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1711307567
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1711307567
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1711307567
transform 1 0 1480 0 1 1170
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1711307567
transform 1 0 1448 0 1 1170
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1711307567
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1711307567
transform 1 0 1400 0 1 1170
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1711307567
transform 1 0 1392 0 1 1170
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1711307567
transform 1 0 1384 0 1 1170
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1711307567
transform 1 0 1328 0 1 1170
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1711307567
transform 1 0 1320 0 1 1170
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1711307567
transform 1 0 1312 0 1 1170
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1711307567
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1711307567
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1711307567
transform 1 0 1240 0 1 1170
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1711307567
transform 1 0 1232 0 1 1170
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1711307567
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1711307567
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1711307567
transform 1 0 1144 0 1 1170
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1711307567
transform 1 0 1136 0 1 1170
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1711307567
transform 1 0 1080 0 1 1170
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1711307567
transform 1 0 1072 0 1 1170
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1711307567
transform 1 0 1064 0 1 1170
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1711307567
transform 1 0 1056 0 1 1170
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1711307567
transform 1 0 1048 0 1 1170
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1711307567
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1711307567
transform 1 0 1000 0 1 1170
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1711307567
transform 1 0 992 0 1 1170
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1711307567
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1711307567
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1711307567
transform 1 0 888 0 1 1170
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1711307567
transform 1 0 880 0 1 1170
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1711307567
transform 1 0 872 0 1 1170
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1711307567
transform 1 0 808 0 1 1170
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1711307567
transform 1 0 800 0 1 1170
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1711307567
transform 1 0 792 0 1 1170
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1711307567
transform 1 0 784 0 1 1170
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1711307567
transform 1 0 728 0 1 1170
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1711307567
transform 1 0 720 0 1 1170
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1711307567
transform 1 0 712 0 1 1170
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1711307567
transform 1 0 680 0 1 1170
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1711307567
transform 1 0 576 0 1 1170
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1711307567
transform 1 0 568 0 1 1170
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1711307567
transform 1 0 464 0 1 1170
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1711307567
transform 1 0 360 0 1 1170
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1711307567
transform 1 0 352 0 1 1170
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1711307567
transform 1 0 344 0 1 1170
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1711307567
transform 1 0 336 0 1 1170
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1711307567
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1711307567
transform 1 0 280 0 1 1170
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1711307567
transform 1 0 272 0 1 1170
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1711307567
transform 1 0 264 0 1 1170
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1711307567
transform 1 0 256 0 1 1170
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1711307567
transform 1 0 248 0 1 1170
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1711307567
transform 1 0 200 0 1 1170
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1711307567
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1711307567
transform 1 0 184 0 1 1170
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1711307567
transform 1 0 176 0 1 1170
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1711307567
transform 1 0 168 0 1 1170
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1711307567
transform 1 0 2752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1711307567
transform 1 0 2744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1711307567
transform 1 0 2736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1711307567
transform 1 0 2728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1711307567
transform 1 0 2720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1711307567
transform 1 0 2712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1711307567
transform 1 0 2704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1711307567
transform 1 0 2696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1711307567
transform 1 0 2688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1711307567
transform 1 0 2680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1711307567
transform 1 0 2624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1711307567
transform 1 0 2616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1711307567
transform 1 0 2608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1711307567
transform 1 0 2600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1711307567
transform 1 0 2568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1711307567
transform 1 0 2560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1711307567
transform 1 0 2552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1711307567
transform 1 0 2544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1711307567
transform 1 0 2536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1711307567
transform 1 0 2528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1711307567
transform 1 0 2520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1711307567
transform 1 0 2512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1711307567
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1711307567
transform 1 0 2472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1711307567
transform 1 0 2464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1711307567
transform 1 0 2456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1711307567
transform 1 0 2448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1711307567
transform 1 0 2344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1711307567
transform 1 0 2336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1711307567
transform 1 0 2328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1711307567
transform 1 0 2320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1711307567
transform 1 0 2312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1711307567
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1711307567
transform 1 0 2296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1711307567
transform 1 0 2288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1711307567
transform 1 0 2184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1711307567
transform 1 0 2176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1711307567
transform 1 0 2168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1711307567
transform 1 0 2144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1711307567
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1711307567
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1711307567
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1711307567
transform 1 0 2072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1711307567
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1711307567
transform 1 0 2056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1711307567
transform 1 0 2048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1711307567
transform 1 0 2040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1711307567
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1711307567
transform 1 0 1976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1711307567
transform 1 0 1952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1711307567
transform 1 0 1896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1711307567
transform 1 0 1888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1711307567
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1711307567
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1711307567
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1711307567
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1711307567
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1711307567
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1711307567
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1711307567
transform 1 0 1736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1711307567
transform 1 0 1728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1711307567
transform 1 0 1720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1711307567
transform 1 0 1712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1711307567
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1711307567
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1711307567
transform 1 0 1688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1711307567
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1711307567
transform 1 0 1672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1711307567
transform 1 0 1664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1711307567
transform 1 0 1656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1711307567
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1711307567
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1711307567
transform 1 0 1632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1711307567
transform 1 0 1624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1711307567
transform 1 0 1616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1711307567
transform 1 0 1584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1711307567
transform 1 0 1576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1711307567
transform 1 0 1544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1711307567
transform 1 0 1536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1711307567
transform 1 0 1528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1711307567
transform 1 0 1520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1711307567
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1711307567
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1711307567
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1711307567
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1711307567
transform 1 0 1392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1711307567
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1711307567
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1711307567
transform 1 0 1320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1711307567
transform 1 0 1312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1711307567
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1711307567
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1711307567
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1711307567
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1711307567
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1711307567
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1711307567
transform 1 0 1136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1711307567
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1711307567
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1711307567
transform 1 0 1112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1711307567
transform 1 0 1104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1711307567
transform 1 0 1000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1711307567
transform 1 0 992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1711307567
transform 1 0 984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1711307567
transform 1 0 952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1711307567
transform 1 0 944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1711307567
transform 1 0 936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1711307567
transform 1 0 832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1711307567
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1711307567
transform 1 0 816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1711307567
transform 1 0 808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1711307567
transform 1 0 776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1711307567
transform 1 0 768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1711307567
transform 1 0 760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1711307567
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1711307567
transform 1 0 648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1711307567
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1711307567
transform 1 0 632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1711307567
transform 1 0 624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1711307567
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1711307567
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1711307567
transform 1 0 560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1711307567
transform 1 0 536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1711307567
transform 1 0 528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1711307567
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1711307567
transform 1 0 512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1711307567
transform 1 0 504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1711307567
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1711307567
transform 1 0 448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1711307567
transform 1 0 440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1711307567
transform 1 0 432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1711307567
transform 1 0 424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1711307567
transform 1 0 416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1711307567
transform 1 0 408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1711307567
transform 1 0 400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1711307567
transform 1 0 392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1711307567
transform 1 0 336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1711307567
transform 1 0 328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1711307567
transform 1 0 320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1711307567
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1711307567
transform 1 0 304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1711307567
transform 1 0 256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1711307567
transform 1 0 248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1711307567
transform 1 0 240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1711307567
transform 1 0 232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1711307567
transform 1 0 224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1711307567
transform 1 0 120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1711307567
transform 1 0 112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1711307567
transform 1 0 104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1711307567
transform 1 0 96 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1711307567
transform 1 0 88 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1711307567
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1711307567
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1711307567
transform 1 0 2752 0 1 970
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1711307567
transform 1 0 2744 0 1 970
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1711307567
transform 1 0 2736 0 1 970
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1711307567
transform 1 0 2728 0 1 970
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1711307567
transform 1 0 2720 0 1 970
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1711307567
transform 1 0 2712 0 1 970
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1711307567
transform 1 0 2704 0 1 970
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1711307567
transform 1 0 2696 0 1 970
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1711307567
transform 1 0 2688 0 1 970
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1711307567
transform 1 0 2680 0 1 970
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1711307567
transform 1 0 2672 0 1 970
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1711307567
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1711307567
transform 1 0 2656 0 1 970
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1711307567
transform 1 0 2648 0 1 970
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1711307567
transform 1 0 2640 0 1 970
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1711307567
transform 1 0 2632 0 1 970
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1711307567
transform 1 0 2624 0 1 970
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1711307567
transform 1 0 2616 0 1 970
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1711307567
transform 1 0 2592 0 1 970
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1711307567
transform 1 0 2584 0 1 970
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1711307567
transform 1 0 2576 0 1 970
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1711307567
transform 1 0 2552 0 1 970
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1711307567
transform 1 0 2544 0 1 970
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1711307567
transform 1 0 2536 0 1 970
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1711307567
transform 1 0 2528 0 1 970
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1711307567
transform 1 0 2504 0 1 970
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1711307567
transform 1 0 2496 0 1 970
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1711307567
transform 1 0 2488 0 1 970
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1711307567
transform 1 0 2456 0 1 970
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1711307567
transform 1 0 2448 0 1 970
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1711307567
transform 1 0 2440 0 1 970
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1711307567
transform 1 0 2432 0 1 970
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1711307567
transform 1 0 2424 0 1 970
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1711307567
transform 1 0 2416 0 1 970
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1711307567
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1711307567
transform 1 0 2400 0 1 970
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1711307567
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1711307567
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1711307567
transform 1 0 2376 0 1 970
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1711307567
transform 1 0 2368 0 1 970
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1711307567
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1711307567
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1711307567
transform 1 0 2328 0 1 970
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1711307567
transform 1 0 2296 0 1 970
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1711307567
transform 1 0 2288 0 1 970
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1711307567
transform 1 0 2256 0 1 970
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1711307567
transform 1 0 2248 0 1 970
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1711307567
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1711307567
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1711307567
transform 1 0 2224 0 1 970
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1711307567
transform 1 0 2216 0 1 970
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1711307567
transform 1 0 2208 0 1 970
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1711307567
transform 1 0 2104 0 1 970
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1711307567
transform 1 0 2096 0 1 970
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1711307567
transform 1 0 2088 0 1 970
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1711307567
transform 1 0 2064 0 1 970
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1711307567
transform 1 0 2056 0 1 970
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1711307567
transform 1 0 2024 0 1 970
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1711307567
transform 1 0 2016 0 1 970
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1711307567
transform 1 0 2008 0 1 970
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1711307567
transform 1 0 1984 0 1 970
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1711307567
transform 1 0 1976 0 1 970
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1711307567
transform 1 0 1968 0 1 970
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1711307567
transform 1 0 1960 0 1 970
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1711307567
transform 1 0 1952 0 1 970
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1711307567
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1711307567
transform 1 0 1920 0 1 970
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1711307567
transform 1 0 1912 0 1 970
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1711307567
transform 1 0 1904 0 1 970
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1711307567
transform 1 0 1896 0 1 970
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1711307567
transform 1 0 1888 0 1 970
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1711307567
transform 1 0 1840 0 1 970
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1711307567
transform 1 0 1832 0 1 970
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1711307567
transform 1 0 1824 0 1 970
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1711307567
transform 1 0 1816 0 1 970
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1711307567
transform 1 0 1808 0 1 970
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1711307567
transform 1 0 1800 0 1 970
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1711307567
transform 1 0 1792 0 1 970
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1711307567
transform 1 0 1592 0 1 970
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1711307567
transform 1 0 1488 0 1 970
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1711307567
transform 1 0 1480 0 1 970
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1711307567
transform 1 0 1448 0 1 970
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1711307567
transform 1 0 1440 0 1 970
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1711307567
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1711307567
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1711307567
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1711307567
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1711307567
transform 1 0 1304 0 1 970
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1711307567
transform 1 0 1296 0 1 970
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1711307567
transform 1 0 1288 0 1 970
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1711307567
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1711307567
transform 1 0 1272 0 1 970
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1711307567
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1711307567
transform 1 0 1256 0 1 970
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1711307567
transform 1 0 1248 0 1 970
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1711307567
transform 1 0 1240 0 1 970
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1711307567
transform 1 0 1040 0 1 970
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1711307567
transform 1 0 1032 0 1 970
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1711307567
transform 1 0 1024 0 1 970
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1711307567
transform 1 0 920 0 1 970
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1711307567
transform 1 0 912 0 1 970
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1711307567
transform 1 0 904 0 1 970
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1711307567
transform 1 0 896 0 1 970
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1711307567
transform 1 0 888 0 1 970
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1711307567
transform 1 0 880 0 1 970
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1711307567
transform 1 0 872 0 1 970
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1711307567
transform 1 0 864 0 1 970
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1711307567
transform 1 0 856 0 1 970
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1711307567
transform 1 0 848 0 1 970
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1711307567
transform 1 0 744 0 1 970
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1711307567
transform 1 0 736 0 1 970
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1711307567
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1711307567
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1711307567
transform 1 0 712 0 1 970
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1711307567
transform 1 0 704 0 1 970
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1711307567
transform 1 0 696 0 1 970
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1711307567
transform 1 0 648 0 1 970
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1711307567
transform 1 0 640 0 1 970
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1711307567
transform 1 0 632 0 1 970
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1711307567
transform 1 0 608 0 1 970
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1711307567
transform 1 0 600 0 1 970
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1711307567
transform 1 0 592 0 1 970
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1711307567
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1711307567
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1711307567
transform 1 0 568 0 1 970
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1711307567
transform 1 0 520 0 1 970
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1711307567
transform 1 0 512 0 1 970
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1711307567
transform 1 0 504 0 1 970
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1711307567
transform 1 0 496 0 1 970
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1711307567
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1711307567
transform 1 0 480 0 1 970
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1711307567
transform 1 0 432 0 1 970
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1711307567
transform 1 0 424 0 1 970
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1711307567
transform 1 0 416 0 1 970
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1711307567
transform 1 0 408 0 1 970
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1711307567
transform 1 0 400 0 1 970
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1711307567
transform 1 0 392 0 1 970
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1711307567
transform 1 0 384 0 1 970
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1711307567
transform 1 0 344 0 1 970
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1711307567
transform 1 0 336 0 1 970
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1711307567
transform 1 0 328 0 1 970
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1711307567
transform 1 0 320 0 1 970
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1711307567
transform 1 0 312 0 1 970
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1711307567
transform 1 0 304 0 1 970
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1711307567
transform 1 0 296 0 1 970
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1711307567
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1711307567
transform 1 0 248 0 1 970
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1711307567
transform 1 0 240 0 1 970
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1711307567
transform 1 0 232 0 1 970
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1711307567
transform 1 0 224 0 1 970
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1711307567
transform 1 0 192 0 1 970
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1711307567
transform 1 0 184 0 1 970
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1711307567
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1711307567
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1711307567
transform 1 0 160 0 1 970
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1711307567
transform 1 0 152 0 1 970
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1711307567
transform 1 0 144 0 1 970
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1711307567
transform 1 0 136 0 1 970
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1711307567
transform 1 0 128 0 1 970
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1711307567
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1711307567
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1711307567
transform 1 0 2656 0 -1 970
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1711307567
transform 1 0 2584 0 -1 970
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1711307567
transform 1 0 2448 0 -1 970
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1711307567
transform 1 0 2440 0 -1 970
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1711307567
transform 1 0 2336 0 -1 970
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1711307567
transform 1 0 2328 0 -1 970
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1711307567
transform 1 0 2320 0 -1 970
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1711307567
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1711307567
transform 1 0 2256 0 -1 970
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1711307567
transform 1 0 2248 0 -1 970
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1711307567
transform 1 0 2240 0 -1 970
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1711307567
transform 1 0 2184 0 -1 970
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1711307567
transform 1 0 2176 0 -1 970
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1711307567
transform 1 0 2168 0 -1 970
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1711307567
transform 1 0 2160 0 -1 970
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1711307567
transform 1 0 2112 0 -1 970
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1711307567
transform 1 0 2104 0 -1 970
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1711307567
transform 1 0 2096 0 -1 970
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1711307567
transform 1 0 2088 0 -1 970
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1711307567
transform 1 0 2056 0 -1 970
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1711307567
transform 1 0 2048 0 -1 970
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1711307567
transform 1 0 2040 0 -1 970
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1711307567
transform 1 0 1992 0 -1 970
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1711307567
transform 1 0 1984 0 -1 970
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1711307567
transform 1 0 1880 0 -1 970
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1711307567
transform 1 0 1872 0 -1 970
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1711307567
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1711307567
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1711307567
transform 1 0 1752 0 -1 970
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1711307567
transform 1 0 1744 0 -1 970
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1711307567
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1711307567
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1711307567
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1711307567
transform 1 0 1648 0 -1 970
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1711307567
transform 1 0 1640 0 -1 970
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1711307567
transform 1 0 1632 0 -1 970
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1711307567
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1711307567
transform 1 0 1576 0 -1 970
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1711307567
transform 1 0 1568 0 -1 970
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1711307567
transform 1 0 1536 0 -1 970
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1711307567
transform 1 0 1528 0 -1 970
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1711307567
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1711307567
transform 1 0 1416 0 -1 970
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1711307567
transform 1 0 1408 0 -1 970
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1711307567
transform 1 0 1400 0 -1 970
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1711307567
transform 1 0 1296 0 -1 970
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1711307567
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1711307567
transform 1 0 1224 0 -1 970
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1711307567
transform 1 0 1216 0 -1 970
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1711307567
transform 1 0 1208 0 -1 970
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1711307567
transform 1 0 1200 0 -1 970
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1711307567
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1711307567
transform 1 0 1168 0 -1 970
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1711307567
transform 1 0 1120 0 -1 970
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1711307567
transform 1 0 1112 0 -1 970
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1711307567
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1711307567
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1711307567
transform 1 0 1088 0 -1 970
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1711307567
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1711307567
transform 1 0 1032 0 -1 970
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1711307567
transform 1 0 1024 0 -1 970
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1711307567
transform 1 0 1016 0 -1 970
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1711307567
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1711307567
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1711307567
transform 1 0 952 0 -1 970
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1711307567
transform 1 0 944 0 -1 970
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1711307567
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1711307567
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1711307567
transform 1 0 848 0 -1 970
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1711307567
transform 1 0 840 0 -1 970
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1711307567
transform 1 0 832 0 -1 970
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1711307567
transform 1 0 760 0 -1 970
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1711307567
transform 1 0 752 0 -1 970
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1711307567
transform 1 0 744 0 -1 970
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1711307567
transform 1 0 736 0 -1 970
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1711307567
transform 1 0 728 0 -1 970
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1711307567
transform 1 0 664 0 -1 970
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1711307567
transform 1 0 656 0 -1 970
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1711307567
transform 1 0 648 0 -1 970
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1711307567
transform 1 0 640 0 -1 970
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1711307567
transform 1 0 584 0 -1 970
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1711307567
transform 1 0 576 0 -1 970
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1711307567
transform 1 0 568 0 -1 970
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1711307567
transform 1 0 520 0 -1 970
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1711307567
transform 1 0 512 0 -1 970
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1711307567
transform 1 0 504 0 -1 970
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1711307567
transform 1 0 496 0 -1 970
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1711307567
transform 1 0 488 0 -1 970
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1711307567
transform 1 0 424 0 -1 970
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1711307567
transform 1 0 416 0 -1 970
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1711307567
transform 1 0 408 0 -1 970
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1711307567
transform 1 0 400 0 -1 970
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1711307567
transform 1 0 344 0 -1 970
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1711307567
transform 1 0 336 0 -1 970
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1711307567
transform 1 0 328 0 -1 970
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1711307567
transform 1 0 320 0 -1 970
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1711307567
transform 1 0 280 0 -1 970
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1711307567
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1711307567
transform 1 0 240 0 -1 970
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1711307567
transform 1 0 232 0 -1 970
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1711307567
transform 1 0 224 0 -1 970
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1711307567
transform 1 0 184 0 -1 970
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1711307567
transform 1 0 176 0 -1 970
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1711307567
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1711307567
transform 1 0 2656 0 1 770
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1711307567
transform 1 0 2648 0 1 770
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1711307567
transform 1 0 2640 0 1 770
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1711307567
transform 1 0 2584 0 1 770
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1711307567
transform 1 0 2576 0 1 770
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1711307567
transform 1 0 2568 0 1 770
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1711307567
transform 1 0 2560 0 1 770
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1711307567
transform 1 0 2512 0 1 770
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1711307567
transform 1 0 2504 0 1 770
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1711307567
transform 1 0 2496 0 1 770
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1711307567
transform 1 0 2456 0 1 770
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1711307567
transform 1 0 2432 0 1 770
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1711307567
transform 1 0 2424 0 1 770
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1711307567
transform 1 0 2416 0 1 770
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1711307567
transform 1 0 2408 0 1 770
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1711307567
transform 1 0 2376 0 1 770
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1711307567
transform 1 0 2368 0 1 770
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1711307567
transform 1 0 2336 0 1 770
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1711307567
transform 1 0 2328 0 1 770
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1711307567
transform 1 0 2304 0 1 770
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1711307567
transform 1 0 2296 0 1 770
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1711307567
transform 1 0 2256 0 1 770
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1711307567
transform 1 0 2248 0 1 770
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1711307567
transform 1 0 2216 0 1 770
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1711307567
transform 1 0 2208 0 1 770
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1711307567
transform 1 0 2176 0 1 770
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1711307567
transform 1 0 2152 0 1 770
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1711307567
transform 1 0 2144 0 1 770
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1711307567
transform 1 0 2136 0 1 770
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1711307567
transform 1 0 2128 0 1 770
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1711307567
transform 1 0 2120 0 1 770
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1711307567
transform 1 0 2064 0 1 770
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1711307567
transform 1 0 1960 0 1 770
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1711307567
transform 1 0 1952 0 1 770
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1711307567
transform 1 0 1944 0 1 770
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1711307567
transform 1 0 1872 0 1 770
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1711307567
transform 1 0 1864 0 1 770
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1711307567
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1711307567
transform 1 0 1752 0 1 770
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1711307567
transform 1 0 1688 0 1 770
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1711307567
transform 1 0 1680 0 1 770
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1711307567
transform 1 0 1672 0 1 770
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1711307567
transform 1 0 1664 0 1 770
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1711307567
transform 1 0 1656 0 1 770
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1711307567
transform 1 0 1592 0 1 770
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1711307567
transform 1 0 1584 0 1 770
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1711307567
transform 1 0 1576 0 1 770
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1711307567
transform 1 0 1568 0 1 770
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1711307567
transform 1 0 1496 0 1 770
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1711307567
transform 1 0 1488 0 1 770
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1711307567
transform 1 0 1480 0 1 770
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1711307567
transform 1 0 1472 0 1 770
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1711307567
transform 1 0 1464 0 1 770
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1711307567
transform 1 0 1416 0 1 770
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1711307567
transform 1 0 1408 0 1 770
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1711307567
transform 1 0 1360 0 1 770
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1711307567
transform 1 0 1352 0 1 770
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1711307567
transform 1 0 1344 0 1 770
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1711307567
transform 1 0 1336 0 1 770
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1711307567
transform 1 0 1296 0 1 770
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1711307567
transform 1 0 1288 0 1 770
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1711307567
transform 1 0 1280 0 1 770
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1711307567
transform 1 0 1232 0 1 770
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1711307567
transform 1 0 1224 0 1 770
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1711307567
transform 1 0 1216 0 1 770
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1711307567
transform 1 0 1208 0 1 770
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1711307567
transform 1 0 1176 0 1 770
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1711307567
transform 1 0 1136 0 1 770
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1711307567
transform 1 0 1128 0 1 770
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1711307567
transform 1 0 1120 0 1 770
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1711307567
transform 1 0 1080 0 1 770
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1711307567
transform 1 0 1072 0 1 770
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1711307567
transform 1 0 1032 0 1 770
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1711307567
transform 1 0 1024 0 1 770
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1711307567
transform 1 0 984 0 1 770
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1711307567
transform 1 0 976 0 1 770
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1711307567
transform 1 0 968 0 1 770
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1711307567
transform 1 0 944 0 1 770
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1711307567
transform 1 0 936 0 1 770
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1711307567
transform 1 0 904 0 1 770
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1711307567
transform 1 0 896 0 1 770
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1711307567
transform 1 0 856 0 1 770
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1711307567
transform 1 0 848 0 1 770
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1711307567
transform 1 0 808 0 1 770
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1711307567
transform 1 0 800 0 1 770
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1711307567
transform 1 0 792 0 1 770
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1711307567
transform 1 0 736 0 1 770
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1711307567
transform 1 0 728 0 1 770
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1711307567
transform 1 0 720 0 1 770
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1711307567
transform 1 0 712 0 1 770
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1711307567
transform 1 0 704 0 1 770
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1711307567
transform 1 0 696 0 1 770
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1711307567
transform 1 0 656 0 1 770
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1711307567
transform 1 0 632 0 1 770
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1711307567
transform 1 0 624 0 1 770
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1711307567
transform 1 0 600 0 1 770
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1711307567
transform 1 0 592 0 1 770
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1711307567
transform 1 0 584 0 1 770
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1711307567
transform 1 0 576 0 1 770
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1711307567
transform 1 0 536 0 1 770
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1711307567
transform 1 0 528 0 1 770
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1711307567
transform 1 0 520 0 1 770
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1711307567
transform 1 0 512 0 1 770
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1711307567
transform 1 0 480 0 1 770
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1711307567
transform 1 0 472 0 1 770
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1711307567
transform 1 0 448 0 1 770
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1711307567
transform 1 0 440 0 1 770
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1711307567
transform 1 0 432 0 1 770
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1711307567
transform 1 0 424 0 1 770
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1711307567
transform 1 0 416 0 1 770
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1711307567
transform 1 0 368 0 1 770
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1711307567
transform 1 0 360 0 1 770
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1711307567
transform 1 0 352 0 1 770
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1711307567
transform 1 0 344 0 1 770
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1711307567
transform 1 0 336 0 1 770
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1711307567
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1711307567
transform 1 0 320 0 1 770
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1711307567
transform 1 0 288 0 1 770
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1711307567
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1711307567
transform 1 0 272 0 1 770
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1711307567
transform 1 0 264 0 1 770
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1711307567
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1711307567
transform 1 0 216 0 1 770
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1711307567
transform 1 0 208 0 1 770
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1711307567
transform 1 0 184 0 1 770
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1711307567
transform 1 0 176 0 1 770
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1711307567
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1711307567
transform 1 0 2656 0 -1 770
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1711307567
transform 1 0 2648 0 -1 770
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1711307567
transform 1 0 2592 0 -1 770
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1711307567
transform 1 0 2584 0 -1 770
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1711307567
transform 1 0 2560 0 -1 770
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1711307567
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1711307567
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1711307567
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1711307567
transform 1 0 2488 0 -1 770
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1711307567
transform 1 0 2424 0 -1 770
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1711307567
transform 1 0 2416 0 -1 770
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1711307567
transform 1 0 2408 0 -1 770
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1711307567
transform 1 0 2400 0 -1 770
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1711307567
transform 1 0 2392 0 -1 770
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1711307567
transform 1 0 2360 0 -1 770
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1711307567
transform 1 0 2328 0 -1 770
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1711307567
transform 1 0 2320 0 -1 770
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1711307567
transform 1 0 2312 0 -1 770
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1711307567
transform 1 0 2304 0 -1 770
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1711307567
transform 1 0 2272 0 -1 770
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1711307567
transform 1 0 2264 0 -1 770
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1711307567
transform 1 0 2256 0 -1 770
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1711307567
transform 1 0 2248 0 -1 770
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1711307567
transform 1 0 2200 0 -1 770
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1711307567
transform 1 0 2192 0 -1 770
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1711307567
transform 1 0 2184 0 -1 770
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1711307567
transform 1 0 2176 0 -1 770
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1711307567
transform 1 0 2136 0 -1 770
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1711307567
transform 1 0 2096 0 -1 770
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1711307567
transform 1 0 2088 0 -1 770
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1711307567
transform 1 0 2080 0 -1 770
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1711307567
transform 1 0 2032 0 -1 770
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1711307567
transform 1 0 2024 0 -1 770
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1711307567
transform 1 0 2016 0 -1 770
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1711307567
transform 1 0 2008 0 -1 770
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1711307567
transform 1 0 1984 0 -1 770
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1711307567
transform 1 0 1952 0 -1 770
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1711307567
transform 1 0 1928 0 -1 770
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1711307567
transform 1 0 1920 0 -1 770
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1711307567
transform 1 0 1912 0 -1 770
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1711307567
transform 1 0 1880 0 -1 770
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1711307567
transform 1 0 1840 0 -1 770
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1711307567
transform 1 0 1832 0 -1 770
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1711307567
transform 1 0 1824 0 -1 770
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1711307567
transform 1 0 1776 0 -1 770
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1711307567
transform 1 0 1768 0 -1 770
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1711307567
transform 1 0 1760 0 -1 770
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1711307567
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1711307567
transform 1 0 1696 0 -1 770
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1711307567
transform 1 0 1688 0 -1 770
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1711307567
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1711307567
transform 1 0 1624 0 -1 770
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1711307567
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1711307567
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1711307567
transform 1 0 1576 0 -1 770
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1711307567
transform 1 0 1536 0 -1 770
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1711307567
transform 1 0 1528 0 -1 770
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1711307567
transform 1 0 1520 0 -1 770
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1711307567
transform 1 0 1512 0 -1 770
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1711307567
transform 1 0 1472 0 -1 770
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1711307567
transform 1 0 1464 0 -1 770
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1711307567
transform 1 0 1456 0 -1 770
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1711307567
transform 1 0 1424 0 -1 770
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1711307567
transform 1 0 1416 0 -1 770
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1711307567
transform 1 0 1408 0 -1 770
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1711307567
transform 1 0 1360 0 -1 770
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1711307567
transform 1 0 1352 0 -1 770
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1711307567
transform 1 0 1344 0 -1 770
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1711307567
transform 1 0 1336 0 -1 770
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1711307567
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1711307567
transform 1 0 1280 0 -1 770
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1711307567
transform 1 0 1272 0 -1 770
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1711307567
transform 1 0 1264 0 -1 770
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1711307567
transform 1 0 1240 0 -1 770
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1711307567
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1711307567
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1711307567
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1711307567
transform 1 0 1152 0 -1 770
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1711307567
transform 1 0 1144 0 -1 770
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1711307567
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1711307567
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1711307567
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1711307567
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1711307567
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1711307567
transform 1 0 1040 0 -1 770
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1711307567
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1711307567
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1711307567
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1711307567
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1711307567
transform 1 0 968 0 -1 770
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1711307567
transform 1 0 960 0 -1 770
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1711307567
transform 1 0 952 0 -1 770
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1711307567
transform 1 0 912 0 -1 770
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1711307567
transform 1 0 904 0 -1 770
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1711307567
transform 1 0 896 0 -1 770
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1711307567
transform 1 0 888 0 -1 770
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1711307567
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1711307567
transform 1 0 832 0 -1 770
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1711307567
transform 1 0 824 0 -1 770
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1711307567
transform 1 0 816 0 -1 770
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1711307567
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1711307567
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1711307567
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1711307567
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1711307567
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1711307567
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1711307567
transform 1 0 688 0 -1 770
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1711307567
transform 1 0 680 0 -1 770
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1711307567
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1711307567
transform 1 0 624 0 -1 770
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1711307567
transform 1 0 616 0 -1 770
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1711307567
transform 1 0 608 0 -1 770
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1711307567
transform 1 0 560 0 -1 770
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1711307567
transform 1 0 552 0 -1 770
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1711307567
transform 1 0 544 0 -1 770
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1711307567
transform 1 0 536 0 -1 770
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1711307567
transform 1 0 512 0 -1 770
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1711307567
transform 1 0 504 0 -1 770
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1711307567
transform 1 0 496 0 -1 770
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1711307567
transform 1 0 488 0 -1 770
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1711307567
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1711307567
transform 1 0 440 0 -1 770
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1711307567
transform 1 0 432 0 -1 770
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1711307567
transform 1 0 424 0 -1 770
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1711307567
transform 1 0 384 0 -1 770
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1711307567
transform 1 0 376 0 -1 770
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1711307567
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1711307567
transform 1 0 360 0 -1 770
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1711307567
transform 1 0 352 0 -1 770
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1711307567
transform 1 0 344 0 -1 770
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1711307567
transform 1 0 296 0 -1 770
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1711307567
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1711307567
transform 1 0 280 0 -1 770
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1711307567
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1711307567
transform 1 0 264 0 -1 770
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1711307567
transform 1 0 256 0 -1 770
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1711307567
transform 1 0 248 0 -1 770
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1711307567
transform 1 0 240 0 -1 770
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1711307567
transform 1 0 232 0 -1 770
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1711307567
transform 1 0 224 0 -1 770
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1711307567
transform 1 0 176 0 -1 770
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1711307567
transform 1 0 168 0 -1 770
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1711307567
transform 1 0 160 0 -1 770
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1711307567
transform 1 0 152 0 -1 770
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1711307567
transform 1 0 144 0 -1 770
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1711307567
transform 1 0 136 0 -1 770
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1711307567
transform 1 0 128 0 -1 770
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1711307567
transform 1 0 120 0 -1 770
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1711307567
transform 1 0 112 0 -1 770
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1711307567
transform 1 0 104 0 -1 770
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1711307567
transform 1 0 96 0 -1 770
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1711307567
transform 1 0 88 0 -1 770
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1711307567
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1711307567
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1711307567
transform 1 0 2696 0 1 570
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1711307567
transform 1 0 2688 0 1 570
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1711307567
transform 1 0 2512 0 1 570
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1711307567
transform 1 0 2504 0 1 570
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1711307567
transform 1 0 2440 0 1 570
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1711307567
transform 1 0 2336 0 1 570
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1711307567
transform 1 0 2328 0 1 570
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1711307567
transform 1 0 2272 0 1 570
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1711307567
transform 1 0 2240 0 1 570
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1711307567
transform 1 0 2232 0 1 570
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1711307567
transform 1 0 2224 0 1 570
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1711307567
transform 1 0 2184 0 1 570
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1711307567
transform 1 0 2176 0 1 570
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1711307567
transform 1 0 2168 0 1 570
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1711307567
transform 1 0 2120 0 1 570
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1711307567
transform 1 0 2112 0 1 570
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1711307567
transform 1 0 2104 0 1 570
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1711307567
transform 1 0 2080 0 1 570
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1711307567
transform 1 0 2072 0 1 570
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1711307567
transform 1 0 2024 0 1 570
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1711307567
transform 1 0 2016 0 1 570
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1711307567
transform 1 0 2008 0 1 570
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1711307567
transform 1 0 1944 0 1 570
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1711307567
transform 1 0 1936 0 1 570
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1711307567
transform 1 0 1928 0 1 570
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1711307567
transform 1 0 1920 0 1 570
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1711307567
transform 1 0 1912 0 1 570
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1711307567
transform 1 0 1856 0 1 570
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1711307567
transform 1 0 1848 0 1 570
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1711307567
transform 1 0 1840 0 1 570
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1711307567
transform 1 0 1832 0 1 570
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1711307567
transform 1 0 1776 0 1 570
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1711307567
transform 1 0 1768 0 1 570
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1711307567
transform 1 0 1760 0 1 570
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1711307567
transform 1 0 1752 0 1 570
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1711307567
transform 1 0 1696 0 1 570
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1711307567
transform 1 0 1688 0 1 570
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1711307567
transform 1 0 1680 0 1 570
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1711307567
transform 1 0 1648 0 1 570
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1711307567
transform 1 0 1640 0 1 570
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1711307567
transform 1 0 1632 0 1 570
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1711307567
transform 1 0 1584 0 1 570
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1711307567
transform 1 0 1576 0 1 570
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1711307567
transform 1 0 1568 0 1 570
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1711307567
transform 1 0 1512 0 1 570
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1711307567
transform 1 0 1504 0 1 570
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1711307567
transform 1 0 1496 0 1 570
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1711307567
transform 1 0 1432 0 1 570
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1711307567
transform 1 0 1424 0 1 570
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1711307567
transform 1 0 1416 0 1 570
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1711307567
transform 1 0 1360 0 1 570
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1711307567
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1711307567
transform 1 0 1312 0 1 570
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1711307567
transform 1 0 1272 0 1 570
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1711307567
transform 1 0 1264 0 1 570
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1711307567
transform 1 0 1256 0 1 570
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1711307567
transform 1 0 1208 0 1 570
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1711307567
transform 1 0 1200 0 1 570
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1711307567
transform 1 0 1192 0 1 570
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1711307567
transform 1 0 1144 0 1 570
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1711307567
transform 1 0 1120 0 1 570
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1711307567
transform 1 0 1112 0 1 570
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1711307567
transform 1 0 1104 0 1 570
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1711307567
transform 1 0 1064 0 1 570
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1711307567
transform 1 0 1056 0 1 570
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1711307567
transform 1 0 1016 0 1 570
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1711307567
transform 1 0 976 0 1 570
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1711307567
transform 1 0 968 0 1 570
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1711307567
transform 1 0 960 0 1 570
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1711307567
transform 1 0 952 0 1 570
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1711307567
transform 1 0 888 0 1 570
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1711307567
transform 1 0 880 0 1 570
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1711307567
transform 1 0 872 0 1 570
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1711307567
transform 1 0 864 0 1 570
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1711307567
transform 1 0 816 0 1 570
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1711307567
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1711307567
transform 1 0 800 0 1 570
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1711307567
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1711307567
transform 1 0 744 0 1 570
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1711307567
transform 1 0 736 0 1 570
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1711307567
transform 1 0 728 0 1 570
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1711307567
transform 1 0 680 0 1 570
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1711307567
transform 1 0 672 0 1 570
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1711307567
transform 1 0 664 0 1 570
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1711307567
transform 1 0 656 0 1 570
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1711307567
transform 1 0 648 0 1 570
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1711307567
transform 1 0 640 0 1 570
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1711307567
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1711307567
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1711307567
transform 1 0 576 0 1 570
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1711307567
transform 1 0 568 0 1 570
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1711307567
transform 1 0 528 0 1 570
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1711307567
transform 1 0 520 0 1 570
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1711307567
transform 1 0 512 0 1 570
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1711307567
transform 1 0 504 0 1 570
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1711307567
transform 1 0 464 0 1 570
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1711307567
transform 1 0 456 0 1 570
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1711307567
transform 1 0 416 0 1 570
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1711307567
transform 1 0 408 0 1 570
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1711307567
transform 1 0 400 0 1 570
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1711307567
transform 1 0 392 0 1 570
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1711307567
transform 1 0 336 0 1 570
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1711307567
transform 1 0 328 0 1 570
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1711307567
transform 1 0 320 0 1 570
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1711307567
transform 1 0 216 0 1 570
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1711307567
transform 1 0 208 0 1 570
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1711307567
transform 1 0 176 0 1 570
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1711307567
transform 1 0 168 0 1 570
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1711307567
transform 1 0 2752 0 -1 570
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1711307567
transform 1 0 2720 0 -1 570
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1711307567
transform 1 0 2712 0 -1 570
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1711307567
transform 1 0 2672 0 -1 570
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1711307567
transform 1 0 2664 0 -1 570
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1711307567
transform 1 0 2656 0 -1 570
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1711307567
transform 1 0 2648 0 -1 570
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1711307567
transform 1 0 2640 0 -1 570
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1711307567
transform 1 0 2632 0 -1 570
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1711307567
transform 1 0 2624 0 -1 570
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1711307567
transform 1 0 2616 0 -1 570
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1711307567
transform 1 0 2608 0 -1 570
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1711307567
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1711307567
transform 1 0 2592 0 -1 570
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1711307567
transform 1 0 2584 0 -1 570
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1711307567
transform 1 0 2544 0 -1 570
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1711307567
transform 1 0 2536 0 -1 570
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1711307567
transform 1 0 2528 0 -1 570
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1711307567
transform 1 0 2520 0 -1 570
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1711307567
transform 1 0 2512 0 -1 570
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1711307567
transform 1 0 2504 0 -1 570
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1711307567
transform 1 0 2496 0 -1 570
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1711307567
transform 1 0 2472 0 -1 570
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1711307567
transform 1 0 2464 0 -1 570
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1711307567
transform 1 0 2456 0 -1 570
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1711307567
transform 1 0 2448 0 -1 570
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1711307567
transform 1 0 2440 0 -1 570
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1711307567
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1711307567
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1711307567
transform 1 0 2416 0 -1 570
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1711307567
transform 1 0 2312 0 -1 570
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1711307567
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1711307567
transform 1 0 2296 0 -1 570
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1711307567
transform 1 0 2264 0 -1 570
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1711307567
transform 1 0 2224 0 -1 570
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1711307567
transform 1 0 2216 0 -1 570
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1711307567
transform 1 0 2208 0 -1 570
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1711307567
transform 1 0 2200 0 -1 570
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1711307567
transform 1 0 2152 0 -1 570
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1711307567
transform 1 0 2144 0 -1 570
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1711307567
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1711307567
transform 1 0 2128 0 -1 570
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1711307567
transform 1 0 2080 0 -1 570
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1711307567
transform 1 0 2072 0 -1 570
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1711307567
transform 1 0 2064 0 -1 570
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1711307567
transform 1 0 2056 0 -1 570
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1711307567
transform 1 0 2024 0 -1 570
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1711307567
transform 1 0 2016 0 -1 570
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1711307567
transform 1 0 2008 0 -1 570
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1711307567
transform 1 0 1960 0 -1 570
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1711307567
transform 1 0 1952 0 -1 570
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1711307567
transform 1 0 1944 0 -1 570
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1711307567
transform 1 0 1936 0 -1 570
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1711307567
transform 1 0 1928 0 -1 570
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1711307567
transform 1 0 1880 0 -1 570
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1711307567
transform 1 0 1872 0 -1 570
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1711307567
transform 1 0 1864 0 -1 570
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1711307567
transform 1 0 1856 0 -1 570
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1711307567
transform 1 0 1808 0 -1 570
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1711307567
transform 1 0 1800 0 -1 570
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1711307567
transform 1 0 1792 0 -1 570
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1711307567
transform 1 0 1744 0 -1 570
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1711307567
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1711307567
transform 1 0 1728 0 -1 570
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1711307567
transform 1 0 1720 0 -1 570
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1711307567
transform 1 0 1712 0 -1 570
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1711307567
transform 1 0 1648 0 -1 570
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1711307567
transform 1 0 1640 0 -1 570
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1711307567
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1711307567
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1711307567
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1711307567
transform 1 0 1576 0 -1 570
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1711307567
transform 1 0 1568 0 -1 570
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1711307567
transform 1 0 1528 0 -1 570
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1711307567
transform 1 0 1520 0 -1 570
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1711307567
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1711307567
transform 1 0 1504 0 -1 570
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1711307567
transform 1 0 1464 0 -1 570
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1711307567
transform 1 0 1456 0 -1 570
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1711307567
transform 1 0 1448 0 -1 570
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1711307567
transform 1 0 1440 0 -1 570
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1711307567
transform 1 0 1432 0 -1 570
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1711307567
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1711307567
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1711307567
transform 1 0 1376 0 -1 570
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1711307567
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1711307567
transform 1 0 1360 0 -1 570
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1711307567
transform 1 0 1352 0 -1 570
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1711307567
transform 1 0 1344 0 -1 570
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1711307567
transform 1 0 1336 0 -1 570
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1711307567
transform 1 0 1328 0 -1 570
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1711307567
transform 1 0 1320 0 -1 570
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1711307567
transform 1 0 1312 0 -1 570
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1711307567
transform 1 0 1280 0 -1 570
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1711307567
transform 1 0 1272 0 -1 570
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1711307567
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1711307567
transform 1 0 1256 0 -1 570
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1711307567
transform 1 0 1248 0 -1 570
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1711307567
transform 1 0 1208 0 -1 570
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1711307567
transform 1 0 1200 0 -1 570
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1711307567
transform 1 0 1160 0 -1 570
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1711307567
transform 1 0 1152 0 -1 570
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1711307567
transform 1 0 1144 0 -1 570
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1711307567
transform 1 0 1040 0 -1 570
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1711307567
transform 1 0 1032 0 -1 570
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1711307567
transform 1 0 928 0 -1 570
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1711307567
transform 1 0 920 0 -1 570
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1711307567
transform 1 0 912 0 -1 570
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1711307567
transform 1 0 872 0 -1 570
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1711307567
transform 1 0 864 0 -1 570
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1711307567
transform 1 0 856 0 -1 570
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1711307567
transform 1 0 816 0 -1 570
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1711307567
transform 1 0 808 0 -1 570
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1711307567
transform 1 0 800 0 -1 570
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1711307567
transform 1 0 792 0 -1 570
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1711307567
transform 1 0 752 0 -1 570
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1711307567
transform 1 0 744 0 -1 570
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1711307567
transform 1 0 736 0 -1 570
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1711307567
transform 1 0 728 0 -1 570
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1711307567
transform 1 0 720 0 -1 570
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1711307567
transform 1 0 616 0 -1 570
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1711307567
transform 1 0 608 0 -1 570
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1711307567
transform 1 0 600 0 -1 570
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1711307567
transform 1 0 496 0 -1 570
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1711307567
transform 1 0 488 0 -1 570
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1711307567
transform 1 0 480 0 -1 570
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1711307567
transform 1 0 472 0 -1 570
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1711307567
transform 1 0 464 0 -1 570
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1711307567
transform 1 0 456 0 -1 570
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1711307567
transform 1 0 448 0 -1 570
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1711307567
transform 1 0 408 0 -1 570
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1711307567
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1711307567
transform 1 0 392 0 -1 570
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1711307567
transform 1 0 384 0 -1 570
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1711307567
transform 1 0 376 0 -1 570
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1711307567
transform 1 0 352 0 -1 570
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1711307567
transform 1 0 344 0 -1 570
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1711307567
transform 1 0 336 0 -1 570
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1711307567
transform 1 0 304 0 -1 570
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1711307567
transform 1 0 296 0 -1 570
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1711307567
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1711307567
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1711307567
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1711307567
transform 1 0 264 0 -1 570
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1711307567
transform 1 0 256 0 -1 570
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1711307567
transform 1 0 248 0 -1 570
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1711307567
transform 1 0 240 0 -1 570
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1711307567
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1711307567
transform 1 0 176 0 -1 570
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1711307567
transform 1 0 168 0 -1 570
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1711307567
transform 1 0 2752 0 1 370
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1711307567
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1711307567
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1711307567
transform 1 0 2424 0 1 370
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1711307567
transform 1 0 2392 0 1 370
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1711307567
transform 1 0 2384 0 1 370
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1711307567
transform 1 0 2376 0 1 370
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1711307567
transform 1 0 2368 0 1 370
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1711307567
transform 1 0 2360 0 1 370
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1711307567
transform 1 0 2352 0 1 370
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1711307567
transform 1 0 2344 0 1 370
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1711307567
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1711307567
transform 1 0 2328 0 1 370
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1711307567
transform 1 0 2320 0 1 370
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1711307567
transform 1 0 2272 0 1 370
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1711307567
transform 1 0 2264 0 1 370
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1711307567
transform 1 0 2256 0 1 370
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1711307567
transform 1 0 2248 0 1 370
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1711307567
transform 1 0 2240 0 1 370
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1711307567
transform 1 0 2184 0 1 370
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1711307567
transform 1 0 2176 0 1 370
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1711307567
transform 1 0 2168 0 1 370
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1711307567
transform 1 0 2136 0 1 370
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1711307567
transform 1 0 2128 0 1 370
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1711307567
transform 1 0 2120 0 1 370
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1711307567
transform 1 0 2112 0 1 370
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1711307567
transform 1 0 2008 0 1 370
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1711307567
transform 1 0 2000 0 1 370
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1711307567
transform 1 0 1968 0 1 370
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1711307567
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1711307567
transform 1 0 1912 0 1 370
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1711307567
transform 1 0 1904 0 1 370
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1711307567
transform 1 0 1896 0 1 370
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1711307567
transform 1 0 1888 0 1 370
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1711307567
transform 1 0 1880 0 1 370
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1711307567
transform 1 0 1832 0 1 370
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1711307567
transform 1 0 1824 0 1 370
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1711307567
transform 1 0 1816 0 1 370
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1711307567
transform 1 0 1808 0 1 370
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1711307567
transform 1 0 1800 0 1 370
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1711307567
transform 1 0 1792 0 1 370
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1711307567
transform 1 0 1768 0 1 370
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1711307567
transform 1 0 1760 0 1 370
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1711307567
transform 1 0 1752 0 1 370
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1711307567
transform 1 0 1712 0 1 370
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1711307567
transform 1 0 1704 0 1 370
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1711307567
transform 1 0 1696 0 1 370
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1711307567
transform 1 0 1688 0 1 370
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1711307567
transform 1 0 1680 0 1 370
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1711307567
transform 1 0 1672 0 1 370
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1711307567
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1711307567
transform 1 0 1656 0 1 370
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1711307567
transform 1 0 1648 0 1 370
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1711307567
transform 1 0 1616 0 1 370
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1711307567
transform 1 0 1608 0 1 370
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1711307567
transform 1 0 1600 0 1 370
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1711307567
transform 1 0 1592 0 1 370
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1711307567
transform 1 0 1560 0 1 370
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1711307567
transform 1 0 1552 0 1 370
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1711307567
transform 1 0 1544 0 1 370
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1711307567
transform 1 0 1536 0 1 370
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1711307567
transform 1 0 1528 0 1 370
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1711307567
transform 1 0 1496 0 1 370
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1711307567
transform 1 0 1488 0 1 370
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1711307567
transform 1 0 1480 0 1 370
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1711307567
transform 1 0 1376 0 1 370
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1711307567
transform 1 0 1272 0 1 370
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1711307567
transform 1 0 1264 0 1 370
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1711307567
transform 1 0 1256 0 1 370
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1711307567
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1711307567
transform 1 0 1192 0 1 370
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1711307567
transform 1 0 1184 0 1 370
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1711307567
transform 1 0 1176 0 1 370
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1711307567
transform 1 0 1120 0 1 370
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1711307567
transform 1 0 1112 0 1 370
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1711307567
transform 1 0 1104 0 1 370
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1711307567
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1711307567
transform 1 0 1088 0 1 370
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1711307567
transform 1 0 1080 0 1 370
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1711307567
transform 1 0 1072 0 1 370
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1711307567
transform 1 0 1040 0 1 370
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1711307567
transform 1 0 1008 0 1 370
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1711307567
transform 1 0 1000 0 1 370
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1711307567
transform 1 0 992 0 1 370
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1711307567
transform 1 0 952 0 1 370
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1711307567
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1711307567
transform 1 0 936 0 1 370
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1711307567
transform 1 0 928 0 1 370
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1711307567
transform 1 0 920 0 1 370
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1711307567
transform 1 0 912 0 1 370
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1711307567
transform 1 0 848 0 1 370
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1711307567
transform 1 0 840 0 1 370
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1711307567
transform 1 0 832 0 1 370
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1711307567
transform 1 0 824 0 1 370
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1711307567
transform 1 0 816 0 1 370
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1711307567
transform 1 0 768 0 1 370
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1711307567
transform 1 0 664 0 1 370
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1711307567
transform 1 0 656 0 1 370
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1711307567
transform 1 0 648 0 1 370
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1711307567
transform 1 0 544 0 1 370
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1711307567
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1711307567
transform 1 0 528 0 1 370
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1711307567
transform 1 0 328 0 1 370
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1711307567
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1711307567
transform 1 0 120 0 1 370
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1711307567
transform 1 0 112 0 1 370
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1711307567
transform 1 0 104 0 1 370
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1711307567
transform 1 0 96 0 1 370
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1711307567
transform 1 0 88 0 1 370
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1711307567
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1711307567
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1711307567
transform 1 0 2656 0 -1 370
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1711307567
transform 1 0 2584 0 -1 370
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1711307567
transform 1 0 2576 0 -1 370
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1711307567
transform 1 0 2536 0 -1 370
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1711307567
transform 1 0 2528 0 -1 370
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1711307567
transform 1 0 2472 0 -1 370
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1711307567
transform 1 0 2464 0 -1 370
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1711307567
transform 1 0 2408 0 -1 370
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1711307567
transform 1 0 2304 0 -1 370
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1711307567
transform 1 0 2296 0 -1 370
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1711307567
transform 1 0 2208 0 -1 370
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1711307567
transform 1 0 2200 0 -1 370
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1711307567
transform 1 0 2096 0 -1 370
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1711307567
transform 1 0 2088 0 -1 370
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1711307567
transform 1 0 2080 0 -1 370
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1711307567
transform 1 0 2048 0 -1 370
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1711307567
transform 1 0 2040 0 -1 370
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1711307567
transform 1 0 2032 0 -1 370
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1711307567
transform 1 0 2000 0 -1 370
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1711307567
transform 1 0 1952 0 -1 370
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1711307567
transform 1 0 1944 0 -1 370
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1711307567
transform 1 0 1936 0 -1 370
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1711307567
transform 1 0 1888 0 -1 370
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1711307567
transform 1 0 1880 0 -1 370
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1711307567
transform 1 0 1872 0 -1 370
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1711307567
transform 1 0 1864 0 -1 370
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1711307567
transform 1 0 1760 0 -1 370
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1711307567
transform 1 0 1520 0 -1 370
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1711307567
transform 1 0 1464 0 -1 370
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1711307567
transform 1 0 1456 0 -1 370
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1711307567
transform 1 0 1400 0 -1 370
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1711307567
transform 1 0 1176 0 -1 370
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1711307567
transform 1 0 1144 0 -1 370
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1711307567
transform 1 0 1040 0 -1 370
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1711307567
transform 1 0 1032 0 -1 370
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1711307567
transform 1 0 912 0 -1 370
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1711307567
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1711307567
transform 1 0 896 0 -1 370
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1711307567
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1711307567
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1711307567
transform 1 0 752 0 -1 370
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1711307567
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1711307567
transform 1 0 712 0 -1 370
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1711307567
transform 1 0 704 0 -1 370
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1711307567
transform 1 0 696 0 -1 370
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1711307567
transform 1 0 688 0 -1 370
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1711307567
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1711307567
transform 1 0 648 0 -1 370
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1711307567
transform 1 0 616 0 -1 370
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1711307567
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1711307567
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1711307567
transform 1 0 592 0 -1 370
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1711307567
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1711307567
transform 1 0 576 0 -1 370
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1711307567
transform 1 0 520 0 -1 370
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1711307567
transform 1 0 512 0 -1 370
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1711307567
transform 1 0 504 0 -1 370
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1711307567
transform 1 0 496 0 -1 370
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1711307567
transform 1 0 488 0 -1 370
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1711307567
transform 1 0 456 0 -1 370
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1711307567
transform 1 0 448 0 -1 370
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1711307567
transform 1 0 440 0 -1 370
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1711307567
transform 1 0 408 0 -1 370
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1711307567
transform 1 0 400 0 -1 370
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1711307567
transform 1 0 392 0 -1 370
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1711307567
transform 1 0 384 0 -1 370
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1711307567
transform 1 0 352 0 -1 370
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1711307567
transform 1 0 344 0 -1 370
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1711307567
transform 1 0 336 0 -1 370
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1711307567
transform 1 0 328 0 -1 370
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1711307567
transform 1 0 320 0 -1 370
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1711307567
transform 1 0 288 0 -1 370
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1711307567
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1711307567
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1711307567
transform 1 0 264 0 -1 370
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1711307567
transform 1 0 232 0 -1 370
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1711307567
transform 1 0 224 0 -1 370
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1711307567
transform 1 0 216 0 -1 370
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1711307567
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1711307567
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1711307567
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1711307567
transform 1 0 160 0 -1 370
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1711307567
transform 1 0 152 0 -1 370
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1711307567
transform 1 0 144 0 -1 370
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1711307567
transform 1 0 136 0 -1 370
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1711307567
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1711307567
transform 1 0 120 0 -1 370
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1711307567
transform 1 0 112 0 -1 370
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1711307567
transform 1 0 104 0 -1 370
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1711307567
transform 1 0 96 0 -1 370
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1711307567
transform 1 0 88 0 -1 370
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1711307567
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1711307567
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1711307567
transform 1 0 2752 0 1 170
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1711307567
transform 1 0 2744 0 1 170
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1711307567
transform 1 0 2736 0 1 170
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1711307567
transform 1 0 2728 0 1 170
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1711307567
transform 1 0 2720 0 1 170
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1711307567
transform 1 0 2712 0 1 170
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1711307567
transform 1 0 2704 0 1 170
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1711307567
transform 1 0 2600 0 1 170
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1711307567
transform 1 0 2592 0 1 170
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1711307567
transform 1 0 2584 0 1 170
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1711307567
transform 1 0 2552 0 1 170
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1711307567
transform 1 0 2512 0 1 170
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1711307567
transform 1 0 2504 0 1 170
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1711307567
transform 1 0 2496 0 1 170
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1711307567
transform 1 0 2488 0 1 170
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1711307567
transform 1 0 2480 0 1 170
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1711307567
transform 1 0 2440 0 1 170
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1711307567
transform 1 0 2432 0 1 170
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1711307567
transform 1 0 2424 0 1 170
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1711307567
transform 1 0 2416 0 1 170
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1711307567
transform 1 0 2408 0 1 170
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1711307567
transform 1 0 2400 0 1 170
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1711307567
transform 1 0 2392 0 1 170
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1711307567
transform 1 0 2384 0 1 170
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1711307567
transform 1 0 2376 0 1 170
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1711307567
transform 1 0 2368 0 1 170
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1711307567
transform 1 0 2360 0 1 170
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1711307567
transform 1 0 2352 0 1 170
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1711307567
transform 1 0 2344 0 1 170
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1711307567
transform 1 0 2304 0 1 170
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1711307567
transform 1 0 2296 0 1 170
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1711307567
transform 1 0 2288 0 1 170
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1711307567
transform 1 0 2280 0 1 170
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1711307567
transform 1 0 2240 0 1 170
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1711307567
transform 1 0 2232 0 1 170
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1711307567
transform 1 0 2224 0 1 170
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1711307567
transform 1 0 2192 0 1 170
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1711307567
transform 1 0 2184 0 1 170
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1711307567
transform 1 0 2176 0 1 170
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1711307567
transform 1 0 2168 0 1 170
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1711307567
transform 1 0 2160 0 1 170
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1711307567
transform 1 0 2152 0 1 170
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1711307567
transform 1 0 2128 0 1 170
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1711307567
transform 1 0 2120 0 1 170
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1711307567
transform 1 0 2112 0 1 170
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1711307567
transform 1 0 2008 0 1 170
box -8 -3 16 105
use FILL  FILL_3130
timestamp 1711307567
transform 1 0 2000 0 1 170
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1711307567
transform 1 0 1992 0 1 170
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1711307567
transform 1 0 1984 0 1 170
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1711307567
transform 1 0 1976 0 1 170
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1711307567
transform 1 0 1928 0 1 170
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1711307567
transform 1 0 1920 0 1 170
box -8 -3 16 105
use FILL  FILL_3136
timestamp 1711307567
transform 1 0 1912 0 1 170
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1711307567
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1711307567
transform 1 0 1800 0 1 170
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1711307567
transform 1 0 1792 0 1 170
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1711307567
transform 1 0 1784 0 1 170
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1711307567
transform 1 0 1776 0 1 170
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1711307567
transform 1 0 1768 0 1 170
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1711307567
transform 1 0 1760 0 1 170
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1711307567
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1711307567
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1711307567
transform 1 0 1736 0 1 170
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1711307567
transform 1 0 1728 0 1 170
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1711307567
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1711307567
transform 1 0 1712 0 1 170
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1711307567
transform 1 0 1704 0 1 170
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1711307567
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1711307567
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1711307567
transform 1 0 1680 0 1 170
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1711307567
transform 1 0 1672 0 1 170
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1711307567
transform 1 0 1664 0 1 170
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1711307567
transform 1 0 1656 0 1 170
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1711307567
transform 1 0 1648 0 1 170
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1711307567
transform 1 0 1640 0 1 170
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1711307567
transform 1 0 1632 0 1 170
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1711307567
transform 1 0 1624 0 1 170
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1711307567
transform 1 0 1584 0 1 170
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1711307567
transform 1 0 1576 0 1 170
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1711307567
transform 1 0 1568 0 1 170
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1711307567
transform 1 0 1560 0 1 170
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1711307567
transform 1 0 1552 0 1 170
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1711307567
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1711307567
transform 1 0 1536 0 1 170
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1711307567
transform 1 0 1528 0 1 170
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1711307567
transform 1 0 1520 0 1 170
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1711307567
transform 1 0 1512 0 1 170
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1711307567
transform 1 0 1504 0 1 170
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1711307567
transform 1 0 1496 0 1 170
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1711307567
transform 1 0 1488 0 1 170
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1711307567
transform 1 0 1480 0 1 170
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1711307567
transform 1 0 1440 0 1 170
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1711307567
transform 1 0 1432 0 1 170
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1711307567
transform 1 0 1408 0 1 170
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1711307567
transform 1 0 1400 0 1 170
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1711307567
transform 1 0 1392 0 1 170
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1711307567
transform 1 0 1360 0 1 170
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1711307567
transform 1 0 1352 0 1 170
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1711307567
transform 1 0 1344 0 1 170
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1711307567
transform 1 0 1336 0 1 170
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1711307567
transform 1 0 1328 0 1 170
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1711307567
transform 1 0 1288 0 1 170
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1711307567
transform 1 0 1280 0 1 170
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1711307567
transform 1 0 1272 0 1 170
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1711307567
transform 1 0 1248 0 1 170
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1711307567
transform 1 0 1240 0 1 170
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1711307567
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1711307567
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1711307567
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1711307567
transform 1 0 1184 0 1 170
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1711307567
transform 1 0 1176 0 1 170
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1711307567
transform 1 0 1168 0 1 170
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1711307567
transform 1 0 1128 0 1 170
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1711307567
transform 1 0 1120 0 1 170
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1711307567
transform 1 0 1112 0 1 170
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1711307567
transform 1 0 1080 0 1 170
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1711307567
transform 1 0 1072 0 1 170
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1711307567
transform 1 0 1064 0 1 170
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1711307567
transform 1 0 1032 0 1 170
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1711307567
transform 1 0 1024 0 1 170
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1711307567
transform 1 0 984 0 1 170
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1711307567
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1711307567
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1711307567
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1711307567
transform 1 0 952 0 1 170
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1711307567
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1711307567
transform 1 0 840 0 1 170
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1711307567
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1711307567
transform 1 0 824 0 1 170
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1711307567
transform 1 0 816 0 1 170
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1711307567
transform 1 0 808 0 1 170
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1711307567
transform 1 0 800 0 1 170
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1711307567
transform 1 0 792 0 1 170
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1711307567
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1711307567
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1711307567
transform 1 0 736 0 1 170
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1711307567
transform 1 0 728 0 1 170
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1711307567
transform 1 0 720 0 1 170
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1711307567
transform 1 0 712 0 1 170
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1711307567
transform 1 0 704 0 1 170
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1711307567
transform 1 0 696 0 1 170
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1711307567
transform 1 0 656 0 1 170
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1711307567
transform 1 0 648 0 1 170
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1711307567
transform 1 0 640 0 1 170
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1711307567
transform 1 0 616 0 1 170
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1711307567
transform 1 0 608 0 1 170
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1711307567
transform 1 0 568 0 1 170
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1711307567
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1711307567
transform 1 0 552 0 1 170
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1711307567
transform 1 0 544 0 1 170
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1711307567
transform 1 0 520 0 1 170
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1711307567
transform 1 0 512 0 1 170
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1711307567
transform 1 0 504 0 1 170
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1711307567
transform 1 0 496 0 1 170
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1711307567
transform 1 0 488 0 1 170
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1711307567
transform 1 0 448 0 1 170
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1711307567
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1711307567
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1711307567
transform 1 0 408 0 1 170
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1711307567
transform 1 0 400 0 1 170
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1711307567
transform 1 0 392 0 1 170
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1711307567
transform 1 0 384 0 1 170
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1711307567
transform 1 0 376 0 1 170
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1711307567
transform 1 0 368 0 1 170
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1711307567
transform 1 0 328 0 1 170
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1711307567
transform 1 0 320 0 1 170
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1711307567
transform 1 0 312 0 1 170
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1711307567
transform 1 0 304 0 1 170
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1711307567
transform 1 0 280 0 1 170
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1711307567
transform 1 0 272 0 1 170
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1711307567
transform 1 0 264 0 1 170
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1711307567
transform 1 0 256 0 1 170
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1711307567
transform 1 0 248 0 1 170
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1711307567
transform 1 0 208 0 1 170
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1711307567
transform 1 0 200 0 1 170
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1711307567
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1711307567
transform 1 0 184 0 1 170
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1711307567
transform 1 0 160 0 1 170
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1711307567
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1711307567
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1711307567
transform 1 0 136 0 1 170
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1711307567
transform 1 0 128 0 1 170
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1711307567
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1711307567
transform 1 0 112 0 1 170
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1711307567
transform 1 0 104 0 1 170
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1711307567
transform 1 0 96 0 1 170
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1711307567
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1711307567
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1711307567
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1711307567
transform 1 0 2656 0 -1 170
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1711307567
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1711307567
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1711307567
transform 1 0 2632 0 -1 170
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1711307567
transform 1 0 2624 0 -1 170
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1711307567
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1711307567
transform 1 0 2560 0 -1 170
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1711307567
transform 1 0 2552 0 -1 170
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1711307567
transform 1 0 2544 0 -1 170
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1711307567
transform 1 0 2536 0 -1 170
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1711307567
transform 1 0 2472 0 -1 170
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1711307567
transform 1 0 2464 0 -1 170
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1711307567
transform 1 0 2456 0 -1 170
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1711307567
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1711307567
transform 1 0 2440 0 -1 170
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1711307567
transform 1 0 2432 0 -1 170
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1711307567
transform 1 0 2360 0 -1 170
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1711307567
transform 1 0 2352 0 -1 170
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1711307567
transform 1 0 2248 0 -1 170
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1711307567
transform 1 0 2240 0 -1 170
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1711307567
transform 1 0 2136 0 -1 170
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1711307567
transform 1 0 2128 0 -1 170
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1711307567
transform 1 0 2096 0 -1 170
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1711307567
transform 1 0 2088 0 -1 170
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1711307567
transform 1 0 2080 0 -1 170
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1711307567
transform 1 0 2072 0 -1 170
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1711307567
transform 1 0 2064 0 -1 170
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1711307567
transform 1 0 2056 0 -1 170
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1711307567
transform 1 0 2048 0 -1 170
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1711307567
transform 1 0 2040 0 -1 170
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1711307567
transform 1 0 1936 0 -1 170
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1711307567
transform 1 0 1928 0 -1 170
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1711307567
transform 1 0 1920 0 -1 170
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1711307567
transform 1 0 1912 0 -1 170
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1711307567
transform 1 0 1864 0 -1 170
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1711307567
transform 1 0 1856 0 -1 170
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1711307567
transform 1 0 1848 0 -1 170
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1711307567
transform 1 0 1840 0 -1 170
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1711307567
transform 1 0 1832 0 -1 170
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1711307567
transform 1 0 1632 0 -1 170
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1711307567
transform 1 0 1624 0 -1 170
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1711307567
transform 1 0 1616 0 -1 170
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1711307567
transform 1 0 1568 0 -1 170
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1711307567
transform 1 0 1560 0 -1 170
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1711307567
transform 1 0 1456 0 -1 170
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1711307567
transform 1 0 1352 0 -1 170
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1711307567
transform 1 0 1248 0 -1 170
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1711307567
transform 1 0 1240 0 -1 170
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1711307567
transform 1 0 1136 0 -1 170
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1711307567
transform 1 0 1128 0 -1 170
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1711307567
transform 1 0 1120 0 -1 170
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1711307567
transform 1 0 1112 0 -1 170
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1711307567
transform 1 0 1088 0 -1 170
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1711307567
transform 1 0 1080 0 -1 170
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1711307567
transform 1 0 1072 0 -1 170
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1711307567
transform 1 0 1064 0 -1 170
box -8 -3 16 105
use FILL  FILL_3329
timestamp 1711307567
transform 1 0 1040 0 -1 170
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1711307567
transform 1 0 1032 0 -1 170
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1711307567
transform 1 0 1024 0 -1 170
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1711307567
transform 1 0 1016 0 -1 170
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1711307567
transform 1 0 912 0 -1 170
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1711307567
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1711307567
transform 1 0 896 0 -1 170
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1711307567
transform 1 0 888 0 -1 170
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1711307567
transform 1 0 880 0 -1 170
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1711307567
transform 1 0 872 0 -1 170
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1711307567
transform 1 0 864 0 -1 170
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1711307567
transform 1 0 760 0 -1 170
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1711307567
transform 1 0 736 0 -1 170
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1711307567
transform 1 0 728 0 -1 170
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1711307567
transform 1 0 720 0 -1 170
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1711307567
transform 1 0 616 0 -1 170
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1711307567
transform 1 0 608 0 -1 170
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1711307567
transform 1 0 600 0 -1 170
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1711307567
transform 1 0 496 0 -1 170
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1711307567
transform 1 0 488 0 -1 170
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1711307567
transform 1 0 480 0 -1 170
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1711307567
transform 1 0 472 0 -1 170
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1711307567
transform 1 0 368 0 -1 170
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1711307567
transform 1 0 360 0 -1 170
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1711307567
transform 1 0 352 0 -1 170
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1711307567
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1711307567
transform 1 0 240 0 -1 170
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1711307567
transform 1 0 232 0 -1 170
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1711307567
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1711307567
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1711307567
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1711307567
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1711307567
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1711307567
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1711307567
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1711307567
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1711307567
transform 1 0 2672 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1711307567
transform 1 0 2680 0 1 2170
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1711307567
transform 1 0 2664 0 -1 2170
box -5 -3 84 105
use INVX2  INVX2_0
timestamp 1711307567
transform 1 0 2744 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1711307567
transform 1 0 2344 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1711307567
transform 1 0 1640 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1711307567
transform 1 0 1336 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1711307567
transform 1 0 1408 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1711307567
transform 1 0 1920 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1711307567
transform 1 0 1648 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1711307567
transform 1 0 2056 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1711307567
transform 1 0 1904 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1711307567
transform 1 0 1648 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1711307567
transform 1 0 896 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1711307567
transform 1 0 1432 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1711307567
transform 1 0 1616 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1711307567
transform 1 0 320 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1711307567
transform 1 0 1048 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1711307567
transform 1 0 1744 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1711307567
transform 1 0 856 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1711307567
transform 1 0 1448 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1711307567
transform 1 0 1904 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1711307567
transform 1 0 1312 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1711307567
transform 1 0 1592 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1711307567
transform 1 0 1640 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1711307567
transform 1 0 1120 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1711307567
transform 1 0 1560 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1711307567
transform 1 0 1768 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1711307567
transform 1 0 1848 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1711307567
transform 1 0 472 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1711307567
transform 1 0 952 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1711307567
transform 1 0 1392 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1711307567
transform 1 0 1136 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1711307567
transform 1 0 1600 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1711307567
transform 1 0 744 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1711307567
transform 1 0 2064 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1711307567
transform 1 0 1008 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1711307567
transform 1 0 1736 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1711307567
transform 1 0 480 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1711307567
transform 1 0 1688 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1711307567
transform 1 0 1904 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1711307567
transform 1 0 2080 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1711307567
transform 1 0 1616 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1711307567
transform 1 0 600 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1711307567
transform 1 0 2064 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1711307567
transform 1 0 976 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1711307567
transform 1 0 1968 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1711307567
transform 1 0 2352 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1711307567
transform 1 0 2376 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1711307567
transform 1 0 960 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1711307567
transform 1 0 1672 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1711307567
transform 1 0 2280 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1711307567
transform 1 0 2160 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1711307567
transform 1 0 1800 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1711307567
transform 1 0 504 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1711307567
transform 1 0 1064 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1711307567
transform 1 0 1712 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1711307567
transform 1 0 2376 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1711307567
transform 1 0 2080 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1711307567
transform 1 0 864 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1711307567
transform 1 0 1680 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1711307567
transform 1 0 1952 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1711307567
transform 1 0 2264 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1711307567
transform 1 0 384 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1711307567
transform 1 0 904 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1711307567
transform 1 0 1472 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1711307567
transform 1 0 2088 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1711307567
transform 1 0 1488 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1711307567
transform 1 0 2528 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1711307567
transform 1 0 2480 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1711307567
transform 1 0 2600 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1711307567
transform 1 0 2664 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1711307567
transform 1 0 2648 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1711307567
transform 1 0 2624 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1711307567
transform 1 0 2712 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1711307567
transform 1 0 2552 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1711307567
transform 1 0 360 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1711307567
transform 1 0 192 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1711307567
transform 1 0 88 0 1 970
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1711307567
transform 1 0 192 0 1 770
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1711307567
transform 1 0 288 0 1 170
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1711307567
transform 1 0 168 0 1 170
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1711307567
transform 1 0 528 0 1 170
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1711307567
transform 1 0 416 0 1 170
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1711307567
transform 1 0 800 0 1 370
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1711307567
transform 1 0 744 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1711307567
transform 1 0 624 0 1 170
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1711307567
transform 1 0 1016 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1711307567
transform 1 0 1048 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1711307567
transform 1 0 1096 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1711307567
transform 1 0 1208 0 1 370
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1711307567
transform 1 0 1256 0 1 170
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1711307567
transform 1 0 1600 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1711307567
transform 1 0 1416 0 1 170
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1711307567
transform 1 0 1504 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1711307567
transform 1 0 1744 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1711307567
transform 1 0 1896 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1711307567
transform 1 0 1864 0 1 370
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1711307567
transform 1 0 1960 0 1 170
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1711307567
transform 1 0 2024 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1711307567
transform 1 0 2072 0 1 770
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1711307567
transform 1 0 2632 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1711307567
transform 1 0 2624 0 1 770
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1711307567
transform 1 0 2512 0 1 970
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1711307567
transform 1 0 2304 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1711307567
transform 1 0 2560 0 1 970
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1711307567
transform 1 0 2600 0 1 970
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1711307567
transform 1 0 2312 0 1 570
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1711307567
transform 1 0 2304 0 1 370
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1711307567
transform 1 0 2416 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1711307567
transform 1 0 2480 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1711307567
transform 1 0 2544 0 1 370
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1711307567
transform 1 0 2520 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1711307567
transform 1 0 2512 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1711307567
transform 1 0 2448 0 1 170
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1711307567
transform 1 0 2464 0 1 170
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1711307567
transform 1 0 1696 0 1 770
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1711307567
transform 1 0 1648 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1711307567
transform 1 0 1584 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1711307567
transform 1 0 1736 0 1 570
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1711307567
transform 1 0 1936 0 1 970
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1711307567
transform 1 0 1816 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1711307567
transform 1 0 2328 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1711307567
transform 1 0 1976 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1711307567
transform 1 0 2472 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1711307567
transform 1 0 2048 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1711307567
transform 1 0 1856 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1711307567
transform 1 0 1864 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1711307567
transform 1 0 2272 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1711307567
transform 1 0 1752 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1711307567
transform 1 0 1736 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1711307567
transform 1 0 1640 0 1 770
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1711307567
transform 1 0 1992 0 1 970
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1711307567
transform 1 0 376 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1711307567
transform 1 0 216 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1711307567
transform 1 0 344 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1711307567
transform 1 0 288 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1711307567
transform 1 0 2192 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1711307567
transform 1 0 264 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1711307567
transform 1 0 192 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1711307567
transform 1 0 456 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1711307567
transform 1 0 352 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1711307567
transform 1 0 248 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1711307567
transform 1 0 248 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1711307567
transform 1 0 416 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1711307567
transform 1 0 456 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1711307567
transform 1 0 512 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1711307567
transform 1 0 520 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1711307567
transform 1 0 472 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1711307567
transform 1 0 568 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1711307567
transform 1 0 432 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1711307567
transform 1 0 456 0 1 770
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1711307567
transform 1 0 616 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1711307567
transform 1 0 584 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1711307567
transform 1 0 328 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1711307567
transform 1 0 608 0 1 770
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1711307567
transform 1 0 472 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1711307567
transform 1 0 712 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1711307567
transform 1 0 728 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1711307567
transform 1 0 800 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1711307567
transform 1 0 616 0 1 970
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1711307567
transform 1 0 736 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1711307567
transform 1 0 544 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1711307567
transform 1 0 632 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1711307567
transform 1 0 768 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1711307567
transform 1 0 896 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1711307567
transform 1 0 640 0 1 770
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1711307567
transform 1 0 696 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1711307567
transform 1 0 992 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1711307567
transform 1 0 520 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1711307567
transform 1 0 2312 0 1 770
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1711307567
transform 1 0 2232 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1711307567
transform 1 0 920 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1711307567
transform 1 0 1072 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1711307567
transform 1 0 1032 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1711307567
transform 1 0 1088 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1711307567
transform 1 0 952 0 1 770
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1711307567
transform 1 0 1176 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1711307567
transform 1 0 1096 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1711307567
transform 1 0 1144 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1711307567
transform 1 0 696 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1711307567
transform 1 0 816 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1711307567
transform 1 0 1272 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1711307567
transform 1 0 1200 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1711307567
transform 1 0 1168 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1711307567
transform 1 0 976 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1711307567
transform 1 0 936 0 1 570
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1711307567
transform 1 0 1088 0 1 770
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1711307567
transform 1 0 1128 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1711307567
transform 1 0 1440 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1711307567
transform 1 0 1104 0 1 770
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1711307567
transform 1 0 976 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1711307567
transform 1 0 1224 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1711307567
transform 1 0 1152 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1711307567
transform 1 0 1368 0 1 570
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1711307567
transform 1 0 1128 0 1 570
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1711307567
transform 1 0 1784 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1711307567
transform 1 0 1392 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1711307567
transform 1 0 1488 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1711307567
transform 1 0 1248 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1711307567
transform 1 0 1504 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1711307567
transform 1 0 1656 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1711307567
transform 1 0 1816 0 1 570
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1711307567
transform 1 0 1592 0 1 570
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1711307567
transform 1 0 1896 0 1 570
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1711307567
transform 1 0 2088 0 1 570
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1711307567
transform 1 0 1992 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1711307567
transform 1 0 1552 0 1 570
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1711307567
transform 1 0 2440 0 1 770
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1711307567
transform 1 0 1736 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1711307567
transform 1 0 1568 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1711307567
transform 1 0 1776 0 1 370
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1711307567
transform 1 0 2072 0 1 970
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1711307567
transform 1 0 2568 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1711307567
transform 1 0 1936 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1711307567
transform 1 0 2160 0 1 770
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1711307567
transform 1 0 2648 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1711307567
transform 1 0 2728 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1711307567
transform 1 0 2704 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1711307567
transform 1 0 2728 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1711307567
transform 1 0 2680 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1711307567
transform 1 0 2624 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1711307567
transform 1 0 2616 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1711307567
transform 1 0 2576 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1711307567
transform 1 0 2536 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1711307567
transform 1 0 1440 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_223
timestamp 1711307567
transform 1 0 136 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1711307567
transform 1 0 128 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_225
timestamp 1711307567
transform 1 0 128 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_226
timestamp 1711307567
transform 1 0 2024 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_227
timestamp 1711307567
transform 1 0 2240 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_228
timestamp 1711307567
transform 1 0 2320 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_229
timestamp 1711307567
transform 1 0 2104 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_230
timestamp 1711307567
transform 1 0 2216 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1711307567
transform 1 0 2704 0 1 570
box -9 -3 26 105
use INVX2  INVX2_232
timestamp 1711307567
transform 1 0 1960 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1711307567
transform 1 0 2448 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_234
timestamp 1711307567
transform 1 0 2064 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_235
timestamp 1711307567
transform 1 0 2144 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_236
timestamp 1711307567
transform 1 0 1032 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_237
timestamp 1711307567
transform 1 0 752 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1711307567
transform 1 0 1176 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_239
timestamp 1711307567
transform 1 0 1760 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1711307567
transform 1 0 2136 0 1 170
box -9 -3 26 105
use INVX2  INVX2_241
timestamp 1711307567
transform 1 0 2304 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_242
timestamp 1711307567
transform 1 0 2352 0 1 970
box -9 -3 26 105
use INVX2  INVX2_243
timestamp 1711307567
transform 1 0 2288 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_244
timestamp 1711307567
transform 1 0 2264 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_245
timestamp 1711307567
transform 1 0 1952 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1711307567
transform 1 0 2720 0 1 570
box -9 -3 26 105
use INVX2  INVX2_247
timestamp 1711307567
transform 1 0 2680 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_248
timestamp 1711307567
transform 1 0 2696 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_249
timestamp 1711307567
transform 1 0 2152 0 -1 1170
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1711307567
transform 1 0 2700 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1711307567
transform 1 0 2692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1711307567
transform 1 0 2708 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1711307567
transform 1 0 2684 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1711307567
transform 1 0 2700 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1711307567
transform 1 0 2604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1711307567
transform 1 0 2532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1711307567
transform 1 0 2396 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1711307567
transform 1 0 2380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1711307567
transform 1 0 2372 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1711307567
transform 1 0 2356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1711307567
transform 1 0 2332 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1711307567
transform 1 0 2316 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1711307567
transform 1 0 2516 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1711307567
transform 1 0 2412 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1711307567
transform 1 0 2380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1711307567
transform 1 0 2364 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1711307567
transform 1 0 2308 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1711307567
transform 1 0 2284 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1711307567
transform 1 0 2452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1711307567
transform 1 0 2404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1711307567
transform 1 0 2372 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1711307567
transform 1 0 2348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1711307567
transform 1 0 2348 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1711307567
transform 1 0 2284 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1711307567
transform 1 0 2388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1711307567
transform 1 0 2068 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1711307567
transform 1 0 1980 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1711307567
transform 1 0 2292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1711307567
transform 1 0 2084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1711307567
transform 1 0 1996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1711307567
transform 1 0 1956 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1711307567
transform 1 0 2324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1711307567
transform 1 0 2276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1711307567
transform 1 0 2060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1711307567
transform 1 0 2004 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1711307567
transform 1 0 1964 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1711307567
transform 1 0 1852 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1711307567
transform 1 0 1836 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1711307567
transform 1 0 2540 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1711307567
transform 1 0 2420 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1711307567
transform 1 0 2164 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1711307567
transform 1 0 2124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1711307567
transform 1 0 2124 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1711307567
transform 1 0 2084 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1711307567
transform 1 0 2012 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1711307567
transform 1 0 1996 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1711307567
transform 1 0 1964 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1711307567
transform 1 0 1924 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1711307567
transform 1 0 1916 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1711307567
transform 1 0 2452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1711307567
transform 1 0 2172 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1711307567
transform 1 0 2172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1711307567
transform 1 0 1700 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1711307567
transform 1 0 1332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1711307567
transform 1 0 1284 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1711307567
transform 1 0 2484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1711307567
transform 1 0 2100 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1711307567
transform 1 0 1732 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1711307567
transform 1 0 1372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1711307567
transform 1 0 1308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1711307567
transform 1 0 1308 0 1 2455
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1711307567
transform 1 0 2564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1711307567
transform 1 0 2332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1711307567
transform 1 0 2260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1711307567
transform 1 0 2436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1711307567
transform 1 0 2316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1711307567
transform 1 0 2756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1711307567
transform 1 0 2596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1711307567
transform 1 0 2596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1711307567
transform 1 0 2684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1711307567
transform 1 0 2588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1711307567
transform 1 0 2564 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1711307567
transform 1 0 2436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1711307567
transform 1 0 2308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1711307567
transform 1 0 2580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1711307567
transform 1 0 2516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1711307567
transform 1 0 2756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1711307567
transform 1 0 2628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1711307567
transform 1 0 2756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1711307567
transform 1 0 2628 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1711307567
transform 1 0 2124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1711307567
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1711307567
transform 1 0 2028 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1711307567
transform 1 0 2108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1711307567
transform 1 0 1996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1711307567
transform 1 0 1964 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1711307567
transform 1 0 2196 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1711307567
transform 1 0 1956 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1711307567
transform 1 0 1868 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1711307567
transform 1 0 2036 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1711307567
transform 1 0 1932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1711307567
transform 1 0 1900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1711307567
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1711307567
transform 1 0 1724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1711307567
transform 1 0 1620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1711307567
transform 1 0 1508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1711307567
transform 1 0 1452 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1711307567
transform 1 0 1420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1711307567
transform 1 0 1604 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1711307567
transform 1 0 1580 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1711307567
transform 1 0 1348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1711307567
transform 1 0 1260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1711307567
transform 1 0 1380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1711307567
transform 1 0 1212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1711307567
transform 1 0 1236 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1711307567
transform 1 0 1100 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1711307567
transform 1 0 716 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1711307567
transform 1 0 628 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1711307567
transform 1 0 860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1711307567
transform 1 0 748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1711307567
transform 1 0 900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1711307567
transform 1 0 804 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1711307567
transform 1 0 468 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1711307567
transform 1 0 420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1711307567
transform 1 0 596 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1711307567
transform 1 0 532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1711307567
transform 1 0 228 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1711307567
transform 1 0 172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1711307567
transform 1 0 348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1711307567
transform 1 0 292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1711307567
transform 1 0 188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1711307567
transform 1 0 92 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1711307567
transform 1 0 428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1711307567
transform 1 0 364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1711307567
transform 1 0 2292 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1711307567
transform 1 0 2252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1711307567
transform 1 0 2756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1711307567
transform 1 0 2660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1711307567
transform 1 0 2748 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1711307567
transform 1 0 2724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1711307567
transform 1 0 2284 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1711307567
transform 1 0 2084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1711307567
transform 1 0 2636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1711307567
transform 1 0 2316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1711307567
transform 1 0 2444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1711307567
transform 1 0 2188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1711307567
transform 1 0 2204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1711307567
transform 1 0 1932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1711307567
transform 1 0 2540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1711307567
transform 1 0 2388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1711307567
transform 1 0 2692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1711307567
transform 1 0 2516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1711307567
transform 1 0 2756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1711307567
transform 1 0 2388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1711307567
transform 1 0 1980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1711307567
transform 1 0 1852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1711307567
transform 1 0 1868 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1711307567
transform 1 0 1708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1711307567
transform 1 0 1900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1711307567
transform 1 0 1716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1711307567
transform 1 0 1860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1711307567
transform 1 0 1756 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1711307567
transform 1 0 1844 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1711307567
transform 1 0 1588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1711307567
transform 1 0 1860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1711307567
transform 1 0 1604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1711307567
transform 1 0 1476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1711307567
transform 1 0 1364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1711307567
transform 1 0 1396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1711307567
transform 1 0 1220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1711307567
transform 1 0 1732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1711307567
transform 1 0 1428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1711307567
transform 1 0 1276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1711307567
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1711307567
transform 1 0 1140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1711307567
transform 1 0 1132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1711307567
transform 1 0 1140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1711307567
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1711307567
transform 1 0 996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1711307567
transform 1 0 860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1711307567
transform 1 0 1028 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1711307567
transform 1 0 972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1711307567
transform 1 0 644 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1711307567
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1711307567
transform 1 0 764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1711307567
transform 1 0 660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1711307567
transform 1 0 732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1711307567
transform 1 0 676 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1711307567
transform 1 0 524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1711307567
transform 1 0 460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1711307567
transform 1 0 596 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1711307567
transform 1 0 380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1711307567
transform 1 0 220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1711307567
transform 1 0 188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1711307567
transform 1 0 332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1711307567
transform 1 0 308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1711307567
transform 1 0 220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1711307567
transform 1 0 188 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1711307567
transform 1 0 164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1711307567
transform 1 0 132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1711307567
transform 1 0 172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1711307567
transform 1 0 172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1711307567
transform 1 0 316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1711307567
transform 1 0 260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1711307567
transform 1 0 2164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1711307567
transform 1 0 2148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1711307567
transform 1 0 2348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1711307567
transform 1 0 2332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1711307567
transform 1 0 2228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1711307567
transform 1 0 2196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1711307567
transform 1 0 2068 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1711307567
transform 1 0 1972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1711307567
transform 1 0 2420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1711307567
transform 1 0 2332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1711307567
transform 1 0 2548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1711307567
transform 1 0 2524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1711307567
transform 1 0 2428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1711307567
transform 1 0 2428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1711307567
transform 1 0 1900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1711307567
transform 1 0 1900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1711307567
transform 1 0 1748 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1711307567
transform 1 0 1748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1711307567
transform 1 0 1700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1711307567
transform 1 0 1700 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1711307567
transform 1 0 1788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1711307567
transform 1 0 1764 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1711307567
transform 1 0 1796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1711307567
transform 1 0 1796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1711307567
transform 1 0 1620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1711307567
transform 1 0 1596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1711307567
transform 1 0 1692 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1711307567
transform 1 0 1644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1711307567
transform 1 0 1404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1711307567
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1711307567
transform 1 0 1292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1711307567
transform 1 0 1276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1711307567
transform 1 0 1468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1711307567
transform 1 0 1436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1711307567
transform 1 0 1308 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1711307567
transform 1 0 1268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1711307567
transform 1 0 1164 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1711307567
transform 1 0 1140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1711307567
transform 1 0 1124 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1711307567
transform 1 0 1124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1711307567
transform 1 0 948 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1711307567
transform 1 0 892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1711307567
transform 1 0 1020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1711307567
transform 1 0 1020 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1711307567
transform 1 0 676 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1711307567
transform 1 0 644 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1711307567
transform 1 0 756 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1711307567
transform 1 0 740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1711307567
transform 1 0 844 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1711307567
transform 1 0 708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1711307567
transform 1 0 572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1711307567
transform 1 0 532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1711307567
transform 1 0 460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1711307567
transform 1 0 420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1711307567
transform 1 0 220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1711307567
transform 1 0 212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1711307567
transform 1 0 388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1711307567
transform 1 0 348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1711307567
transform 1 0 300 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1711307567
transform 1 0 276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1711307567
transform 1 0 172 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1711307567
transform 1 0 172 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1711307567
transform 1 0 244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1711307567
transform 1 0 204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1711307567
transform 1 0 332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1711307567
transform 1 0 196 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1711307567
transform 1 0 2548 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1711307567
transform 1 0 2500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1711307567
transform 1 0 2500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1711307567
transform 1 0 2676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1711307567
transform 1 0 2644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1711307567
transform 1 0 2628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1711307567
transform 1 0 2628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1711307567
transform 1 0 2684 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1711307567
transform 1 0 2652 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1711307567
transform 1 0 2644 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1711307567
transform 1 0 2620 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1711307567
transform 1 0 2556 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1711307567
transform 1 0 2556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1711307567
transform 1 0 2516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1711307567
transform 1 0 2500 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1711307567
transform 1 0 2716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1711307567
transform 1 0 2668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1711307567
transform 1 0 2668 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1711307567
transform 1 0 2644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1711307567
transform 1 0 2604 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1711307567
transform 1 0 2500 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1711307567
transform 1 0 2476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1711307567
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1711307567
transform 1 0 2684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1711307567
transform 1 0 2604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1711307567
transform 1 0 2452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1711307567
transform 1 0 2420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1711307567
transform 1 0 2700 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1711307567
transform 1 0 2644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1711307567
transform 1 0 2612 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1711307567
transform 1 0 2460 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1711307567
transform 1 0 2372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1711307567
transform 1 0 2348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1711307567
transform 1 0 2660 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1711307567
transform 1 0 2532 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1711307567
transform 1 0 2532 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1711307567
transform 1 0 2284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1711307567
transform 1 0 2260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1711307567
transform 1 0 2596 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1711307567
transform 1 0 2532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1711307567
transform 1 0 2524 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1711307567
transform 1 0 2500 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1711307567
transform 1 0 2492 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1711307567
transform 1 0 2388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1711307567
transform 1 0 2348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1711307567
transform 1 0 2252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1711307567
transform 1 0 2252 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1711307567
transform 1 0 2708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1711307567
transform 1 0 2540 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1711307567
transform 1 0 2468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1711307567
transform 1 0 2284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1711307567
transform 1 0 2244 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1711307567
transform 1 0 2756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1711307567
transform 1 0 2596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1711307567
transform 1 0 2572 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1711307567
transform 1 0 2516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1711307567
transform 1 0 2484 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1711307567
transform 1 0 2356 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1711307567
transform 1 0 2284 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1711307567
transform 1 0 2252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1711307567
transform 1 0 2756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1711307567
transform 1 0 2668 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1711307567
transform 1 0 2628 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1711307567
transform 1 0 2628 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1711307567
transform 1 0 2620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1711307567
transform 1 0 2612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1711307567
transform 1 0 2604 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1711307567
transform 1 0 2620 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1711307567
transform 1 0 2596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1711307567
transform 1 0 2756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1711307567
transform 1 0 2644 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1711307567
transform 1 0 2380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1711307567
transform 1 0 2332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1711307567
transform 1 0 2308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1711307567
transform 1 0 1876 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1711307567
transform 1 0 1852 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1711307567
transform 1 0 1780 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1711307567
transform 1 0 1668 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1711307567
transform 1 0 1644 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1711307567
transform 1 0 1588 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1711307567
transform 1 0 1548 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1711307567
transform 1 0 1188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1711307567
transform 1 0 1164 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1711307567
transform 1 0 540 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1711307567
transform 1 0 532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1711307567
transform 1 0 492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1711307567
transform 1 0 1028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1711307567
transform 1 0 980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1711307567
transform 1 0 820 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1711307567
transform 1 0 812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1711307567
transform 1 0 788 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1711307567
transform 1 0 764 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1711307567
transform 1 0 764 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1711307567
transform 1 0 748 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1711307567
transform 1 0 668 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1711307567
transform 1 0 660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1711307567
transform 1 0 524 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1711307567
transform 1 0 524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1711307567
transform 1 0 1532 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1711307567
transform 1 0 1500 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1711307567
transform 1 0 1484 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1711307567
transform 1 0 1428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1711307567
transform 1 0 1924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1711307567
transform 1 0 1868 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1711307567
transform 1 0 1868 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1711307567
transform 1 0 1836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1711307567
transform 1 0 1828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1711307567
transform 1 0 1644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1711307567
transform 1 0 860 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1711307567
transform 1 0 836 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1711307567
transform 1 0 2060 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1711307567
transform 1 0 2036 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1711307567
transform 1 0 1932 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1711307567
transform 1 0 1860 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1711307567
transform 1 0 1828 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1711307567
transform 1 0 1972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1711307567
transform 1 0 1892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1711307567
transform 1 0 1892 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1711307567
transform 1 0 1820 0 1 2485
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1711307567
transform 1 0 1820 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1711307567
transform 1 0 1892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1711307567
transform 1 0 1812 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1711307567
transform 1 0 1676 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1711307567
transform 1 0 1676 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1711307567
transform 1 0 996 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1711307567
transform 1 0 780 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1711307567
transform 1 0 956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1711307567
transform 1 0 908 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1711307567
transform 1 0 908 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1711307567
transform 1 0 884 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1711307567
transform 1 0 1932 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1711307567
transform 1 0 1508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1711307567
transform 1 0 1436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1711307567
transform 1 0 836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1711307567
transform 1 0 1676 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1711307567
transform 1 0 1660 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1711307567
transform 1 0 1412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1711307567
transform 1 0 1076 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1711307567
transform 1 0 524 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1711307567
transform 1 0 356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1711307567
transform 1 0 340 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1711307567
transform 1 0 1052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1711307567
transform 1 0 1028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1711307567
transform 1 0 860 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1711307567
transform 1 0 772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1711307567
transform 1 0 1924 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1711307567
transform 1 0 1788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1711307567
transform 1 0 1748 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1711307567
transform 1 0 1268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1711307567
transform 1 0 1252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1711307567
transform 1 0 932 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1711307567
transform 1 0 908 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1711307567
transform 1 0 1516 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1711307567
transform 1 0 1436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1711307567
transform 1 0 1388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1711307567
transform 1 0 1332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1711307567
transform 1 0 1300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1711307567
transform 1 0 1916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1711307567
transform 1 0 1844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1711307567
transform 1 0 1516 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1711307567
transform 1 0 1316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1711307567
transform 1 0 1228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1711307567
transform 1 0 1644 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1711307567
transform 1 0 1628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1711307567
transform 1 0 1612 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1711307567
transform 1 0 1604 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1711307567
transform 1 0 564 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1711307567
transform 1 0 380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1711307567
transform 1 0 356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1711307567
transform 1 0 316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1711307567
transform 1 0 1676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1711307567
transform 1 0 1660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1711307567
transform 1 0 1620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1711307567
transform 1 0 1612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1711307567
transform 1 0 1596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1711307567
transform 1 0 1572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1711307567
transform 1 0 1332 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1711307567
transform 1 0 1132 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1711307567
transform 1 0 1076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1711307567
transform 1 0 1044 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1711307567
transform 1 0 1604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1711307567
transform 1 0 1572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1711307567
transform 1 0 628 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1711307567
transform 1 0 484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1711307567
transform 1 0 1796 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1711307567
transform 1 0 1796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1711307567
transform 1 0 1748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1711307567
transform 1 0 1716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1711307567
transform 1 0 1460 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1711307567
transform 1 0 1388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1711307567
transform 1 0 1860 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1711307567
transform 1 0 1860 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1711307567
transform 1 0 1860 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1711307567
transform 1 0 1828 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1711307567
transform 1 0 1388 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1711307567
transform 1 0 988 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1711307567
transform 1 0 548 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1711307567
transform 1 0 412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1711307567
transform 1 0 388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1711307567
transform 1 0 572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1711307567
transform 1 0 532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1711307567
transform 1 0 484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1711307567
transform 1 0 468 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1711307567
transform 1 0 1156 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1711307567
transform 1 0 1156 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1711307567
transform 1 0 1108 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1711307567
transform 1 0 908 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1711307567
transform 1 0 884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1711307567
transform 1 0 2028 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1711307567
transform 1 0 1748 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1711307567
transform 1 0 1420 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1711307567
transform 1 0 1388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1711307567
transform 1 0 1084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1711307567
transform 1 0 1356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1711307567
transform 1 0 1148 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1711307567
transform 1 0 1060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1711307567
transform 1 0 1692 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1711307567
transform 1 0 1588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1711307567
transform 1 0 1236 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1711307567
transform 1 0 780 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1711307567
transform 1 0 524 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1711307567
transform 1 0 836 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1711307567
transform 1 0 796 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1711307567
transform 1 0 780 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1711307567
transform 1 0 772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1711307567
transform 1 0 748 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1711307567
transform 1 0 748 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1711307567
transform 1 0 2116 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1711307567
transform 1 0 2044 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1711307567
transform 1 0 1988 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1711307567
transform 1 0 1252 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1711307567
transform 1 0 1212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1711307567
transform 1 0 1052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1711307567
transform 1 0 1004 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1711307567
transform 1 0 980 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1711307567
transform 1 0 1716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1711307567
transform 1 0 1676 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1711307567
transform 1 0 804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1711307567
transform 1 0 636 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1711307567
transform 1 0 516 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1711307567
transform 1 0 508 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1711307567
transform 1 0 1788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1711307567
transform 1 0 1716 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1711307567
transform 1 0 1900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1711307567
transform 1 0 1876 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1711307567
transform 1 0 2084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1711307567
transform 1 0 2060 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1711307567
transform 1 0 2012 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1711307567
transform 1 0 1732 0 1 1895
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1711307567
transform 1 0 1724 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1711307567
transform 1 0 1692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1711307567
transform 1 0 1596 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1711307567
transform 1 0 1260 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1711307567
transform 1 0 1188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1711307567
transform 1 0 1172 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1711307567
transform 1 0 1172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1711307567
transform 1 0 732 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1711307567
transform 1 0 708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1711307567
transform 1 0 628 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1711307567
transform 1 0 628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1711307567
transform 1 0 596 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1711307567
transform 1 0 588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1711307567
transform 1 0 548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1711307567
transform 1 0 2060 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1711307567
transform 1 0 2044 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1711307567
transform 1 0 1140 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1711307567
transform 1 0 1124 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1711307567
transform 1 0 988 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1711307567
transform 1 0 812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1711307567
transform 1 0 812 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1711307567
transform 1 0 772 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1711307567
transform 1 0 764 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1711307567
transform 1 0 764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1711307567
transform 1 0 2020 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1711307567
transform 1 0 2020 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1711307567
transform 1 0 1980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1711307567
transform 1 0 1876 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1711307567
transform 1 0 1876 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1711307567
transform 1 0 2332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1711307567
transform 1 0 2332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1711307567
transform 1 0 2308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1711307567
transform 1 0 2268 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1711307567
transform 1 0 2228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1711307567
transform 1 0 2388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1711307567
transform 1 0 2380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1711307567
transform 1 0 2300 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1711307567
transform 1 0 2292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1711307567
transform 1 0 2220 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1711307567
transform 1 0 1108 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1711307567
transform 1 0 1020 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1711307567
transform 1 0 956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1711307567
transform 1 0 1740 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1711307567
transform 1 0 1692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1711307567
transform 1 0 2252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1711307567
transform 1 0 2036 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1711307567
transform 1 0 2036 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1711307567
transform 1 0 1188 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1711307567
transform 1 0 820 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1711307567
transform 1 0 572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1711307567
transform 1 0 2172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1711307567
transform 1 0 2004 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1711307567
transform 1 0 1684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1711307567
transform 1 0 1140 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1711307567
transform 1 0 604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1711307567
transform 1 0 1892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1711307567
transform 1 0 1796 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1711307567
transform 1 0 1220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1711307567
transform 1 0 820 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1711307567
transform 1 0 1700 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1711307567
transform 1 0 1668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1711307567
transform 1 0 2364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1711307567
transform 1 0 2356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1711307567
transform 1 0 2284 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1711307567
transform 1 0 2252 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1711307567
transform 1 0 2236 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1711307567
transform 1 0 2092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1711307567
transform 1 0 1916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1711307567
transform 1 0 1708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1711307567
transform 1 0 844 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1711307567
transform 1 0 716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1711307567
transform 1 0 1668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1711307567
transform 1 0 1628 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1711307567
transform 1 0 1964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1711307567
transform 1 0 1892 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1711307567
transform 1 0 1188 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1711307567
transform 1 0 852 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1711307567
transform 1 0 2276 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1711307567
transform 1 0 2036 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1711307567
transform 1 0 1228 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1711307567
transform 1 0 788 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1711307567
transform 1 0 596 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1711307567
transform 1 0 980 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1711307567
transform 1 0 892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1711307567
transform 1 0 892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1711307567
transform 1 0 1604 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1711307567
transform 1 0 1492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1711307567
transform 1 0 1476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1711307567
transform 1 0 2076 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1711307567
transform 1 0 2076 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1711307567
transform 1 0 1684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1711307567
transform 1 0 1084 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1711307567
transform 1 0 700 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1711307567
transform 1 0 2524 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1711307567
transform 1 0 2508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1711307567
transform 1 0 2628 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1711307567
transform 1 0 2628 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1711307567
transform 1 0 2596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1711307567
transform 1 0 2572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1711307567
transform 1 0 2668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1711307567
transform 1 0 2636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1711307567
transform 1 0 2612 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1711307567
transform 1 0 2580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1711307567
transform 1 0 2644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1711307567
transform 1 0 2628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1711307567
transform 1 0 2596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1711307567
transform 1 0 2572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1711307567
transform 1 0 2636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1711307567
transform 1 0 2636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1711307567
transform 1 0 2724 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1711307567
transform 1 0 2724 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1711307567
transform 1 0 2700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1711307567
transform 1 0 2700 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1711307567
transform 1 0 2740 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1711307567
transform 1 0 2652 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1711307567
transform 1 0 2572 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1711307567
transform 1 0 2556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1711307567
transform 1 0 2524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1711307567
transform 1 0 204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1711307567
transform 1 0 204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1711307567
transform 1 0 196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1711307567
transform 1 0 124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1711307567
transform 1 0 100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1711307567
transform 1 0 236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1711307567
transform 1 0 236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1711307567
transform 1 0 268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1711307567
transform 1 0 268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1711307567
transform 1 0 188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1711307567
transform 1 0 188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1711307567
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1711307567
transform 1 0 548 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1711307567
transform 1 0 436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1711307567
transform 1 0 436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1711307567
transform 1 0 756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1711307567
transform 1 0 748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1711307567
transform 1 0 748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1711307567
transform 1 0 644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1711307567
transform 1 0 644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1711307567
transform 1 0 1068 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1711307567
transform 1 0 1028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1711307567
transform 1 0 972 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1711307567
transform 1 0 1068 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1711307567
transform 1 0 1060 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1711307567
transform 1 0 1004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1711307567
transform 1 0 1108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1711307567
transform 1 0 1108 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1711307567
transform 1 0 1180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1711307567
transform 1 0 1156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1711307567
transform 1 0 1612 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1711307567
transform 1 0 1604 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1711307567
transform 1 0 1516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1711307567
transform 1 0 1484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1711307567
transform 1 0 1740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1711307567
transform 1 0 1732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1711307567
transform 1 0 2084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1711307567
transform 1 0 2084 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1711307567
transform 1 0 2708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1711307567
transform 1 0 2644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1711307567
transform 1 0 2612 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1711307567
transform 1 0 2652 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1711307567
transform 1 0 2644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1711307567
transform 1 0 2604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1711307567
transform 1 0 2540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1711307567
transform 1 0 2524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1711307567
transform 1 0 2468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1711307567
transform 1 0 2316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1711307567
transform 1 0 2284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1711307567
transform 1 0 2284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1711307567
transform 1 0 2532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1711307567
transform 1 0 2516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1711307567
transform 1 0 2604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1711307567
transform 1 0 2604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1711307567
transform 1 0 2332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1711307567
transform 1 0 2324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1711307567
transform 1 0 2292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1711307567
transform 1 0 2316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1711307567
transform 1 0 2284 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1711307567
transform 1 0 2580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1711307567
transform 1 0 2436 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1711307567
transform 1 0 2428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1711307567
transform 1 0 2596 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1711307567
transform 1 0 2556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1711307567
transform 1 0 2548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1711307567
transform 1 0 2428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1711307567
transform 1 0 2524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1711307567
transform 1 0 2508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1711307567
transform 1 0 2508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1711307567
transform 1 0 2516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1711307567
transform 1 0 2492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1711307567
transform 1 0 2468 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1711307567
transform 1 0 2436 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1711307567
transform 1 0 2540 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1711307567
transform 1 0 2516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1711307567
transform 1 0 2468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1711307567
transform 1 0 2580 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1711307567
transform 1 0 2532 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1711307567
transform 1 0 2476 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1711307567
transform 1 0 2476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1711307567
transform 1 0 2476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1711307567
transform 1 0 1628 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1711307567
transform 1 0 1260 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1711307567
transform 1 0 1580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1711307567
transform 1 0 1540 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1711307567
transform 1 0 1508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1711307567
transform 1 0 1204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1711307567
transform 1 0 1820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1711307567
transform 1 0 1788 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1711307567
transform 1 0 1716 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1711307567
transform 1 0 1980 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1711307567
transform 1 0 1964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1711307567
transform 1 0 1900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1711307567
transform 1 0 1900 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1711307567
transform 1 0 2020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1711307567
transform 1 0 2012 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1711307567
transform 1 0 1884 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1711307567
transform 1 0 1868 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1711307567
transform 1 0 1860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1711307567
transform 1 0 1828 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1711307567
transform 1 0 1868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1711307567
transform 1 0 1844 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1711307567
transform 1 0 1772 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1711307567
transform 1 0 1764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1711307567
transform 1 0 1852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1711307567
transform 1 0 1716 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1711307567
transform 1 0 1660 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1711307567
transform 1 0 1652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1711307567
transform 1 0 1540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1711307567
transform 1 0 1484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1711307567
transform 1 0 332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1711307567
transform 1 0 308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1711307567
transform 1 0 228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1711307567
transform 1 0 212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1711307567
transform 1 0 364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1711307567
transform 1 0 220 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1711307567
transform 1 0 828 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1711307567
transform 1 0 668 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1711307567
transform 1 0 372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1711307567
transform 1 0 364 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1711307567
transform 1 0 316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1711307567
transform 1 0 308 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1711307567
transform 1 0 268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1711307567
transform 1 0 268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1711307567
transform 1 0 484 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1711307567
transform 1 0 348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1711307567
transform 1 0 332 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1711307567
transform 1 0 292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1711307567
transform 1 0 420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1711307567
transform 1 0 380 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1711307567
transform 1 0 364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1711307567
transform 1 0 668 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1711307567
transform 1 0 580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1711307567
transform 1 0 548 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1711307567
transform 1 0 604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1711307567
transform 1 0 524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1711307567
transform 1 0 508 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1711307567
transform 1 0 364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1711307567
transform 1 0 684 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1711307567
transform 1 0 524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1711307567
transform 1 0 508 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1711307567
transform 1 0 428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1711307567
transform 1 0 412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1711307567
transform 1 0 660 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1711307567
transform 1 0 628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1711307567
transform 1 0 604 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1711307567
transform 1 0 604 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1711307567
transform 1 0 324 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1711307567
transform 1 0 308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1711307567
transform 1 0 764 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1711307567
transform 1 0 740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1711307567
transform 1 0 692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1711307567
transform 1 0 660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1711307567
transform 1 0 636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1711307567
transform 1 0 636 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1711307567
transform 1 0 1372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1711307567
transform 1 0 796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1711307567
transform 1 0 772 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1711307567
transform 1 0 660 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1711307567
transform 1 0 1300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1711307567
transform 1 0 828 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1711307567
transform 1 0 860 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1711307567
transform 1 0 732 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1711307567
transform 1 0 732 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1711307567
transform 1 0 724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1711307567
transform 1 0 652 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1711307567
transform 1 0 572 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1711307567
transform 1 0 516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1711307567
transform 1 0 836 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1711307567
transform 1 0 804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1711307567
transform 1 0 724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1711307567
transform 1 0 676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1711307567
transform 1 0 636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1711307567
transform 1 0 636 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1711307567
transform 1 0 636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1711307567
transform 1 0 692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1711307567
transform 1 0 692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1711307567
transform 1 0 644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1711307567
transform 1 0 644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1711307567
transform 1 0 612 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1711307567
transform 1 0 604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1711307567
transform 1 0 564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1711307567
transform 1 0 564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1711307567
transform 1 0 1676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1711307567
transform 1 0 1652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1711307567
transform 1 0 1628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1711307567
transform 1 0 1388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1711307567
transform 1 0 1028 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1711307567
transform 1 0 1004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1711307567
transform 1 0 836 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1711307567
transform 1 0 508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1711307567
transform 1 0 508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1711307567
transform 1 0 468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1711307567
transform 1 0 396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1711307567
transform 1 0 396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1711307567
transform 1 0 2228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1711307567
transform 1 0 2212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1711307567
transform 1 0 2180 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1711307567
transform 1 0 2140 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1711307567
transform 1 0 1412 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1711307567
transform 1 0 1116 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1711307567
transform 1 0 1108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1711307567
transform 1 0 1492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1711307567
transform 1 0 1004 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1711307567
transform 1 0 852 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1711307567
transform 1 0 804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1711307567
transform 1 0 1356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1711307567
transform 1 0 1108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1711307567
transform 1 0 1100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1711307567
transform 1 0 1092 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1711307567
transform 1 0 1092 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1711307567
transform 1 0 1276 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1711307567
transform 1 0 1140 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1711307567
transform 1 0 1108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1711307567
transform 1 0 1236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1711307567
transform 1 0 1148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1711307567
transform 1 0 996 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1711307567
transform 1 0 868 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1711307567
transform 1 0 684 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1711307567
transform 1 0 684 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1711307567
transform 1 0 868 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1711307567
transform 1 0 860 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1711307567
transform 1 0 1212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1711307567
transform 1 0 1140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1711307567
transform 1 0 1076 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1711307567
transform 1 0 996 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1711307567
transform 1 0 1100 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1711307567
transform 1 0 980 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1711307567
transform 1 0 876 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1711307567
transform 1 0 804 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1711307567
transform 1 0 764 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1711307567
transform 1 0 1132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1711307567
transform 1 0 1124 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1711307567
transform 1 0 1084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1711307567
transform 1 0 1476 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1711307567
transform 1 0 1476 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1711307567
transform 1 0 980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1711307567
transform 1 0 980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1711307567
transform 1 0 956 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1711307567
transform 1 0 956 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1711307567
transform 1 0 828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1711307567
transform 1 0 828 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1711307567
transform 1 0 1164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1711307567
transform 1 0 1164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1711307567
transform 1 0 1132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1711307567
transform 1 0 1108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1711307567
transform 1 0 1492 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1711307567
transform 1 0 1364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1711307567
transform 1 0 1548 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1711307567
transform 1 0 1316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1711307567
transform 1 0 1252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1711307567
transform 1 0 1212 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1711307567
transform 1 0 1148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1711307567
transform 1 0 1148 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1711307567
transform 1 0 1860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1711307567
transform 1 0 1804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1711307567
transform 1 0 1796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1711307567
transform 1 0 1460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1711307567
transform 1 0 1436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1711307567
transform 1 0 1452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1711307567
transform 1 0 1332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1711307567
transform 1 0 1532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1711307567
transform 1 0 1516 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1711307567
transform 1 0 1492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1711307567
transform 1 0 1484 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1711307567
transform 1 0 1452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1711307567
transform 1 0 1836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1711307567
transform 1 0 1756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1711307567
transform 1 0 1612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1711307567
transform 1 0 1532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1711307567
transform 1 0 2196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1711307567
transform 1 0 2164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1711307567
transform 1 0 2124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1711307567
transform 1 0 2124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1711307567
transform 1 0 1580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1711307567
transform 1 0 1580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1711307567
transform 1 0 1516 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1711307567
transform 1 0 1412 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1711307567
transform 1 0 1412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1711307567
transform 1 0 1388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1711307567
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1711307567
transform 1 0 2500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1711307567
transform 1 0 2500 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1711307567
transform 1 0 2452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1711307567
transform 1 0 2436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1711307567
transform 1 0 1908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1711307567
transform 1 0 1740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1711307567
transform 1 0 1540 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1711307567
transform 1 0 1548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1711307567
transform 1 0 1372 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1711307567
transform 1 0 1332 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1711307567
transform 1 0 1324 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1711307567
transform 1 0 2620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1711307567
transform 1 0 2604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1711307567
transform 1 0 2580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1711307567
transform 1 0 2580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1711307567
transform 1 0 1916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1711307567
transform 1 0 1540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1711307567
transform 1 0 2116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1711307567
transform 1 0 2108 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1711307567
transform 1 0 2740 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1711307567
transform 1 0 2668 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1711307567
transform 1 0 2748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1711307567
transform 1 0 2732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1711307567
transform 1 0 2644 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1711307567
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1711307567
transform 1 0 2556 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1711307567
transform 1 0 2692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1711307567
transform 1 0 2612 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1711307567
transform 1 0 2732 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1711307567
transform 1 0 2692 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1711307567
transform 1 0 2668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1711307567
transform 1 0 2644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1711307567
transform 1 0 2540 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1711307567
transform 1 0 2668 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1711307567
transform 1 0 2644 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1711307567
transform 1 0 2620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1711307567
transform 1 0 2548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1711307567
transform 1 0 2692 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1711307567
transform 1 0 2564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1711307567
transform 1 0 2516 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1711307567
transform 1 0 2572 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1711307567
transform 1 0 2564 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1711307567
transform 1 0 2548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1711307567
transform 1 0 2548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1711307567
transform 1 0 2500 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1711307567
transform 1 0 2500 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1711307567
transform 1 0 1460 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1711307567
transform 1 0 1452 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1711307567
transform 1 0 148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1711307567
transform 1 0 148 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1711307567
transform 1 0 140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1711307567
transform 1 0 140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1711307567
transform 1 0 140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1711307567
transform 1 0 140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1711307567
transform 1 0 2028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1711307567
transform 1 0 2028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1711307567
transform 1 0 2212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1711307567
transform 1 0 2140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1711307567
transform 1 0 2292 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1711307567
transform 1 0 2292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1711307567
transform 1 0 2108 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1711307567
transform 1 0 2108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1711307567
transform 1 0 2740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1711307567
transform 1 0 2732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1711307567
transform 1 0 2724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1711307567
transform 1 0 2756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1711307567
transform 1 0 2700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1711307567
transform 1 0 2684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1711307567
transform 1 0 2756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1711307567
transform 1 0 2724 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1711307567
transform 1 0 2732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1711307567
transform 1 0 2676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1711307567
transform 1 0 2156 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1711307567
transform 1 0 2116 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1711307567
transform 1 0 2028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1711307567
transform 1 0 2028 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1711307567
transform 1 0 1980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1711307567
transform 1 0 1956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1711307567
transform 1 0 1636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1711307567
transform 1 0 1540 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1711307567
transform 1 0 1476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1711307567
transform 1 0 1372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1711307567
transform 1 0 1292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1711307567
transform 1 0 1268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1711307567
transform 1 0 1156 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1711307567
transform 1 0 2700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1711307567
transform 1 0 2676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1711307567
transform 1 0 932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1711307567
transform 1 0 932 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1711307567
transform 1 0 812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1711307567
transform 1 0 780 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1711307567
transform 1 0 636 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1711307567
transform 1 0 516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1711307567
transform 1 0 388 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1711307567
transform 1 0 348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1711307567
transform 1 0 268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1711307567
transform 1 0 148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1711307567
transform 1 0 92 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1711307567
transform 1 0 92 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1711307567
transform 1 0 84 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1711307567
transform 1 0 2708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1711307567
transform 1 0 2668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1711307567
transform 1 0 2660 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1711307567
transform 1 0 2572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1711307567
transform 1 0 2484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1711307567
transform 1 0 2484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1711307567
transform 1 0 2476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1711307567
transform 1 0 2460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1711307567
transform 1 0 2452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1711307567
transform 1 0 2436 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1711307567
transform 1 0 2404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1711307567
transform 1 0 2372 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1711307567
transform 1 0 2364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1711307567
transform 1 0 2308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1711307567
transform 1 0 2244 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1711307567
transform 1 0 2212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1711307567
transform 1 0 2676 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1711307567
transform 1 0 2676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1711307567
transform 1 0 2620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1711307567
transform 1 0 2612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1711307567
transform 1 0 2556 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1711307567
transform 1 0 2460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1711307567
transform 1 0 2460 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1711307567
transform 1 0 2364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1711307567
transform 1 0 2324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1711307567
transform 1 0 2268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1711307567
transform 1 0 2204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1711307567
transform 1 0 2124 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1711307567
transform 1 0 2068 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1711307567
transform 1 0 1900 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1711307567
transform 1 0 1820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1711307567
transform 1 0 1788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1711307567
transform 1 0 1780 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1711307567
transform 1 0 1780 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1711307567
transform 1 0 1748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1711307567
transform 1 0 1652 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1711307567
transform 1 0 1564 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1711307567
transform 1 0 1396 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1711307567
transform 1 0 1316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1711307567
transform 1 0 1196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1711307567
transform 1 0 1060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1711307567
transform 1 0 1060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1711307567
transform 1 0 860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1711307567
transform 1 0 1484 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1711307567
transform 1 0 1436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1711307567
transform 1 0 948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1711307567
transform 1 0 684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1711307567
transform 1 0 636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1711307567
transform 1 0 564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1711307567
transform 1 0 516 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1711307567
transform 1 0 444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1711307567
transform 1 0 244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1711307567
transform 1 0 236 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1711307567
transform 1 0 140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1711307567
transform 1 0 140 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1711307567
transform 1 0 84 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1711307567
transform 1 0 84 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1711307567
transform 1 0 2444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1711307567
transform 1 0 2348 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1711307567
transform 1 0 2252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1711307567
transform 1 0 2196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1711307567
transform 1 0 2108 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1711307567
transform 1 0 2084 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1711307567
transform 1 0 1988 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1711307567
transform 1 0 1820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1711307567
transform 1 0 1716 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1711307567
transform 1 0 1708 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1711307567
transform 1 0 1620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1711307567
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1711307567
transform 1 0 1572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1711307567
transform 1 0 1508 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1711307567
transform 1 0 1436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1711307567
transform 1 0 1356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1711307567
transform 1 0 1316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1711307567
transform 1 0 1228 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1711307567
transform 1 0 1156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1711307567
transform 1 0 1060 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1711307567
transform 1 0 1020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1711307567
transform 1 0 940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1711307567
transform 1 0 852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1711307567
transform 1 0 764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1711307567
transform 1 0 676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1711307567
transform 1 0 596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1711307567
transform 1 0 484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1711307567
transform 1 0 380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1711307567
transform 1 0 2540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1711307567
transform 1 0 2476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1711307567
transform 1 0 2420 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1711307567
transform 1 0 2372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1711307567
transform 1 0 2324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1711307567
transform 1 0 2292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1711307567
transform 1 0 2204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1711307567
transform 1 0 1476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1711307567
transform 1 0 308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1711307567
transform 1 0 220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1711307567
transform 1 0 132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1711307567
transform 1 0 108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1711307567
transform 1 0 92 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1711307567
transform 1 0 92 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1711307567
transform 1 0 2028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1711307567
transform 1 0 1532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1711307567
transform 1 0 1516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1711307567
transform 1 0 1460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1711307567
transform 1 0 1524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1711307567
transform 1 0 1492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1711307567
transform 1 0 1436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1711307567
transform 1 0 1420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1711307567
transform 1 0 2548 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1711307567
transform 1 0 2452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1711307567
transform 1 0 2396 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1711307567
transform 1 0 2356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1711307567
transform 1 0 2292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1711307567
transform 1 0 2284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1711307567
transform 1 0 2284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1711307567
transform 1 0 2276 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1711307567
transform 1 0 2228 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1711307567
transform 1 0 2140 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1711307567
transform 1 0 2092 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1711307567
transform 1 0 2012 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1711307567
transform 1 0 1764 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1711307567
transform 1 0 1444 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1711307567
transform 1 0 204 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1711307567
transform 1 0 188 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1711307567
transform 1 0 172 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1711307567
transform 1 0 2652 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1711307567
transform 1 0 2628 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1711307567
transform 1 0 2596 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1711307567
transform 1 0 2580 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1711307567
transform 1 0 2508 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1711307567
transform 1 0 2492 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1711307567
transform 1 0 2468 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1711307567
transform 1 0 2468 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1711307567
transform 1 0 2372 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1711307567
transform 1 0 2364 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1711307567
transform 1 0 2356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1711307567
transform 1 0 2356 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1711307567
transform 1 0 2324 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1711307567
transform 1 0 2292 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1711307567
transform 1 0 2252 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1711307567
transform 1 0 2196 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1711307567
transform 1 0 2172 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1711307567
transform 1 0 2060 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1711307567
transform 1 0 2004 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1711307567
transform 1 0 2116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1711307567
transform 1 0 2052 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1711307567
transform 1 0 1940 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1711307567
transform 1 0 1852 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1711307567
transform 1 0 1844 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1711307567
transform 1 0 1724 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1711307567
transform 1 0 1564 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1711307567
transform 1 0 1436 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1711307567
transform 1 0 1332 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1711307567
transform 1 0 1172 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1711307567
transform 1 0 1084 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1711307567
transform 1 0 1068 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1711307567
transform 1 0 1060 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1711307567
transform 1 0 1052 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1711307567
transform 1 0 1044 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1711307567
transform 1 0 2396 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1711307567
transform 1 0 2380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1711307567
transform 1 0 2364 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1711307567
transform 1 0 772 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1711307567
transform 1 0 692 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1711307567
transform 1 0 604 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1711307567
transform 1 0 500 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1711307567
transform 1 0 396 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1711307567
transform 1 0 388 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1711307567
transform 1 0 308 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1711307567
transform 1 0 188 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1711307567
transform 1 0 172 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1711307567
transform 1 0 172 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1711307567
transform 1 0 164 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1711307567
transform 1 0 132 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1711307567
transform 1 0 108 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1711307567
transform 1 0 1940 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1711307567
transform 1 0 1740 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1711307567
transform 1 0 1732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1711307567
transform 1 0 1652 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1711307567
transform 1 0 1556 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1711307567
transform 1 0 1548 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1711307567
transform 1 0 1228 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1711307567
transform 1 0 1044 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1711307567
transform 1 0 924 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1711307567
transform 1 0 844 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1711307567
transform 1 0 476 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1711307567
transform 1 0 428 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1711307567
transform 1 0 396 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1711307567
transform 1 0 2300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1711307567
transform 1 0 2292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1711307567
transform 1 0 2236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1711307567
transform 1 0 2220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1711307567
transform 1 0 1892 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1711307567
transform 1 0 1612 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1711307567
transform 1 0 1380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1711307567
transform 1 0 1356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1711307567
transform 1 0 1164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1711307567
transform 1 0 980 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1711307567
transform 1 0 804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1711307567
transform 1 0 708 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1711307567
transform 1 0 636 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1711307567
transform 1 0 340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1711307567
transform 1 0 2620 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1711307567
transform 1 0 2300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1711307567
transform 1 0 2268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1711307567
transform 1 0 2268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1711307567
transform 1 0 2212 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1711307567
transform 1 0 2212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1711307567
transform 1 0 2172 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1711307567
transform 1 0 2140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1711307567
transform 1 0 2132 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1711307567
transform 1 0 2116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1711307567
transform 1 0 2076 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1711307567
transform 1 0 2044 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1711307567
transform 1 0 2044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1711307567
transform 1 0 1852 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1711307567
transform 1 0 1812 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1711307567
transform 1 0 1796 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1711307567
transform 1 0 1380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1711307567
transform 1 0 1364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1711307567
transform 1 0 1300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1711307567
transform 1 0 1132 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1711307567
transform 1 0 1068 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1711307567
transform 1 0 916 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1711307567
transform 1 0 756 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1711307567
transform 1 0 668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1711307567
transform 1 0 652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1711307567
transform 1 0 468 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1711307567
transform 1 0 388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1711307567
transform 1 0 220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1711307567
transform 1 0 196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1711307567
transform 1 0 196 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1711307567
transform 1 0 2020 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1711307567
transform 1 0 1996 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1711307567
transform 1 0 1956 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1711307567
transform 1 0 1932 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1711307567
transform 1 0 1876 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1711307567
transform 1 0 1828 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1711307567
transform 1 0 1660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1711307567
transform 1 0 2044 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1711307567
transform 1 0 1924 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1711307567
transform 1 0 1852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1711307567
transform 1 0 1772 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1711307567
transform 1 0 1676 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1711307567
transform 1 0 1580 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1711307567
transform 1 0 1572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1711307567
transform 1 0 1420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1711307567
transform 1 0 1380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1711307567
transform 1 0 1212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1711307567
transform 1 0 1204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1711307567
transform 1 0 1140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1711307567
transform 1 0 2308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1711307567
transform 1 0 2012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1711307567
transform 1 0 1012 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1711307567
transform 1 0 940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1711307567
transform 1 0 860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1711307567
transform 1 0 636 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1711307567
transform 1 0 636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1711307567
transform 1 0 596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1711307567
transform 1 0 2196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1711307567
transform 1 0 1956 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1711307567
transform 1 0 420 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1711307567
transform 1 0 340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1711307567
transform 1 0 300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1711307567
transform 1 0 220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1711307567
transform 1 0 196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1711307567
transform 1 0 140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1711307567
transform 1 0 1940 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1711307567
transform 1 0 1844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1711307567
transform 1 0 244 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1711307567
transform 1 0 220 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1711307567
transform 1 0 2492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1711307567
transform 1 0 2364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1711307567
transform 1 0 2348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1711307567
transform 1 0 2116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1711307567
transform 1 0 2036 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1711307567
transform 1 0 1868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1711307567
transform 1 0 1860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1711307567
transform 1 0 1804 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1711307567
transform 1 0 1724 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1711307567
transform 1 0 1716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1711307567
transform 1 0 2212 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1711307567
transform 1 0 2164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1711307567
transform 1 0 2108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1711307567
transform 1 0 1956 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1711307567
transform 1 0 1812 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1711307567
transform 1 0 1628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1711307567
transform 1 0 1628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1711307567
transform 1 0 1452 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1711307567
transform 1 0 1396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1711307567
transform 1 0 1268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1711307567
transform 1 0 1260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1711307567
transform 1 0 700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1711307567
transform 1 0 684 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1711307567
transform 1 0 612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1711307567
transform 1 0 484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1711307567
transform 1 0 404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1711307567
transform 1 0 332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1711307567
transform 1 0 316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1711307567
transform 1 0 292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1711307567
transform 1 0 236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1711307567
transform 1 0 236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1711307567
transform 1 0 188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1711307567
transform 1 0 2172 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1711307567
transform 1 0 2164 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1711307567
transform 1 0 2132 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1711307567
transform 1 0 2108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1711307567
transform 1 0 2076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1711307567
transform 1 0 1988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1711307567
transform 1 0 1836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1711307567
transform 1 0 1740 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1711307567
transform 1 0 1708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1711307567
transform 1 0 1500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1711307567
transform 1 0 1420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1711307567
transform 1 0 1316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1711307567
transform 1 0 1276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1711307567
transform 1 0 1276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1711307567
transform 1 0 1084 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1711307567
transform 1 0 1068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1711307567
transform 1 0 1052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1711307567
transform 1 0 996 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1711307567
transform 1 0 996 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1711307567
transform 1 0 852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1711307567
transform 1 0 764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1711307567
transform 1 0 716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1711307567
transform 1 0 692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1711307567
transform 1 0 588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1711307567
transform 1 0 492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1711307567
transform 1 0 316 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1711307567
transform 1 0 316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1711307567
transform 1 0 276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1711307567
transform 1 0 276 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1711307567
transform 1 0 2068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1711307567
transform 1 0 2060 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1711307567
transform 1 0 2028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1711307567
transform 1 0 1996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1711307567
transform 1 0 1924 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1711307567
transform 1 0 1908 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1711307567
transform 1 0 1836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1711307567
transform 1 0 1636 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1711307567
transform 1 0 1572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1711307567
transform 1 0 1020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1711307567
transform 1 0 924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1711307567
transform 1 0 468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1711307567
transform 1 0 460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1711307567
transform 1 0 2012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1711307567
transform 1 0 1996 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1711307567
transform 1 0 1972 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1711307567
transform 1 0 1940 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1711307567
transform 1 0 1932 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1711307567
transform 1 0 1884 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1711307567
transform 1 0 1812 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1711307567
transform 1 0 1804 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1711307567
transform 1 0 1796 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1711307567
transform 1 0 1732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1711307567
transform 1 0 1596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1711307567
transform 1 0 1548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1711307567
transform 1 0 1012 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1711307567
transform 1 0 1012 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1711307567
transform 1 0 996 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1711307567
transform 1 0 996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1711307567
transform 1 0 900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1711307567
transform 1 0 876 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1711307567
transform 1 0 444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1711307567
transform 1 0 300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1711307567
transform 1 0 2444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1711307567
transform 1 0 2236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1711307567
transform 1 0 1988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1711307567
transform 1 0 388 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1711307567
transform 1 0 364 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1711307567
transform 1 0 1996 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1711307567
transform 1 0 1972 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1711307567
transform 1 0 1644 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1711307567
transform 1 0 1588 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1711307567
transform 1 0 1524 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1711307567
transform 1 0 1428 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1711307567
transform 1 0 1324 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1711307567
transform 1 0 1300 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1711307567
transform 1 0 1172 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1711307567
transform 1 0 1172 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1711307567
transform 1 0 1036 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1711307567
transform 1 0 924 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1711307567
transform 1 0 780 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1711307567
transform 1 0 684 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1711307567
transform 1 0 572 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1711307567
transform 1 0 484 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1711307567
transform 1 0 380 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1711307567
transform 1 0 364 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1711307567
transform 1 0 316 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1711307567
transform 1 0 316 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1711307567
transform 1 0 284 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1711307567
transform 1 0 2292 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1711307567
transform 1 0 2284 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1711307567
transform 1 0 2220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1711307567
transform 1 0 1596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1711307567
transform 1 0 1436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1711307567
transform 1 0 1276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1711307567
transform 1 0 1228 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1711307567
transform 1 0 1116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1711307567
transform 1 0 956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1711307567
transform 1 0 948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1711307567
transform 1 0 836 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1711307567
transform 1 0 708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1711307567
transform 1 0 644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1711307567
transform 1 0 580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1711307567
transform 1 0 2564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1711307567
transform 1 0 2444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1711307567
transform 1 0 2276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1711307567
transform 1 0 2212 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1711307567
transform 1 0 2092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1711307567
transform 1 0 1716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1711307567
transform 1 0 1452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1711307567
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1711307567
transform 1 0 412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1711307567
transform 1 0 308 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1711307567
transform 1 0 228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1711307567
transform 1 0 212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1711307567
transform 1 0 212 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1711307567
transform 1 0 212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1711307567
transform 1 0 196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1711307567
transform 1 0 2620 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1711307567
transform 1 0 2564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1711307567
transform 1 0 2564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1711307567
transform 1 0 2548 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1711307567
transform 1 0 2500 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1711307567
transform 1 0 2308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1711307567
transform 1 0 2212 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1711307567
transform 1 0 1996 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1711307567
transform 1 0 1988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1711307567
transform 1 0 1948 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1711307567
transform 1 0 1924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1711307567
transform 1 0 1892 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1711307567
transform 1 0 2124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1711307567
transform 1 0 2076 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1711307567
transform 1 0 2068 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1711307567
transform 1 0 2060 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1711307567
transform 1 0 1980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1711307567
transform 1 0 1908 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1711307567
transform 1 0 1836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1711307567
transform 1 0 1820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1711307567
transform 1 0 1300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1711307567
transform 1 0 1228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1711307567
transform 1 0 1012 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1711307567
transform 1 0 964 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1711307567
transform 1 0 748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1711307567
transform 1 0 732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1711307567
transform 1 0 676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1711307567
transform 1 0 676 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1711307567
transform 1 0 2284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1711307567
transform 1 0 2148 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1711307567
transform 1 0 1900 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1711307567
transform 1 0 1572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1711307567
transform 1 0 1452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1711307567
transform 1 0 452 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1711307567
transform 1 0 388 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1711307567
transform 1 0 1724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1711307567
transform 1 0 1708 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1711307567
transform 1 0 1476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1711307567
transform 1 0 1476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1711307567
transform 1 0 1020 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1711307567
transform 1 0 1004 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1711307567
transform 1 0 988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1711307567
transform 1 0 964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1711307567
transform 1 0 532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1711307567
transform 1 0 532 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1711307567
transform 1 0 1572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1711307567
transform 1 0 1540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1711307567
transform 1 0 1028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1711307567
transform 1 0 996 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1711307567
transform 1 0 2668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1711307567
transform 1 0 2652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1711307567
transform 1 0 1868 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1711307567
transform 1 0 1612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1711307567
transform 1 0 1780 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1711307567
transform 1 0 356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1711307567
transform 1 0 2188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1711307567
transform 1 0 2140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1711307567
transform 1 0 2116 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1711307567
transform 1 0 1780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1711307567
transform 1 0 1708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1711307567
transform 1 0 1676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1711307567
transform 1 0 876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1711307567
transform 1 0 724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1711307567
transform 1 0 540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1711307567
transform 1 0 2188 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1711307567
transform 1 0 2156 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1711307567
transform 1 0 796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1711307567
transform 1 0 748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1711307567
transform 1 0 628 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1711307567
transform 1 0 540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1711307567
transform 1 0 548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1711307567
transform 1 0 364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1711307567
transform 1 0 340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1711307567
transform 1 0 300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1711307567
transform 1 0 692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1711307567
transform 1 0 684 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1711307567
transform 1 0 452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1711307567
transform 1 0 452 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1711307567
transform 1 0 1572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1711307567
transform 1 0 1444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1711307567
transform 1 0 780 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1711307567
transform 1 0 588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1711307567
transform 1 0 1500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1711307567
transform 1 0 1428 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1711307567
transform 1 0 804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1711307567
transform 1 0 580 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1711307567
transform 1 0 1900 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1711307567
transform 1 0 1796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1711307567
transform 1 0 1156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1711307567
transform 1 0 716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1711307567
transform 1 0 388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1711307567
transform 1 0 772 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1711307567
transform 1 0 716 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1711307567
transform 1 0 676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1711307567
transform 1 0 604 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1711307567
transform 1 0 596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1711307567
transform 1 0 596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1711307567
transform 1 0 1508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1711307567
transform 1 0 1284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1711307567
transform 1 0 1284 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1711307567
transform 1 0 1252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1711307567
transform 1 0 1244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1711307567
transform 1 0 1140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1711307567
transform 1 0 1428 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1711307567
transform 1 0 1364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1711307567
transform 1 0 1308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1711307567
transform 1 0 1292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1711307567
transform 1 0 1220 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1711307567
transform 1 0 2324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1711307567
transform 1 0 1612 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1711307567
transform 1 0 1548 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1711307567
transform 1 0 1548 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1711307567
transform 1 0 1508 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1711307567
transform 1 0 1436 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1711307567
transform 1 0 1348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1711307567
transform 1 0 1164 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1711307567
transform 1 0 1156 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1711307567
transform 1 0 884 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1711307567
transform 1 0 828 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1711307567
transform 1 0 756 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1711307567
transform 1 0 484 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1711307567
transform 1 0 428 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1711307567
transform 1 0 380 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1711307567
transform 1 0 340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1711307567
transform 1 0 340 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1711307567
transform 1 0 324 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1711307567
transform 1 0 300 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1711307567
transform 1 0 284 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1711307567
transform 1 0 284 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1711307567
transform 1 0 1356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1711307567
transform 1 0 1076 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1711307567
transform 1 0 2220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1711307567
transform 1 0 2180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1711307567
transform 1 0 2108 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1711307567
transform 1 0 508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1711307567
transform 1 0 420 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1711307567
transform 1 0 356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1711307567
transform 1 0 2276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1711307567
transform 1 0 2220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1711307567
transform 1 0 2204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1711307567
transform 1 0 2204 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1711307567
transform 1 0 2164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1711307567
transform 1 0 1980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1711307567
transform 1 0 1756 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1711307567
transform 1 0 1380 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1711307567
transform 1 0 764 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1711307567
transform 1 0 548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1711307567
transform 1 0 1948 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1711307567
transform 1 0 1852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1711307567
transform 1 0 1228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1711307567
transform 1 0 732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1711307567
transform 1 0 420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1711307567
transform 1 0 2284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1711307567
transform 1 0 2260 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1711307567
transform 1 0 2036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1711307567
transform 1 0 2036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1711307567
transform 1 0 1684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1711307567
transform 1 0 1564 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1711307567
transform 1 0 1556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1711307567
transform 1 0 1460 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1711307567
transform 1 0 1380 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1711307567
transform 1 0 948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1711307567
transform 1 0 948 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1711307567
transform 1 0 540 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1711307567
transform 1 0 492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1711307567
transform 1 0 348 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1711307567
transform 1 0 2732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1711307567
transform 1 0 2724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1711307567
transform 1 0 2724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1711307567
transform 1 0 2700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1711307567
transform 1 0 2684 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1711307567
transform 1 0 2684 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1711307567
transform 1 0 2556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1711307567
transform 1 0 2044 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1711307567
transform 1 0 2020 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1711307567
transform 1 0 1996 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1711307567
transform 1 0 1180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1711307567
transform 1 0 1172 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1711307567
transform 1 0 1164 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1711307567
transform 1 0 1148 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1711307567
transform 1 0 884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1711307567
transform 1 0 788 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1711307567
transform 1 0 764 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1711307567
transform 1 0 700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1711307567
transform 1 0 692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1711307567
transform 1 0 620 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1711307567
transform 1 0 540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1711307567
transform 1 0 244 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1711307567
transform 1 0 244 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1711307567
transform 1 0 2740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1711307567
transform 1 0 2652 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1711307567
transform 1 0 2580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1711307567
transform 1 0 2564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1711307567
transform 1 0 2732 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1711307567
transform 1 0 2668 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1711307567
transform 1 0 2748 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1711307567
transform 1 0 2740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1711307567
transform 1 0 2740 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1711307567
transform 1 0 2708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1711307567
transform 1 0 2636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1711307567
transform 1 0 2612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1711307567
transform 1 0 2588 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1711307567
transform 1 0 2532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1711307567
transform 1 0 2596 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1711307567
transform 1 0 2292 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1711307567
transform 1 0 2588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1711307567
transform 1 0 2508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1711307567
transform 1 0 2524 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1711307567
transform 1 0 2412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1711307567
transform 1 0 2524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1711307567
transform 1 0 2452 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1711307567
transform 1 0 2532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1711307567
transform 1 0 2532 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1711307567
transform 1 0 2716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1711307567
transform 1 0 2708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1711307567
transform 1 0 2564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1711307567
transform 1 0 2468 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1711307567
transform 1 0 2020 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1711307567
transform 1 0 2012 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1711307567
transform 1 0 1996 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1711307567
transform 1 0 1892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1711307567
transform 1 0 1876 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1711307567
transform 1 0 1860 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1711307567
transform 1 0 2500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1711307567
transform 1 0 2500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1711307567
transform 1 0 2348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1711307567
transform 1 0 2308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1711307567
transform 1 0 2412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1711307567
transform 1 0 2412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1711307567
transform 1 0 2316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1711307567
transform 1 0 2276 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1711307567
transform 1 0 2228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1711307567
transform 1 0 2204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1711307567
transform 1 0 2444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1711307567
transform 1 0 2404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1711307567
transform 1 0 2628 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1711307567
transform 1 0 2588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1711307567
transform 1 0 2220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1711307567
transform 1 0 1964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1711307567
transform 1 0 2468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1711307567
transform 1 0 2236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1711307567
transform 1 0 2372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1711307567
transform 1 0 2204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1711307567
transform 1 0 1868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1711307567
transform 1 0 1868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1711307567
transform 1 0 1660 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1711307567
transform 1 0 1660 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1711307567
transform 1 0 1740 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1711307567
transform 1 0 1740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1711307567
transform 1 0 1748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1711307567
transform 1 0 1540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1711307567
transform 1 0 1548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1711307567
transform 1 0 1540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1711307567
transform 1 0 1636 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1711307567
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1711307567
transform 1 0 1340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1711307567
transform 1 0 1340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1711307567
transform 1 0 1204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1711307567
transform 1 0 1204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1711307567
transform 1 0 1388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1711307567
transform 1 0 1388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1711307567
transform 1 0 1260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1711307567
transform 1 0 1260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1711307567
transform 1 0 1084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1711307567
transform 1 0 924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1711307567
transform 1 0 1092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1711307567
transform 1 0 1044 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1711307567
transform 1 0 876 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1711307567
transform 1 0 852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1711307567
transform 1 0 972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1711307567
transform 1 0 972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1711307567
transform 1 0 628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1711307567
transform 1 0 628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1711307567
transform 1 0 708 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1711307567
transform 1 0 708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1711307567
transform 1 0 796 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1711307567
transform 1 0 796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1711307567
transform 1 0 516 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1711307567
transform 1 0 484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1711307567
transform 1 0 404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1711307567
transform 1 0 396 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1711307567
transform 1 0 436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1711307567
transform 1 0 180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1711307567
transform 1 0 396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1711307567
transform 1 0 356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1711307567
transform 1 0 316 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1711307567
transform 1 0 268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1711307567
transform 1 0 1452 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1711307567
transform 1 0 1444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1711307567
transform 1 0 1428 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1711307567
transform 1 0 1428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1711307567
transform 1 0 1428 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1711307567
transform 1 0 1420 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1711307567
transform 1 0 1476 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1711307567
transform 1 0 1476 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1711307567
transform 1 0 1420 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1711307567
transform 1 0 1380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1711307567
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1711307567
transform 1 0 1452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1711307567
transform 1 0 1468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1711307567
transform 1 0 1460 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1711307567
transform 1 0 1436 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1711307567
transform 1 0 1428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1711307567
transform 1 0 1628 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1711307567
transform 1 0 1452 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1711307567
transform 1 0 1468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1711307567
transform 1 0 1068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1711307567
transform 1 0 1028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1711307567
transform 1 0 572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1711307567
transform 1 0 572 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1711307567
transform 1 0 1228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1711307567
transform 1 0 1124 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1711307567
transform 1 0 1724 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1711307567
transform 1 0 1668 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1711307567
transform 1 0 1604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1711307567
transform 1 0 1628 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1711307567
transform 1 0 692 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1711307567
transform 1 0 612 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1711307567
transform 1 0 516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1711307567
transform 1 0 572 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1711307567
transform 1 0 492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1711307567
transform 1 0 292 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1711307567
transform 1 0 588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1711307567
transform 1 0 564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1711307567
transform 1 0 540 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1711307567
transform 1 0 340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1711307567
transform 1 0 292 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1711307567
transform 1 0 572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1711307567
transform 1 0 532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1711307567
transform 1 0 476 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1711307567
transform 1 0 500 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1711307567
transform 1 0 484 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1711307567
transform 1 0 1508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1711307567
transform 1 0 1084 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1711307567
transform 1 0 468 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1711307567
transform 1 0 476 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1711307567
transform 1 0 436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1711307567
transform 1 0 396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1711307567
transform 1 0 1476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1711307567
transform 1 0 1140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1711307567
transform 1 0 548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1711307567
transform 1 0 492 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1711307567
transform 1 0 484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1711307567
transform 1 0 452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1711307567
transform 1 0 436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1711307567
transform 1 0 428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1711307567
transform 1 0 404 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1711307567
transform 1 0 356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1711307567
transform 1 0 340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1711307567
transform 1 0 260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1711307567
transform 1 0 244 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1711307567
transform 1 0 412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1711307567
transform 1 0 316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1711307567
transform 1 0 260 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1711307567
transform 1 0 1804 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1711307567
transform 1 0 1708 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1711307567
transform 1 0 1772 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1711307567
transform 1 0 1740 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1711307567
transform 1 0 2204 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1711307567
transform 1 0 2164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1711307567
transform 1 0 1740 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1711307567
transform 1 0 1636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1711307567
transform 1 0 1524 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1711307567
transform 1 0 1492 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1711307567
transform 1 0 1476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1711307567
transform 1 0 1756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1711307567
transform 1 0 1756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1711307567
transform 1 0 1740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1711307567
transform 1 0 2132 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1711307567
transform 1 0 1772 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1711307567
transform 1 0 1652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1711307567
transform 1 0 1844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1711307567
transform 1 0 1796 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1711307567
transform 1 0 1780 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1711307567
transform 1 0 1940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1711307567
transform 1 0 1860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1711307567
transform 1 0 2084 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1711307567
transform 1 0 1948 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1711307567
transform 1 0 1924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1711307567
transform 1 0 2132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1711307567
transform 1 0 1964 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1711307567
transform 1 0 1964 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1711307567
transform 1 0 1308 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1711307567
transform 1 0 1028 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1711307567
transform 1 0 1412 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1711307567
transform 1 0 1332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1711307567
transform 1 0 1356 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1711307567
transform 1 0 1324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1711307567
transform 1 0 1484 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1711307567
transform 1 0 1388 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1711307567
transform 1 0 1700 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1711307567
transform 1 0 1692 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1711307567
transform 1 0 1676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1711307567
transform 1 0 1644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1711307567
transform 1 0 1644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1711307567
transform 1 0 1628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1711307567
transform 1 0 1628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1711307567
transform 1 0 1628 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1711307567
transform 1 0 1580 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1711307567
transform 1 0 1420 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1711307567
transform 1 0 1372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1711307567
transform 1 0 1484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1711307567
transform 1 0 1484 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1711307567
transform 1 0 1436 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1711307567
transform 1 0 1444 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1711307567
transform 1 0 1420 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1711307567
transform 1 0 1404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1711307567
transform 1 0 1284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1711307567
transform 1 0 1284 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1711307567
transform 1 0 1668 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1711307567
transform 1 0 1556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1711307567
transform 1 0 1436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1711307567
transform 1 0 1244 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1711307567
transform 1 0 1220 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1711307567
transform 1 0 1348 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1711307567
transform 1 0 1284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1711307567
transform 1 0 1396 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1711307567
transform 1 0 1396 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1711307567
transform 1 0 1580 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1711307567
transform 1 0 1484 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1711307567
transform 1 0 1484 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1711307567
transform 1 0 1324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1711307567
transform 1 0 1308 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1711307567
transform 1 0 1252 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1711307567
transform 1 0 1204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1711307567
transform 1 0 1260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1711307567
transform 1 0 1148 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1711307567
transform 1 0 988 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1711307567
transform 1 0 956 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1711307567
transform 1 0 1412 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1711307567
transform 1 0 1372 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1711307567
transform 1 0 1364 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1711307567
transform 1 0 1196 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1711307567
transform 1 0 996 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1711307567
transform 1 0 980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1711307567
transform 1 0 972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1711307567
transform 1 0 852 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1711307567
transform 1 0 844 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1711307567
transform 1 0 836 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1711307567
transform 1 0 820 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1711307567
transform 1 0 796 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1711307567
transform 1 0 772 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1711307567
transform 1 0 764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1711307567
transform 1 0 756 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1711307567
transform 1 0 996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1711307567
transform 1 0 980 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1711307567
transform 1 0 812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1711307567
transform 1 0 932 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1711307567
transform 1 0 724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1711307567
transform 1 0 1052 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1711307567
transform 1 0 972 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1711307567
transform 1 0 1068 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1711307567
transform 1 0 1028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1711307567
transform 1 0 1004 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1711307567
transform 1 0 1068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1711307567
transform 1 0 1052 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1711307567
transform 1 0 1036 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1711307567
transform 1 0 724 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1711307567
transform 1 0 668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1711307567
transform 1 0 644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1711307567
transform 1 0 740 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1711307567
transform 1 0 740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1711307567
transform 1 0 716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1711307567
transform 1 0 700 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1711307567
transform 1 0 1260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1711307567
transform 1 0 1156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1711307567
transform 1 0 1140 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1711307567
transform 1 0 1356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1711307567
transform 1 0 860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1711307567
transform 1 0 1396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1711307567
transform 1 0 1316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1711307567
transform 1 0 1412 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1711307567
transform 1 0 1412 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1711307567
transform 1 0 1428 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1711307567
transform 1 0 1404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1711307567
transform 1 0 1356 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1711307567
transform 1 0 1268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1711307567
transform 1 0 1388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1711307567
transform 1 0 1388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1711307567
transform 1 0 1364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1711307567
transform 1 0 1364 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1711307567
transform 1 0 1188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1711307567
transform 1 0 1132 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1711307567
transform 1 0 1676 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1711307567
transform 1 0 1668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1711307567
transform 1 0 1596 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1711307567
transform 1 0 1532 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1711307567
transform 1 0 1348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1711307567
transform 1 0 1340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1711307567
transform 1 0 1332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1711307567
transform 1 0 1404 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1711307567
transform 1 0 1404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1711307567
transform 1 0 1596 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1711307567
transform 1 0 1588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1711307567
transform 1 0 1548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1711307567
transform 1 0 1396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1711307567
transform 1 0 1500 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1711307567
transform 1 0 1492 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1711307567
transform 1 0 1476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1711307567
transform 1 0 1468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1711307567
transform 1 0 1452 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1711307567
transform 1 0 1236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1711307567
transform 1 0 1188 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1711307567
transform 1 0 1172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1711307567
transform 1 0 636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1711307567
transform 1 0 572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1711307567
transform 1 0 1212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1711307567
transform 1 0 1212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1711307567
transform 1 0 1164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1711307567
transform 1 0 1052 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1711307567
transform 1 0 1052 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1711307567
transform 1 0 1292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1711307567
transform 1 0 1268 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1711307567
transform 1 0 1676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1711307567
transform 1 0 1604 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1711307567
transform 1 0 1444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1711307567
transform 1 0 1284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1711307567
transform 1 0 1308 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1711307567
transform 1 0 1156 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1711307567
transform 1 0 940 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1711307567
transform 1 0 940 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1711307567
transform 1 0 1452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1711307567
transform 1 0 1420 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1711307567
transform 1 0 1540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1711307567
transform 1 0 1452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1711307567
transform 1 0 2004 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1711307567
transform 1 0 1796 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1711307567
transform 1 0 1732 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1711307567
transform 1 0 1516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1711307567
transform 1 0 1540 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1711307567
transform 1 0 572 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1711307567
transform 1 0 1132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1711307567
transform 1 0 1092 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1711307567
transform 1 0 828 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1711307567
transform 1 0 620 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1711307567
transform 1 0 604 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1711307567
transform 1 0 580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1711307567
transform 1 0 556 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1711307567
transform 1 0 556 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1711307567
transform 1 0 564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1711307567
transform 1 0 532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1711307567
transform 1 0 460 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1711307567
transform 1 0 428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1711307567
transform 1 0 1396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1711307567
transform 1 0 1276 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1711307567
transform 1 0 1268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1711307567
transform 1 0 1204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1711307567
transform 1 0 1436 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1711307567
transform 1 0 1412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1711307567
transform 1 0 1516 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1711307567
transform 1 0 1372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1711307567
transform 1 0 1300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1711307567
transform 1 0 1300 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1711307567
transform 1 0 1300 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1711307567
transform 1 0 1044 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1711307567
transform 1 0 1012 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1711307567
transform 1 0 1996 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1711307567
transform 1 0 1988 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1711307567
transform 1 0 1908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1711307567
transform 1 0 1668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1711307567
transform 1 0 1428 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1711307567
transform 1 0 1388 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1711307567
transform 1 0 1700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1711307567
transform 1 0 1660 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1711307567
transform 1 0 1644 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1711307567
transform 1 0 1420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1711307567
transform 1 0 804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1711307567
transform 1 0 708 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1711307567
transform 1 0 932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1711307567
transform 1 0 868 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1711307567
transform 1 0 980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1711307567
transform 1 0 948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1711307567
transform 1 0 940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1711307567
transform 1 0 796 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1711307567
transform 1 0 636 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1711307567
transform 1 0 636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1711307567
transform 1 0 972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1711307567
transform 1 0 964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1711307567
transform 1 0 956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1711307567
transform 1 0 1044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1711307567
transform 1 0 1020 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1711307567
transform 1 0 1436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1711307567
transform 1 0 1316 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1711307567
transform 1 0 1268 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1711307567
transform 1 0 1044 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1711307567
transform 1 0 1020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1711307567
transform 1 0 1036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1711307567
transform 1 0 948 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1711307567
transform 1 0 940 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1711307567
transform 1 0 932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1711307567
transform 1 0 1604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1711307567
transform 1 0 868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1711307567
transform 1 0 892 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1711307567
transform 1 0 844 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1711307567
transform 1 0 788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1711307567
transform 1 0 372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1711307567
transform 1 0 1988 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1711307567
transform 1 0 1940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1711307567
transform 1 0 1820 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1711307567
transform 1 0 1732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1711307567
transform 1 0 1652 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1711307567
transform 1 0 396 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1711307567
transform 1 0 340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1711307567
transform 1 0 364 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1711307567
transform 1 0 356 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1711307567
transform 1 0 1828 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1711307567
transform 1 0 1596 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1711307567
transform 1 0 1612 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1711307567
transform 1 0 1556 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1711307567
transform 1 0 1524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1711307567
transform 1 0 1820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1711307567
transform 1 0 1804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1711307567
transform 1 0 1804 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1711307567
transform 1 0 2028 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1711307567
transform 1 0 1812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1711307567
transform 1 0 1804 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1711307567
transform 1 0 1708 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1711307567
transform 1 0 1692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1711307567
transform 1 0 1556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1711307567
transform 1 0 1876 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1711307567
transform 1 0 1852 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1711307567
transform 1 0 668 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1711307567
transform 1 0 668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1711307567
transform 1 0 748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1711307567
transform 1 0 700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1711307567
transform 1 0 724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1711307567
transform 1 0 604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1711307567
transform 1 0 468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1711307567
transform 1 0 452 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1711307567
transform 1 0 764 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1711307567
transform 1 0 732 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1711307567
transform 1 0 732 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1711307567
transform 1 0 692 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1711307567
transform 1 0 1268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1711307567
transform 1 0 772 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1711307567
transform 1 0 556 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1711307567
transform 1 0 412 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1711307567
transform 1 0 260 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1711307567
transform 1 0 228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1711307567
transform 1 0 180 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1711307567
transform 1 0 804 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1711307567
transform 1 0 596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1711307567
transform 1 0 484 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1711307567
transform 1 0 852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1711307567
transform 1 0 652 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1711307567
transform 1 0 1380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1711307567
transform 1 0 1372 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1711307567
transform 1 0 1292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1711307567
transform 1 0 1052 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1711307567
transform 1 0 1036 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1711307567
transform 1 0 1316 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1711307567
transform 1 0 1316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1711307567
transform 1 0 1284 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1711307567
transform 1 0 876 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1711307567
transform 1 0 940 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1711307567
transform 1 0 844 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1711307567
transform 1 0 860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1711307567
transform 1 0 708 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1711307567
transform 1 0 628 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1711307567
transform 1 0 580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1711307567
transform 1 0 716 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1711307567
transform 1 0 700 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1711307567
transform 1 0 676 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1711307567
transform 1 0 500 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1711307567
transform 1 0 332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1711307567
transform 1 0 1220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1711307567
transform 1 0 716 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1711307567
transform 1 0 508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1711307567
transform 1 0 364 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1711307567
transform 1 0 340 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1711307567
transform 1 0 300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1711307567
transform 1 0 884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1711307567
transform 1 0 580 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1711307567
transform 1 0 1660 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1711307567
transform 1 0 1644 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1711307567
transform 1 0 1436 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1711307567
transform 1 0 844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1711307567
transform 1 0 1004 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1711307567
transform 1 0 908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1711307567
transform 1 0 868 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1711307567
transform 1 0 964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1711307567
transform 1 0 964 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1711307567
transform 1 0 900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1711307567
transform 1 0 892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1711307567
transform 1 0 892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1711307567
transform 1 0 708 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1711307567
transform 1 0 660 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1711307567
transform 1 0 1564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1711307567
transform 1 0 900 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1711307567
transform 1 0 908 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1711307567
transform 1 0 844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1711307567
transform 1 0 916 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1711307567
transform 1 0 916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1711307567
transform 1 0 1220 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1711307567
transform 1 0 948 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1711307567
transform 1 0 1236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1711307567
transform 1 0 1204 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1711307567
transform 1 0 1332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1711307567
transform 1 0 1212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1711307567
transform 1 0 1244 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1711307567
transform 1 0 956 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1711307567
transform 1 0 900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1711307567
transform 1 0 772 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1711307567
transform 1 0 652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1711307567
transform 1 0 604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1711307567
transform 1 0 748 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1711307567
transform 1 0 460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1711307567
transform 1 0 412 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1711307567
transform 1 0 396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1711307567
transform 1 0 412 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1711307567
transform 1 0 300 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1711307567
transform 1 0 292 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1711307567
transform 1 0 276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1711307567
transform 1 0 332 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1711307567
transform 1 0 324 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1711307567
transform 1 0 324 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1711307567
transform 1 0 324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1711307567
transform 1 0 1828 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1711307567
transform 1 0 1556 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1711307567
transform 1 0 1572 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1711307567
transform 1 0 1532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1711307567
transform 1 0 1532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1711307567
transform 1 0 1804 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1711307567
transform 1 0 1804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1711307567
transform 1 0 1924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1711307567
transform 1 0 1868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1711307567
transform 1 0 2052 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1711307567
transform 1 0 1884 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1711307567
transform 1 0 1836 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1711307567
transform 1 0 1836 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1711307567
transform 1 0 1772 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1711307567
transform 1 0 1996 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1711307567
transform 1 0 1916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1711307567
transform 1 0 2068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1711307567
transform 1 0 1948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1711307567
transform 1 0 1932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1711307567
transform 1 0 1260 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1711307567
transform 1 0 1260 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1711307567
transform 1 0 1348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1711307567
transform 1 0 1276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1711307567
transform 1 0 1276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1711307567
transform 1 0 1244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1711307567
transform 1 0 1468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1711307567
transform 1 0 1348 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1711307567
transform 1 0 1228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1711307567
transform 1 0 692 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1711307567
transform 1 0 460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1711307567
transform 1 0 436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1711307567
transform 1 0 1340 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1711307567
transform 1 0 1316 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1711307567
transform 1 0 1324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1711307567
transform 1 0 1316 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1711307567
transform 1 0 1508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1711307567
transform 1 0 1372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1711307567
transform 1 0 1788 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1711307567
transform 1 0 1628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1711307567
transform 1 0 1468 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1711307567
transform 1 0 1492 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1711307567
transform 1 0 588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1711307567
transform 1 0 580 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1711307567
transform 1 0 572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1711307567
transform 1 0 444 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1711307567
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1711307567
transform 1 0 1276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1711307567
transform 1 0 1172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1711307567
transform 1 0 1172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1711307567
transform 1 0 1340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1711307567
transform 1 0 1324 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1711307567
transform 1 0 1676 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1711307567
transform 1 0 1660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1711307567
transform 1 0 1572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1711307567
transform 1 0 1380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1711307567
transform 1 0 788 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1711307567
transform 1 0 708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1711307567
transform 1 0 652 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1711307567
transform 1 0 1564 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1711307567
transform 1 0 1548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1711307567
transform 1 0 1452 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1711307567
transform 1 0 1308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1711307567
transform 1 0 2092 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1711307567
transform 1 0 2068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1711307567
transform 1 0 2036 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1711307567
transform 1 0 1708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1711307567
transform 1 0 1876 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1711307567
transform 1 0 1756 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1711307567
transform 1 0 1652 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1711307567
transform 1 0 1948 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1711307567
transform 1 0 1780 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1711307567
transform 1 0 1588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1711307567
transform 1 0 1524 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1711307567
transform 1 0 1444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1711307567
transform 1 0 1708 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1711307567
transform 1 0 1636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1711307567
transform 1 0 1636 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1711307567
transform 1 0 2052 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1711307567
transform 1 0 1732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1711307567
transform 1 0 1708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1711307567
transform 1 0 212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1711307567
transform 1 0 140 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1711307567
transform 1 0 276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1711307567
transform 1 0 180 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1711307567
transform 1 0 268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1711307567
transform 1 0 188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1711307567
transform 1 0 316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1711307567
transform 1 0 292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1711307567
transform 1 0 532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1711307567
transform 1 0 308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1711307567
transform 1 0 268 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1711307567
transform 1 0 300 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1711307567
transform 1 0 212 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1711307567
transform 1 0 1948 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1711307567
transform 1 0 212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1711307567
transform 1 0 188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1711307567
transform 1 0 188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1711307567
transform 1 0 132 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1711307567
transform 1 0 244 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1711307567
transform 1 0 164 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1711307567
transform 1 0 236 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1711307567
transform 1 0 172 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1711307567
transform 1 0 284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1711307567
transform 1 0 252 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1711307567
transform 1 0 324 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1711307567
transform 1 0 300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1711307567
transform 1 0 252 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1711307567
transform 1 0 252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1711307567
transform 1 0 220 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1711307567
transform 1 0 548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1711307567
transform 1 0 276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1711307567
transform 1 0 276 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1711307567
transform 1 0 172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1711307567
transform 1 0 124 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1711307567
transform 1 0 180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1711307567
transform 1 0 148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1711307567
transform 1 0 212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1711307567
transform 1 0 156 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1711307567
transform 1 0 308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1711307567
transform 1 0 228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1711307567
transform 1 0 188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1711307567
transform 1 0 188 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1711307567
transform 1 0 276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1711307567
transform 1 0 236 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1711307567
transform 1 0 268 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1711307567
transform 1 0 260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1711307567
transform 1 0 1108 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1711307567
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1711307567
transform 1 0 308 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1711307567
transform 1 0 276 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1711307567
transform 1 0 548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1711307567
transform 1 0 388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1711307567
transform 1 0 268 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1711307567
transform 1 0 236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1711307567
transform 1 0 324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1711307567
transform 1 0 324 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1711307567
transform 1 0 2420 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1711307567
transform 1 0 1788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1711307567
transform 1 0 1756 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1711307567
transform 1 0 1956 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1711307567
transform 1 0 1956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1711307567
transform 1 0 1740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1711307567
transform 1 0 660 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1711307567
transform 1 0 660 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1711307567
transform 1 0 636 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1711307567
transform 1 0 636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1711307567
transform 1 0 620 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1711307567
transform 1 0 620 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1711307567
transform 1 0 604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1711307567
transform 1 0 380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1711307567
transform 1 0 300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1711307567
transform 1 0 332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1711307567
transform 1 0 308 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1711307567
transform 1 0 268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1711307567
transform 1 0 252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1711307567
transform 1 0 2348 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1711307567
transform 1 0 1996 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1711307567
transform 1 0 1620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1711307567
transform 1 0 972 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1711307567
transform 1 0 668 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1711307567
transform 1 0 476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1711307567
transform 1 0 452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1711307567
transform 1 0 436 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1711307567
transform 1 0 420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1711307567
transform 1 0 348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1711307567
transform 1 0 348 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1711307567
transform 1 0 380 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1711307567
transform 1 0 372 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1711307567
transform 1 0 300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1711307567
transform 1 0 300 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1711307567
transform 1 0 500 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1711307567
transform 1 0 356 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1711307567
transform 1 0 2372 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1711307567
transform 1 0 1940 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1711307567
transform 1 0 1940 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1711307567
transform 1 0 660 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1711307567
transform 1 0 524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1711307567
transform 1 0 1988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1711307567
transform 1 0 1900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1711307567
transform 1 0 1540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1711307567
transform 1 0 1052 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1711307567
transform 1 0 644 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1711307567
transform 1 0 484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1711307567
transform 1 0 396 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1711307567
transform 1 0 428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1711307567
transform 1 0 412 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1711307567
transform 1 0 540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1711307567
transform 1 0 476 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1711307567
transform 1 0 476 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1711307567
transform 1 0 444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1711307567
transform 1 0 444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1711307567
transform 1 0 492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1711307567
transform 1 0 468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1711307567
transform 1 0 2084 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1711307567
transform 1 0 1988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1711307567
transform 1 0 1572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1711307567
transform 1 0 1124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1711307567
transform 1 0 668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1711307567
transform 1 0 748 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1711307567
transform 1 0 748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1711307567
transform 1 0 700 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1711307567
transform 1 0 604 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1711307567
transform 1 0 396 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1711307567
transform 1 0 372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1711307567
transform 1 0 348 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1711307567
transform 1 0 324 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1711307567
transform 1 0 884 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1711307567
transform 1 0 572 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1711307567
transform 1 0 556 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1711307567
transform 1 0 516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1711307567
transform 1 0 484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1711307567
transform 1 0 404 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1711307567
transform 1 0 2132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1711307567
transform 1 0 2060 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1711307567
transform 1 0 1612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1711307567
transform 1 0 1124 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1711307567
transform 1 0 644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1711307567
transform 1 0 612 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1711307567
transform 1 0 532 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1711307567
transform 1 0 444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1711307567
transform 1 0 476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1711307567
transform 1 0 452 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1711307567
transform 1 0 452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1711307567
transform 1 0 452 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1711307567
transform 1 0 580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1711307567
transform 1 0 500 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1711307567
transform 1 0 764 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1711307567
transform 1 0 692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1711307567
transform 1 0 508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1711307567
transform 1 0 460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1711307567
transform 1 0 420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1711307567
transform 1 0 788 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1711307567
transform 1 0 788 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1711307567
transform 1 0 820 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1711307567
transform 1 0 820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1711307567
transform 1 0 796 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1711307567
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1711307567
transform 1 0 732 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1711307567
transform 1 0 1852 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1711307567
transform 1 0 1676 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1711307567
transform 1 0 1580 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1711307567
transform 1 0 1484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1711307567
transform 1 0 1156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1711307567
transform 1 0 1140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1711307567
transform 1 0 764 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1711307567
transform 1 0 756 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1711307567
transform 1 0 788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1711307567
transform 1 0 748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1711307567
transform 1 0 716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1711307567
transform 1 0 612 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1711307567
transform 1 0 812 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1711307567
transform 1 0 732 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1711307567
transform 1 0 684 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1711307567
transform 1 0 684 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1711307567
transform 1 0 724 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1711307567
transform 1 0 716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1711307567
transform 1 0 772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1711307567
transform 1 0 772 0 1 1845
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1711307567
transform 1 0 764 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1711307567
transform 1 0 868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1711307567
transform 1 0 732 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1711307567
transform 1 0 644 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1711307567
transform 1 0 684 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1711307567
transform 1 0 676 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1711307567
transform 1 0 700 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1711307567
transform 1 0 668 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1711307567
transform 1 0 732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1711307567
transform 1 0 724 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1711307567
transform 1 0 724 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1711307567
transform 1 0 788 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1711307567
transform 1 0 748 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1711307567
transform 1 0 644 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1711307567
transform 1 0 620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1711307567
transform 1 0 620 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1711307567
transform 1 0 620 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1711307567
transform 1 0 900 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1711307567
transform 1 0 796 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1711307567
transform 1 0 612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1711307567
transform 1 0 708 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1711307567
transform 1 0 612 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1711307567
transform 1 0 580 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1711307567
transform 1 0 564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1711307567
transform 1 0 556 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1711307567
transform 1 0 628 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1711307567
transform 1 0 596 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1711307567
transform 1 0 996 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1711307567
transform 1 0 964 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1711307567
transform 1 0 988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1711307567
transform 1 0 972 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1711307567
transform 1 0 1012 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1711307567
transform 1 0 932 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1711307567
transform 1 0 876 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1711307567
transform 1 0 916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1711307567
transform 1 0 916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1711307567
transform 1 0 964 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1711307567
transform 1 0 964 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1711307567
transform 1 0 860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1711307567
transform 1 0 820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1711307567
transform 1 0 820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1711307567
transform 1 0 812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1711307567
transform 1 0 852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1711307567
transform 1 0 844 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1711307567
transform 1 0 1076 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1711307567
transform 1 0 1052 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1711307567
transform 1 0 892 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1711307567
transform 1 0 1996 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1711307567
transform 1 0 1116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1711307567
transform 1 0 1116 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1711307567
transform 1 0 1052 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1711307567
transform 1 0 972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1711307567
transform 1 0 956 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1711307567
transform 1 0 1076 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1711307567
transform 1 0 1028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1711307567
transform 1 0 1020 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1711307567
transform 1 0 1020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1711307567
transform 1 0 1116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1711307567
transform 1 0 1028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1711307567
transform 1 0 988 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1711307567
transform 1 0 980 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1711307567
transform 1 0 1156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1711307567
transform 1 0 1092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1711307567
transform 1 0 924 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1711307567
transform 1 0 900 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1711307567
transform 1 0 972 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1711307567
transform 1 0 956 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1711307567
transform 1 0 1052 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1711307567
transform 1 0 980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1711307567
transform 1 0 1140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1711307567
transform 1 0 1100 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1711307567
transform 1 0 1068 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1711307567
transform 1 0 1052 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1711307567
transform 1 0 1180 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1711307567
transform 1 0 1108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1711307567
transform 1 0 1108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1711307567
transform 1 0 1228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1711307567
transform 1 0 1204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1711307567
transform 1 0 1196 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1711307567
transform 1 0 1156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1711307567
transform 1 0 1244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1711307567
transform 1 0 1236 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1711307567
transform 1 0 1236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1711307567
transform 1 0 1164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1711307567
transform 1 0 1068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1711307567
transform 1 0 1148 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1711307567
transform 1 0 1012 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1711307567
transform 1 0 1492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1711307567
transform 1 0 1212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1711307567
transform 1 0 1164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1711307567
transform 1 0 1356 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1711307567
transform 1 0 1348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1711307567
transform 1 0 1172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1711307567
transform 1 0 1124 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1711307567
transform 1 0 1172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1711307567
transform 1 0 1172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1711307567
transform 1 0 1140 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1711307567
transform 1 0 1140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1711307567
transform 1 0 868 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1711307567
transform 1 0 868 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1711307567
transform 1 0 1308 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1711307567
transform 1 0 1268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1711307567
transform 1 0 1276 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1711307567
transform 1 0 1276 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1711307567
transform 1 0 1236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1711307567
transform 1 0 1204 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1711307567
transform 1 0 1172 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1711307567
transform 1 0 1108 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1711307567
transform 1 0 1100 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1711307567
transform 1 0 900 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1711307567
transform 1 0 900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1711307567
transform 1 0 1236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1711307567
transform 1 0 1228 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1711307567
transform 1 0 1140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1711307567
transform 1 0 1004 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1711307567
transform 1 0 1204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1711307567
transform 1 0 1116 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1711307567
transform 1 0 980 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1711307567
transform 1 0 1092 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1711307567
transform 1 0 1060 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1711307567
transform 1 0 1084 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1711307567
transform 1 0 948 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1711307567
transform 1 0 940 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1711307567
transform 1 0 1020 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1711307567
transform 1 0 988 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1711307567
transform 1 0 1332 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1711307567
transform 1 0 1316 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1711307567
transform 1 0 1452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1711307567
transform 1 0 1220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1711307567
transform 1 0 1212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1711307567
transform 1 0 1340 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1711307567
transform 1 0 1284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1711307567
transform 1 0 1156 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1711307567
transform 1 0 1308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1711307567
transform 1 0 1308 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1711307567
transform 1 0 1292 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1711307567
transform 1 0 1236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1711307567
transform 1 0 1132 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1711307567
transform 1 0 1236 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1711307567
transform 1 0 1236 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1711307567
transform 1 0 1596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1711307567
transform 1 0 1596 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1711307567
transform 1 0 1564 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1711307567
transform 1 0 1564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1711307567
transform 1 0 1580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1711307567
transform 1 0 1564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1711307567
transform 1 0 1532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1711307567
transform 1 0 1500 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1711307567
transform 1 0 1500 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1711307567
transform 1 0 1564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1711307567
transform 1 0 1540 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1711307567
transform 1 0 1668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1711307567
transform 1 0 1588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1711307567
transform 1 0 1588 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1711307567
transform 1 0 1556 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1711307567
transform 1 0 1516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1711307567
transform 1 0 1516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1711307567
transform 1 0 1980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1711307567
transform 1 0 1604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1711307567
transform 1 0 1596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1711307567
transform 1 0 1588 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1711307567
transform 1 0 1572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1711307567
transform 1 0 1556 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1711307567
transform 1 0 2292 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1711307567
transform 1 0 2108 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1711307567
transform 1 0 2084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1711307567
transform 1 0 1884 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1711307567
transform 1 0 1540 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1711307567
transform 1 0 1540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1711307567
transform 1 0 1508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1711307567
transform 1 0 1508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1711307567
transform 1 0 1580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1711307567
transform 1 0 1508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1711307567
transform 1 0 1524 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1711307567
transform 1 0 1444 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1711307567
transform 1 0 1452 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1711307567
transform 1 0 1444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1711307567
transform 1 0 2324 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1711307567
transform 1 0 2180 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1711307567
transform 1 0 2164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1711307567
transform 1 0 1596 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1711307567
transform 1 0 1572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1711307567
transform 1 0 1740 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1711307567
transform 1 0 1716 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1711307567
transform 1 0 1708 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1711307567
transform 1 0 1548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1711307567
transform 1 0 1748 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1711307567
transform 1 0 1700 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1711307567
transform 1 0 1772 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1711307567
transform 1 0 1764 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1711307567
transform 1 0 1652 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1711307567
transform 1 0 2244 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1711307567
transform 1 0 2212 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1711307567
transform 1 0 2092 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1711307567
transform 1 0 1628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1711307567
transform 1 0 1588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1711307567
transform 1 0 1900 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1711307567
transform 1 0 1724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1711307567
transform 1 0 1724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1711307567
transform 1 0 1716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1711307567
transform 1 0 1628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1711307567
transform 1 0 1716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1711307567
transform 1 0 1708 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1711307567
transform 1 0 1844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1711307567
transform 1 0 1772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1711307567
transform 1 0 1716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1711307567
transform 1 0 2396 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1711307567
transform 1 0 2284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1711307567
transform 1 0 1636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1711307567
transform 1 0 1628 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1711307567
transform 1 0 1860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1711307567
transform 1 0 1860 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1711307567
transform 1 0 1884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1711307567
transform 1 0 1796 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1711307567
transform 1 0 1924 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1711307567
transform 1 0 1692 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1711307567
transform 1 0 1684 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1711307567
transform 1 0 1860 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1711307567
transform 1 0 1828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1711307567
transform 1 0 1876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1711307567
transform 1 0 1852 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1711307567
transform 1 0 1772 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1711307567
transform 1 0 1772 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1711307567
transform 1 0 1772 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1711307567
transform 1 0 1812 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1711307567
transform 1 0 1796 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1711307567
transform 1 0 2196 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1711307567
transform 1 0 2108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1711307567
transform 1 0 1924 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1711307567
transform 1 0 1924 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1711307567
transform 1 0 2068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1711307567
transform 1 0 1996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1711307567
transform 1 0 1988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1711307567
transform 1 0 2116 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1711307567
transform 1 0 1972 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1711307567
transform 1 0 1956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1711307567
transform 1 0 2100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1711307567
transform 1 0 2084 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1711307567
transform 1 0 1964 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1711307567
transform 1 0 1932 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1711307567
transform 1 0 1916 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1711307567
transform 1 0 2004 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1711307567
transform 1 0 1988 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1711307567
transform 1 0 2220 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1711307567
transform 1 0 2188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1711307567
transform 1 0 1980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1711307567
transform 1 0 1916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1711307567
transform 1 0 2116 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1711307567
transform 1 0 2044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1711307567
transform 1 0 2028 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1711307567
transform 1 0 1972 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1711307567
transform 1 0 2124 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1711307567
transform 1 0 2124 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1711307567
transform 1 0 2052 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1711307567
transform 1 0 2172 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1711307567
transform 1 0 2068 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1711307567
transform 1 0 2196 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1711307567
transform 1 0 2180 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1711307567
transform 1 0 2020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1711307567
transform 1 0 1988 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1711307567
transform 1 0 1972 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1711307567
transform 1 0 2060 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1711307567
transform 1 0 2044 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1711307567
transform 1 0 1916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1711307567
transform 1 0 1852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1711307567
transform 1 0 1900 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1711307567
transform 1 0 1892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1711307567
transform 1 0 1940 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1711307567
transform 1 0 1908 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1711307567
transform 1 0 1852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1711307567
transform 1 0 1788 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1711307567
transform 1 0 1820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1711307567
transform 1 0 1820 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1711307567
transform 1 0 1836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1711307567
transform 1 0 1820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1711307567
transform 1 0 1924 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1711307567
transform 1 0 1908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1711307567
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1711307567
transform 1 0 1868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1711307567
transform 1 0 1828 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1711307567
transform 1 0 1756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1711307567
transform 1 0 2020 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1711307567
transform 1 0 2020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1711307567
transform 1 0 2012 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1711307567
transform 1 0 1988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1711307567
transform 1 0 1996 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1711307567
transform 1 0 1900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1711307567
transform 1 0 2196 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1711307567
transform 1 0 1980 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1711307567
transform 1 0 1844 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1711307567
transform 1 0 1980 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1711307567
transform 1 0 1964 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1711307567
transform 1 0 2012 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1711307567
transform 1 0 1972 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1711307567
transform 1 0 2036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1711307567
transform 1 0 1964 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1711307567
transform 1 0 2060 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1711307567
transform 1 0 2028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1711307567
transform 1 0 2228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1711307567
transform 1 0 2212 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1711307567
transform 1 0 2148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1711307567
transform 1 0 2140 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1711307567
transform 1 0 2084 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1711307567
transform 1 0 2036 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1711307567
transform 1 0 1972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1711307567
transform 1 0 1972 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1711307567
transform 1 0 1956 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1711307567
transform 1 0 2236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1711307567
transform 1 0 2236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1711307567
transform 1 0 2212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1711307567
transform 1 0 2084 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1711307567
transform 1 0 1844 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1711307567
transform 1 0 1620 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1711307567
transform 1 0 1556 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1711307567
transform 1 0 1508 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1711307567
transform 1 0 2244 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1711307567
transform 1 0 2140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1711307567
transform 1 0 1908 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1711307567
transform 1 0 2204 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1711307567
transform 1 0 2204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1711307567
transform 1 0 2196 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1711307567
transform 1 0 2196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1711307567
transform 1 0 2140 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1711307567
transform 1 0 2140 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1711307567
transform 1 0 2292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1711307567
transform 1 0 2268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1711307567
transform 1 0 2228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1711307567
transform 1 0 2156 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1711307567
transform 1 0 2268 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1711307567
transform 1 0 2268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1711307567
transform 1 0 2308 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1711307567
transform 1 0 2268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1711307567
transform 1 0 2220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1711307567
transform 1 0 2180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1711307567
transform 1 0 1884 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1711307567
transform 1 0 1580 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1711307567
transform 1 0 1524 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1711307567
transform 1 0 1476 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1711307567
transform 1 0 2244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1711307567
transform 1 0 2220 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1711307567
transform 1 0 2236 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1711307567
transform 1 0 2220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1711307567
transform 1 0 2092 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1711307567
transform 1 0 2092 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1711307567
transform 1 0 2076 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1711307567
transform 1 0 1980 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1711307567
transform 1 0 2076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1711307567
transform 1 0 2044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1711307567
transform 1 0 2204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1711307567
transform 1 0 2148 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1711307567
transform 1 0 2084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1711307567
transform 1 0 2108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1711307567
transform 1 0 2060 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1711307567
transform 1 0 2108 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1711307567
transform 1 0 2076 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1711307567
transform 1 0 2716 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1711307567
transform 1 0 2684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1711307567
transform 1 0 2644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1711307567
transform 1 0 2636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1711307567
transform 1 0 2596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1711307567
transform 1 0 2596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1711307567
transform 1 0 2660 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1711307567
transform 1 0 2628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1711307567
transform 1 0 2556 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1711307567
transform 1 0 2540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1711307567
transform 1 0 2596 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1711307567
transform 1 0 2580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1711307567
transform 1 0 2724 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1711307567
transform 1 0 2708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1711307567
transform 1 0 2652 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1711307567
transform 1 0 2572 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1711307567
transform 1 0 2572 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1711307567
transform 1 0 2564 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1711307567
transform 1 0 2564 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1711307567
transform 1 0 2580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1711307567
transform 1 0 2524 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1711307567
transform 1 0 2740 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1711307567
transform 1 0 2708 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1711307567
transform 1 0 2644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1711307567
transform 1 0 2636 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1711307567
transform 1 0 2604 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1711307567
transform 1 0 2572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1711307567
transform 1 0 2724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1711307567
transform 1 0 2676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1711307567
transform 1 0 2660 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1711307567
transform 1 0 2660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1711307567
transform 1 0 2620 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1711307567
transform 1 0 2588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1711307567
transform 1 0 2668 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1711307567
transform 1 0 2540 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1711307567
transform 1 0 2716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1711307567
transform 1 0 2596 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1711307567
transform 1 0 2652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1711307567
transform 1 0 2596 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1711307567
transform 1 0 2612 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1711307567
transform 1 0 2588 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1711307567
transform 1 0 2716 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1711307567
transform 1 0 2716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1711307567
transform 1 0 2588 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1711307567
transform 1 0 2540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1711307567
transform 1 0 2708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1711307567
transform 1 0 2572 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1711307567
transform 1 0 2724 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1711307567
transform 1 0 2604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1711307567
transform 1 0 2668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1711307567
transform 1 0 2628 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1711307567
transform 1 0 2628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1711307567
transform 1 0 2604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1711307567
transform 1 0 2412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1711307567
transform 1 0 2308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1711307567
transform 1 0 2356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1711307567
transform 1 0 2316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1711307567
transform 1 0 2292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1711307567
transform 1 0 2252 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1711307567
transform 1 0 2588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1711307567
transform 1 0 2588 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1711307567
transform 1 0 2388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1711307567
transform 1 0 2388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1711307567
transform 1 0 2212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1711307567
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1711307567
transform 1 0 2500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1711307567
transform 1 0 2500 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1711307567
transform 1 0 2644 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1711307567
transform 1 0 2644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1711307567
transform 1 0 2716 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1711307567
transform 1 0 2716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1711307567
transform 1 0 2044 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1711307567
transform 1 0 1948 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1711307567
transform 1 0 1988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1711307567
transform 1 0 1812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1711307567
transform 1 0 1908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1711307567
transform 1 0 1868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1711307567
transform 1 0 1860 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1711307567
transform 1 0 1828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1711307567
transform 1 0 1836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1711307567
transform 1 0 1796 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1711307567
transform 1 0 1804 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1711307567
transform 1 0 1740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1711307567
transform 1 0 1444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1711307567
transform 1 0 1444 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1711307567
transform 1 0 1364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1711307567
transform 1 0 1364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1711307567
transform 1 0 1676 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1711307567
transform 1 0 1596 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1711307567
transform 1 0 1228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1711307567
transform 1 0 1228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1711307567
transform 1 0 1092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1711307567
transform 1 0 1092 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1711307567
transform 1 0 1100 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1711307567
transform 1 0 1100 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1711307567
transform 1 0 1028 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1711307567
transform 1 0 908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1711307567
transform 1 0 1044 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1711307567
transform 1 0 972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1711307567
transform 1 0 588 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1711307567
transform 1 0 588 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1711307567
transform 1 0 740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1711307567
transform 1 0 732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1711307567
transform 1 0 772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1711307567
transform 1 0 684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1711307567
transform 1 0 468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1711307567
transform 1 0 460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1711307567
transform 1 0 540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1711307567
transform 1 0 540 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1711307567
transform 1 0 180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1711307567
transform 1 0 180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1711307567
transform 1 0 268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1711307567
transform 1 0 268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1711307567
transform 1 0 188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1711307567
transform 1 0 188 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1711307567
transform 1 0 108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1711307567
transform 1 0 108 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1711307567
transform 1 0 180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1711307567
transform 1 0 132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1711307567
transform 1 0 284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1711307567
transform 1 0 284 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1711307567
transform 1 0 2348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1711307567
transform 1 0 2300 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1711307567
transform 1 0 2308 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1711307567
transform 1 0 2252 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1711307567
transform 1 0 2252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1711307567
transform 1 0 2228 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1711307567
transform 1 0 2188 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1711307567
transform 1 0 2156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1711307567
transform 1 0 2076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1711307567
transform 1 0 1996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1711307567
transform 1 0 2236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1711307567
transform 1 0 2204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1711307567
transform 1 0 2196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1711307567
transform 1 0 2308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1711307567
transform 1 0 2268 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1711307567
transform 1 0 2220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1711307567
transform 1 0 2204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1711307567
transform 1 0 2164 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1711307567
transform 1 0 2484 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1711307567
transform 1 0 2140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1711307567
transform 1 0 2172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1711307567
transform 1 0 2132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1711307567
transform 1 0 2132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1711307567
transform 1 0 2116 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1711307567
transform 1 0 2084 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1711307567
transform 1 0 1956 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1711307567
transform 1 0 1884 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1711307567
transform 1 0 2172 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1711307567
transform 1 0 2132 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1711307567
transform 1 0 2076 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1711307567
transform 1 0 1964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1711307567
transform 1 0 2132 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1711307567
transform 1 0 2060 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1711307567
transform 1 0 2132 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1711307567
transform 1 0 2052 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1711307567
transform 1 0 2292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1711307567
transform 1 0 2268 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1711307567
transform 1 0 2244 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1711307567
transform 1 0 2228 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1711307567
transform 1 0 2004 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1711307567
transform 1 0 1988 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1711307567
transform 1 0 2148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1711307567
transform 1 0 2084 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1711307567
transform 1 0 2132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1711307567
transform 1 0 2132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1711307567
transform 1 0 2068 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1711307567
transform 1 0 2036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1711307567
transform 1 0 1980 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1711307567
transform 1 0 1980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1711307567
transform 1 0 1932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1711307567
transform 1 0 1932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1711307567
transform 1 0 1908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1711307567
transform 1 0 1908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1711307567
transform 1 0 2028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1711307567
transform 1 0 1980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1711307567
transform 1 0 2108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1711307567
transform 1 0 2100 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1711307567
transform 1 0 2116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1711307567
transform 1 0 1940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1711307567
transform 1 0 2180 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1711307567
transform 1 0 2180 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1711307567
transform 1 0 2012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1711307567
transform 1 0 1916 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1711307567
transform 1 0 2052 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1711307567
transform 1 0 2052 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1711307567
transform 1 0 1916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1711307567
transform 1 0 1812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1711307567
transform 1 0 1804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1711307567
transform 1 0 1796 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1711307567
transform 1 0 1916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1711307567
transform 1 0 1844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1711307567
transform 1 0 1820 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1711307567
transform 1 0 1780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1711307567
transform 1 0 1700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1711307567
transform 1 0 1492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1711307567
transform 1 0 1940 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1711307567
transform 1 0 1836 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1711307567
transform 1 0 1820 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1711307567
transform 1 0 1708 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1711307567
transform 1 0 1636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1711307567
transform 1 0 1636 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1711307567
transform 1 0 1972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1711307567
transform 1 0 1892 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1711307567
transform 1 0 1900 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1711307567
transform 1 0 1900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1711307567
transform 1 0 1860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1711307567
transform 1 0 1788 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1711307567
transform 1 0 1708 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1711307567
transform 1 0 1684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1711307567
transform 1 0 1548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1711307567
transform 1 0 2420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1711307567
transform 1 0 2364 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1711307567
transform 1 0 2356 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1711307567
transform 1 0 2268 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1711307567
transform 1 0 1732 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1711307567
transform 1 0 1580 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1711307567
transform 1 0 1828 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1711307567
transform 1 0 1660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1711307567
transform 1 0 1884 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1711307567
transform 1 0 1868 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1711307567
transform 1 0 1756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1711307567
transform 1 0 1652 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1711307567
transform 1 0 1508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1711307567
transform 1 0 1380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1711307567
transform 1 0 1748 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1711307567
transform 1 0 1724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1711307567
transform 1 0 1628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1711307567
transform 1 0 1628 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1711307567
transform 1 0 1908 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1711307567
transform 1 0 1652 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1711307567
transform 1 0 1500 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1711307567
transform 1 0 1492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1711307567
transform 1 0 1508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1711307567
transform 1 0 1508 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1711307567
transform 1 0 1772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1711307567
transform 1 0 1532 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1711307567
transform 1 0 1476 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1711307567
transform 1 0 1436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1711307567
transform 1 0 1428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1711307567
transform 1 0 1412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1711307567
transform 1 0 1836 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1711307567
transform 1 0 1468 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1711307567
transform 1 0 1620 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1711307567
transform 1 0 1612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1711307567
transform 1 0 1572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1711307567
transform 1 0 1572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1711307567
transform 1 0 1692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1711307567
transform 1 0 1564 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1711307567
transform 1 0 1500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1711307567
transform 1 0 1468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1711307567
transform 1 0 1468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1711307567
transform 1 0 1396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1711307567
transform 1 0 1364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1711307567
transform 1 0 1316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1711307567
transform 1 0 1244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1711307567
transform 1 0 1188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1711307567
transform 1 0 1180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1711307567
transform 1 0 1084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1711307567
transform 1 0 1428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1711307567
transform 1 0 1092 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1711307567
transform 1 0 996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1711307567
transform 1 0 940 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1711307567
transform 1 0 876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1711307567
transform 1 0 876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1711307567
transform 1 0 796 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1711307567
transform 1 0 756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1711307567
transform 1 0 1740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1711307567
transform 1 0 1732 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1711307567
transform 1 0 1716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1711307567
transform 1 0 1612 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1711307567
transform 1 0 1460 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1711307567
transform 1 0 1612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1711307567
transform 1 0 1596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1711307567
transform 1 0 1580 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1711307567
transform 1 0 1324 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1711307567
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1711307567
transform 1 0 1348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1711307567
transform 1 0 1284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1711307567
transform 1 0 1348 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1711307567
transform 1 0 1308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1711307567
transform 1 0 1420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1711307567
transform 1 0 1276 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1711307567
transform 1 0 1188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1711307567
transform 1 0 1172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1711307567
transform 1 0 1164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1711307567
transform 1 0 1252 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1711307567
transform 1 0 1252 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1711307567
transform 1 0 1308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1711307567
transform 1 0 1292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1711307567
transform 1 0 1308 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1711307567
transform 1 0 1236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1711307567
transform 1 0 1164 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1711307567
transform 1 0 1164 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1711307567
transform 1 0 1260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1711307567
transform 1 0 1156 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1711307567
transform 1 0 1244 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1711307567
transform 1 0 1180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1711307567
transform 1 0 1164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1711307567
transform 1 0 1036 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1711307567
transform 1 0 1204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1711307567
transform 1 0 1156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1711307567
transform 1 0 1196 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1711307567
transform 1 0 1172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1711307567
transform 1 0 1452 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1711307567
transform 1 0 1340 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1711307567
transform 1 0 1332 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1711307567
transform 1 0 1020 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1711307567
transform 1 0 1020 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1711307567
transform 1 0 1020 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1711307567
transform 1 0 924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1711307567
transform 1 0 916 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1711307567
transform 1 0 1076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1711307567
transform 1 0 1060 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1711307567
transform 1 0 964 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1711307567
transform 1 0 892 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1711307567
transform 1 0 892 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1711307567
transform 1 0 820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1711307567
transform 1 0 796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1711307567
transform 1 0 764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1711307567
transform 1 0 1388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1711307567
transform 1 0 1308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1711307567
transform 1 0 1172 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1711307567
transform 1 0 1108 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1711307567
transform 1 0 1076 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1711307567
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1711307567
transform 1 0 1556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1711307567
transform 1 0 1580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1711307567
transform 1 0 1548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1711307567
transform 1 0 1012 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1711307567
transform 1 0 1012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1711307567
transform 1 0 1012 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1711307567
transform 1 0 916 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1711307567
transform 1 0 692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1711307567
transform 1 0 692 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1711307567
transform 1 0 796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1711307567
transform 1 0 668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1711307567
transform 1 0 788 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1711307567
transform 1 0 772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1711307567
transform 1 0 772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1711307567
transform 1 0 772 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1711307567
transform 1 0 852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1711307567
transform 1 0 756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1711307567
transform 1 0 868 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1711307567
transform 1 0 860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1711307567
transform 1 0 900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1711307567
transform 1 0 892 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1711307567
transform 1 0 916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1711307567
transform 1 0 892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1711307567
transform 1 0 908 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1711307567
transform 1 0 844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1711307567
transform 1 0 876 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1711307567
transform 1 0 868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1711307567
transform 1 0 844 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1711307567
transform 1 0 796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1711307567
transform 1 0 892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1711307567
transform 1 0 876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1711307567
transform 1 0 900 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1711307567
transform 1 0 692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1711307567
transform 1 0 644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1711307567
transform 1 0 940 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1711307567
transform 1 0 612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1711307567
transform 1 0 612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1711307567
transform 1 0 956 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1711307567
transform 1 0 940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1711307567
transform 1 0 1516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1711307567
transform 1 0 948 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1711307567
transform 1 0 756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1711307567
transform 1 0 748 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1711307567
transform 1 0 700 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1711307567
transform 1 0 700 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1711307567
transform 1 0 492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1711307567
transform 1 0 492 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1711307567
transform 1 0 500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1711307567
transform 1 0 468 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1711307567
transform 1 0 708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1711307567
transform 1 0 532 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1711307567
transform 1 0 604 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1711307567
transform 1 0 596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1711307567
transform 1 0 564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1711307567
transform 1 0 548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1711307567
transform 1 0 660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1711307567
transform 1 0 580 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1711307567
transform 1 0 284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1711307567
transform 1 0 284 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1711307567
transform 1 0 420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1711307567
transform 1 0 300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1711307567
transform 1 0 588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1711307567
transform 1 0 452 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1711307567
transform 1 0 388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1711307567
transform 1 0 388 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1711307567
transform 1 0 460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1711307567
transform 1 0 364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1711307567
transform 1 0 620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1711307567
transform 1 0 468 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1711307567
transform 1 0 812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1711307567
transform 1 0 524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1711307567
transform 1 0 1316 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1711307567
transform 1 0 828 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1711307567
transform 1 0 812 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1711307567
transform 1 0 788 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1711307567
transform 1 0 772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1711307567
transform 1 0 332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1711307567
transform 1 0 284 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1711307567
transform 1 0 452 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1711307567
transform 1 0 340 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1711307567
transform 1 0 572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1711307567
transform 1 0 492 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1711307567
transform 1 0 492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1711307567
transform 1 0 436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1711307567
transform 1 0 436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1711307567
transform 1 0 628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1711307567
transform 1 0 564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1711307567
transform 1 0 564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1711307567
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1711307567
transform 1 0 468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1711307567
transform 1 0 292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1711307567
transform 1 0 244 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1711307567
transform 1 0 460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1711307567
transform 1 0 340 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1711307567
transform 1 0 332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1711307567
transform 1 0 308 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1711307567
transform 1 0 412 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1711307567
transform 1 0 348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1711307567
transform 1 0 548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1711307567
transform 1 0 436 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1711307567
transform 1 0 452 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1711307567
transform 1 0 428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1711307567
transform 1 0 396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1711307567
transform 1 0 372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1711307567
transform 1 0 548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1711307567
transform 1 0 428 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1711307567
transform 1 0 788 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1711307567
transform 1 0 612 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1711307567
transform 1 0 588 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1711307567
transform 1 0 372 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1711307567
transform 1 0 356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1711307567
transform 1 0 2660 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1711307567
transform 1 0 2628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1711307567
transform 1 0 2580 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1711307567
transform 1 0 2572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1711307567
transform 1 0 2596 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1711307567
transform 1 0 2596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1711307567
transform 1 0 2556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1711307567
transform 1 0 2556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1711307567
transform 1 0 2532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1711307567
transform 1 0 2468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1711307567
transform 1 0 2452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1711307567
transform 1 0 2452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1711307567
transform 1 0 2468 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1711307567
transform 1 0 2436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1711307567
transform 1 0 2620 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1711307567
transform 1 0 2540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1711307567
transform 1 0 2548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1711307567
transform 1 0 2436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1711307567
transform 1 0 2372 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1711307567
transform 1 0 2364 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1711307567
transform 1 0 1532 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1711307567
transform 1 0 2404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1711307567
transform 1 0 2388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1711307567
transform 1 0 2628 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1711307567
transform 1 0 2532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1711307567
transform 1 0 2540 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1711307567
transform 1 0 2428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1711307567
transform 1 0 2388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1711307567
transform 1 0 2372 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1711307567
transform 1 0 1508 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1711307567
transform 1 0 1508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1711307567
transform 1 0 1564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1711307567
transform 1 0 1524 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1711307567
transform 1 0 1564 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1711307567
transform 1 0 1340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1711307567
transform 1 0 2460 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1711307567
transform 1 0 2180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1711307567
transform 1 0 1940 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1711307567
transform 1 0 764 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1711307567
transform 1 0 748 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1711307567
transform 1 0 308 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1711307567
transform 1 0 276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1711307567
transform 1 0 804 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1711307567
transform 1 0 796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1711307567
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1711307567
transform 1 0 1164 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1711307567
transform 1 0 1068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1711307567
transform 1 0 1012 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1711307567
transform 1 0 1916 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1711307567
transform 1 0 1908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1711307567
transform 1 0 2340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1711307567
transform 1 0 2260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1711307567
transform 1 0 2388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1711307567
transform 1 0 2308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1711307567
transform 1 0 2388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1711307567
transform 1 0 2300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1711307567
transform 1 0 2524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1711307567
transform 1 0 2484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1711307567
transform 1 0 2116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1711307567
transform 1 0 2004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1711307567
transform 1 0 2060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1711307567
transform 1 0 2060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1711307567
transform 1 0 2068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1711307567
transform 1 0 2068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1711307567
transform 1 0 2156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1711307567
transform 1 0 2156 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1711307567
transform 1 0 2004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1711307567
transform 1 0 2004 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1711307567
transform 1 0 1756 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1711307567
transform 1 0 1684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1711307567
transform 1 0 1564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1711307567
transform 1 0 1500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1711307567
transform 1 0 1476 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1711307567
transform 1 0 1412 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1711307567
transform 1 0 1620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1711307567
transform 1 0 1524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1711307567
transform 1 0 1324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1711307567
transform 1 0 1316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1711307567
transform 1 0 1316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1711307567
transform 1 0 1276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1711307567
transform 1 0 1180 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1711307567
transform 1 0 1180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1711307567
transform 1 0 1020 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1711307567
transform 1 0 980 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1711307567
transform 1 0 988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1711307567
transform 1 0 980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1711307567
transform 1 0 692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1711307567
transform 1 0 684 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1711307567
transform 1 0 812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1711307567
transform 1 0 812 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1711307567
transform 1 0 892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1711307567
transform 1 0 852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1711307567
transform 1 0 484 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1711307567
transform 1 0 436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1711307567
transform 1 0 604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1711307567
transform 1 0 564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1711307567
transform 1 0 244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1711307567
transform 1 0 196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1711307567
transform 1 0 364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1711307567
transform 1 0 316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1711307567
transform 1 0 260 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1711307567
transform 1 0 132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1711307567
transform 1 0 228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1711307567
transform 1 0 124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1711307567
transform 1 0 236 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1711307567
transform 1 0 132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1711307567
transform 1 0 444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1711307567
transform 1 0 396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1711307567
transform 1 0 2700 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1711307567
transform 1 0 2660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1711307567
transform 1 0 2636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1711307567
transform 1 0 2636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1711307567
transform 1 0 2700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1711307567
transform 1 0 2620 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1711307567
transform 1 0 2700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1711307567
transform 1 0 2628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1711307567
transform 1 0 2652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1711307567
transform 1 0 2548 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1711307567
transform 1 0 2492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1711307567
transform 1 0 2436 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1711307567
transform 1 0 2180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1711307567
transform 1 0 2140 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1711307567
transform 1 0 2700 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1711307567
transform 1 0 2660 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1711307567
transform 1 0 2692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1711307567
transform 1 0 2660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1711307567
transform 1 0 2628 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1711307567
transform 1 0 2556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1711307567
transform 1 0 2620 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1711307567
transform 1 0 2588 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1711307567
transform 1 0 2604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1711307567
transform 1 0 2604 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1711307567
transform 1 0 2620 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1711307567
transform 1 0 2604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1711307567
transform 1 0 2412 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1711307567
transform 1 0 2140 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1711307567
transform 1 0 2500 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1711307567
transform 1 0 2484 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1711307567
transform 1 0 2460 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1711307567
transform 1 0 2452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1711307567
transform 1 0 2540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1711307567
transform 1 0 2476 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1711307567
transform 1 0 2476 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1711307567
transform 1 0 2420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1711307567
transform 1 0 2244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1711307567
transform 1 0 2244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1711307567
transform 1 0 2636 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1711307567
transform 1 0 2620 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1711307567
transform 1 0 2620 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1711307567
transform 1 0 2284 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1711307567
transform 1 0 2268 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1711307567
transform 1 0 1732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1711307567
transform 1 0 1668 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1711307567
transform 1 0 1292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1711307567
transform 1 0 2540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1711307567
transform 1 0 2508 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1711307567
transform 1 0 2412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1711307567
transform 1 0 2412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1711307567
transform 1 0 2340 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1711307567
transform 1 0 1964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1711307567
transform 1 0 1876 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1711307567
transform 1 0 1740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1711307567
transform 1 0 1732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1711307567
transform 1 0 1156 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1711307567
transform 1 0 1068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1711307567
transform 1 0 996 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1711307567
transform 1 0 884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1711307567
transform 1 0 1740 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1711307567
transform 1 0 1724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1711307567
transform 1 0 1684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1711307567
transform 1 0 1332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1711307567
transform 1 0 1884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1711307567
transform 1 0 1868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1711307567
transform 1 0 2404 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1711307567
transform 1 0 2332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1711307567
transform 1 0 2532 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1711307567
transform 1 0 2476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1711307567
transform 1 0 2404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1711307567
transform 1 0 2268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1711307567
transform 1 0 1972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1711307567
transform 1 0 1948 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1711307567
transform 1 0 1916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1711307567
transform 1 0 380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1711307567
transform 1 0 372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1711307567
transform 1 0 308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1711307567
transform 1 0 292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1711307567
transform 1 0 292 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1711307567
transform 1 0 228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1711307567
transform 1 0 220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1711307567
transform 1 0 2204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1711307567
transform 1 0 2172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1711307567
transform 1 0 2172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1711307567
transform 1 0 284 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1711307567
transform 1 0 276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1711307567
transform 1 0 268 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1711307567
transform 1 0 148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1711307567
transform 1 0 300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1711307567
transform 1 0 268 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1711307567
transform 1 0 252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1711307567
transform 1 0 228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1711307567
transform 1 0 436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1711307567
transform 1 0 428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1711307567
transform 1 0 324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1711307567
transform 1 0 476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1711307567
transform 1 0 356 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1711307567
transform 1 0 204 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1711307567
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1711307567
transform 1 0 508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1711307567
transform 1 0 460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1711307567
transform 1 0 396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1711307567
transform 1 0 548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1711307567
transform 1 0 484 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1711307567
transform 1 0 484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1711307567
transform 1 0 476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1711307567
transform 1 0 476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1711307567
transform 1 0 708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1711307567
transform 1 0 692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1711307567
transform 1 0 676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1711307567
transform 1 0 620 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1711307567
transform 1 0 604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1711307567
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1711307567
transform 1 0 988 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1711307567
transform 1 0 916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1711307567
transform 1 0 900 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1711307567
transform 1 0 2636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1711307567
transform 1 0 2332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1711307567
transform 1 0 2316 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1711307567
transform 1 0 2220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1711307567
transform 1 0 916 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1711307567
transform 1 0 876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1711307567
transform 1 0 1060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1711307567
transform 1 0 956 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1711307567
transform 1 0 940 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1711307567
transform 1 0 924 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1711307567
transform 1 0 924 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1711307567
transform 1 0 1172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1711307567
transform 1 0 1148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1711307567
transform 1 0 1276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1711307567
transform 1 0 1252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1711307567
transform 1 0 1548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1711307567
transform 1 0 1444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1711307567
transform 1 0 1076 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1711307567
transform 1 0 884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1711307567
transform 1 0 1380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1711307567
transform 1 0 1260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1711307567
transform 1 0 1108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1711307567
transform 1 0 828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1711307567
transform 1 0 1484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1711307567
transform 1 0 1388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1711307567
transform 1 0 1204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1711307567
transform 1 0 1204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1711307567
transform 1 0 740 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1711307567
transform 1 0 1620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1711307567
transform 1 0 1604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1711307567
transform 1 0 1500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1711307567
transform 1 0 1252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1711307567
transform 1 0 1180 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1711307567
transform 1 0 996 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1711307567
transform 1 0 1676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1711307567
transform 1 0 1644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1711307567
transform 1 0 1604 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1711307567
transform 1 0 1564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1711307567
transform 1 0 1180 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1711307567
transform 1 0 1780 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1711307567
transform 1 0 1780 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1711307567
transform 1 0 1660 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1711307567
transform 1 0 1644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1711307567
transform 1 0 1628 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1711307567
transform 1 0 1220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1711307567
transform 1 0 2156 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1711307567
transform 1 0 2100 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1711307567
transform 1 0 2076 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1711307567
transform 1 0 2404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1711307567
transform 1 0 2404 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1711307567
transform 1 0 2452 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1711307567
transform 1 0 1516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1711307567
transform 1 0 2228 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1711307567
transform 1 0 2212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1711307567
transform 1 0 2212 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1711307567
transform 1 0 2172 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1711307567
transform 1 0 2140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1711307567
transform 1 0 2108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1711307567
transform 1 0 2108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1711307567
transform 1 0 2308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1711307567
transform 1 0 2276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1711307567
transform 1 0 2260 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1711307567
transform 1 0 2100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1711307567
transform 1 0 2556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1711307567
transform 1 0 2308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1711307567
transform 1 0 2260 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1711307567
transform 1 0 2236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1711307567
transform 1 0 2204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1711307567
transform 1 0 2204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1711307567
transform 1 0 2172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1711307567
transform 1 0 2212 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1711307567
transform 1 0 2188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1711307567
transform 1 0 2020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1711307567
transform 1 0 2020 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1711307567
transform 1 0 2020 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1711307567
transform 1 0 2244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1711307567
transform 1 0 2156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1711307567
transform 1 0 2148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1711307567
transform 1 0 1980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1711307567
transform 1 0 1892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1711307567
transform 1 0 1884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1711307567
transform 1 0 2484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1711307567
transform 1 0 2476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1711307567
transform 1 0 2444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1711307567
transform 1 0 2116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1711307567
transform 1 0 2100 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1711307567
transform 1 0 1892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1711307567
transform 1 0 1756 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1711307567
transform 1 0 2468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1711307567
transform 1 0 2340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1711307567
transform 1 0 2188 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1711307567
transform 1 0 1924 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1711307567
transform 1 0 1908 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1711307567
transform 1 0 1820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1711307567
transform 1 0 2068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1711307567
transform 1 0 2060 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1711307567
transform 1 0 1924 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1711307567
transform 1 0 1916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1711307567
transform 1 0 1780 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1711307567
transform 1 0 1676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1711307567
transform 1 0 1924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1711307567
transform 1 0 1740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1711307567
transform 1 0 1716 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1711307567
transform 1 0 1940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1711307567
transform 1 0 1804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1711307567
transform 1 0 1732 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1711307567
transform 1 0 1708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1711307567
transform 1 0 1708 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1711307567
transform 1 0 1884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1711307567
transform 1 0 1884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1711307567
transform 1 0 1852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1711307567
transform 1 0 1844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1711307567
transform 1 0 1876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1711307567
transform 1 0 1708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1711307567
transform 1 0 1668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1711307567
transform 1 0 1348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1711307567
transform 1 0 1284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1711307567
transform 1 0 1260 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1711307567
transform 1 0 1252 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1711307567
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1711307567
transform 1 0 1228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1711307567
transform 1 0 1196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1711307567
transform 1 0 1180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1711307567
transform 1 0 1140 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1711307567
transform 1 0 1140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1711307567
transform 1 0 1212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1711307567
transform 1 0 1148 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1711307567
transform 1 0 1132 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1711307567
transform 1 0 1124 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1711307567
transform 1 0 1108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1711307567
transform 1 0 1292 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1711307567
transform 1 0 1284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1711307567
transform 1 0 1252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1711307567
transform 1 0 1044 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1711307567
transform 1 0 900 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1711307567
transform 1 0 700 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1711307567
transform 1 0 1220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1711307567
transform 1 0 1180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1711307567
transform 1 0 1116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1711307567
transform 1 0 1100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1711307567
transform 1 0 1076 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1711307567
transform 1 0 1052 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1711307567
transform 1 0 756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1711307567
transform 1 0 652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1711307567
transform 1 0 1116 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1711307567
transform 1 0 940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1711307567
transform 1 0 828 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1711307567
transform 1 0 572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1711307567
transform 1 0 1156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1711307567
transform 1 0 1004 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1711307567
transform 1 0 1004 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1711307567
transform 1 0 972 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1711307567
transform 1 0 964 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1711307567
transform 1 0 932 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1711307567
transform 1 0 804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1711307567
transform 1 0 612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1711307567
transform 1 0 924 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1711307567
transform 1 0 924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1711307567
transform 1 0 732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1711307567
transform 1 0 716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1711307567
transform 1 0 444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1711307567
transform 1 0 780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1711307567
transform 1 0 780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1711307567
transform 1 0 780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1711307567
transform 1 0 684 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1711307567
transform 1 0 540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1711307567
transform 1 0 452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1711307567
transform 1 0 868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1711307567
transform 1 0 844 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1711307567
transform 1 0 812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1711307567
transform 1 0 596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1711307567
transform 1 0 596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1711307567
transform 1 0 572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1711307567
transform 1 0 540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1711307567
transform 1 0 852 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1711307567
transform 1 0 804 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1711307567
transform 1 0 724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1711307567
transform 1 0 700 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1711307567
transform 1 0 628 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1711307567
transform 1 0 540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1711307567
transform 1 0 476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1711307567
transform 1 0 460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1711307567
transform 1 0 484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1711307567
transform 1 0 468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1711307567
transform 1 0 436 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1711307567
transform 1 0 580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1711307567
transform 1 0 572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1711307567
transform 1 0 556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1711307567
transform 1 0 500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1711307567
transform 1 0 556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1711307567
transform 1 0 540 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1711307567
transform 1 0 476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1711307567
transform 1 0 468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1711307567
transform 1 0 260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1711307567
transform 1 0 252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1711307567
transform 1 0 284 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1711307567
transform 1 0 284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1711307567
transform 1 0 396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1711307567
transform 1 0 388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1711307567
transform 1 0 356 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1711307567
transform 1 0 2668 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1711307567
transform 1 0 2652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1711307567
transform 1 0 2724 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1711307567
transform 1 0 2708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1711307567
transform 1 0 2468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1711307567
transform 1 0 2452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1711307567
transform 1 0 1500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1711307567
transform 1 0 1476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1711307567
transform 1 0 2692 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1711307567
transform 1 0 2676 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1711307567
transform 1 0 2676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1711307567
transform 1 0 2604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1711307567
transform 1 0 2500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1711307567
transform 1 0 2356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1711307567
transform 1 0 2356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1711307567
transform 1 0 2332 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1711307567
transform 1 0 2700 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1711307567
transform 1 0 2604 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1711307567
transform 1 0 2532 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1711307567
transform 1 0 2372 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1711307567
transform 1 0 2340 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1711307567
transform 1 0 2316 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1711307567
transform 1 0 2516 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1711307567
transform 1 0 2412 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1711307567
transform 1 0 2380 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1711307567
transform 1 0 2372 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1711307567
transform 1 0 2308 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1711307567
transform 1 0 2284 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1711307567
transform 1 0 2452 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1711307567
transform 1 0 2396 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1711307567
transform 1 0 2364 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1711307567
transform 1 0 2348 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1711307567
transform 1 0 2348 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1711307567
transform 1 0 2284 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1711307567
transform 1 0 2388 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1711307567
transform 1 0 2076 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1711307567
transform 1 0 1988 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1711307567
transform 1 0 2292 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1711307567
transform 1 0 2084 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1711307567
transform 1 0 1996 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1711307567
transform 1 0 2324 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1711307567
transform 1 0 2276 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1711307567
transform 1 0 2076 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1711307567
transform 1 0 2060 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1711307567
transform 1 0 2004 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1711307567
transform 1 0 1964 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1711307567
transform 1 0 1852 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1711307567
transform 1 0 2540 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1711307567
transform 1 0 2420 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1711307567
transform 1 0 2124 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1711307567
transform 1 0 2084 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1711307567
transform 1 0 1996 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1711307567
transform 1 0 1964 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1711307567
transform 1 0 1916 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1711307567
transform 1 0 2452 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1711307567
transform 1 0 2172 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1711307567
transform 1 0 1700 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1711307567
transform 1 0 1332 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1711307567
transform 1 0 2484 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1711307567
transform 1 0 2100 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1711307567
transform 1 0 2100 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1711307567
transform 1 0 1724 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1711307567
transform 1 0 1372 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1711307567
transform 1 0 1372 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1711307567
transform 1 0 1308 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1711307567
transform 1 0 2548 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1711307567
transform 1 0 2332 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1711307567
transform 1 0 2260 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1711307567
transform 1 0 2436 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1711307567
transform 1 0 2316 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1711307567
transform 1 0 2756 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1711307567
transform 1 0 2596 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1711307567
transform 1 0 2684 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1711307567
transform 1 0 2588 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1711307567
transform 1 0 2436 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1711307567
transform 1 0 2308 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1711307567
transform 1 0 2580 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1711307567
transform 1 0 2516 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1711307567
transform 1 0 2756 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1711307567
transform 1 0 2628 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1711307567
transform 1 0 2756 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1711307567
transform 1 0 2620 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1711307567
transform 1 0 2124 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1711307567
transform 1 0 2028 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1711307567
transform 1 0 2108 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1711307567
transform 1 0 1988 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1711307567
transform 1 0 2196 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1711307567
transform 1 0 1956 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1711307567
transform 1 0 1868 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1711307567
transform 1 0 2036 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1711307567
transform 1 0 1932 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1711307567
transform 1 0 1612 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1711307567
transform 1 0 1508 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1711307567
transform 1 0 1348 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1711307567
transform 1 0 1260 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1711307567
transform 1 0 1380 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1711307567
transform 1 0 1212 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1711307567
transform 1 0 1236 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1711307567
transform 1 0 1100 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1711307567
transform 1 0 716 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1711307567
transform 1 0 628 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1711307567
transform 1 0 860 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1711307567
transform 1 0 748 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1711307567
transform 1 0 900 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1711307567
transform 1 0 804 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1711307567
transform 1 0 596 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1711307567
transform 1 0 532 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1711307567
transform 1 0 188 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1711307567
transform 1 0 92 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1711307567
transform 1 0 428 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1711307567
transform 1 0 364 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1711307567
transform 1 0 2756 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1711307567
transform 1 0 2660 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1711307567
transform 1 0 2284 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1711307567
transform 1 0 2084 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1711307567
transform 1 0 2628 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1711307567
transform 1 0 2324 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1711307567
transform 1 0 2444 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1711307567
transform 1 0 2188 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1711307567
transform 1 0 2204 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1711307567
transform 1 0 1940 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1711307567
transform 1 0 2540 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1711307567
transform 1 0 2388 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1711307567
transform 1 0 2676 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1711307567
transform 1 0 2524 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1711307567
transform 1 0 2756 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1711307567
transform 1 0 2388 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1711307567
transform 1 0 1972 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1711307567
transform 1 0 1852 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1711307567
transform 1 0 1868 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1711307567
transform 1 0 1708 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1711307567
transform 1 0 1900 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1711307567
transform 1 0 1716 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1711307567
transform 1 0 1860 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1711307567
transform 1 0 1756 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1711307567
transform 1 0 1844 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1711307567
transform 1 0 1596 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1711307567
transform 1 0 1860 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1711307567
transform 1 0 1764 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1711307567
transform 1 0 1764 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1711307567
transform 1 0 1604 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1711307567
transform 1 0 1476 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1711307567
transform 1 0 1364 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1711307567
transform 1 0 1372 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1711307567
transform 1 0 1220 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1711307567
transform 1 0 1708 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1711307567
transform 1 0 1524 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1711307567
transform 1 0 1524 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1711307567
transform 1 0 1428 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1711307567
transform 1 0 1124 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1711307567
transform 1 0 1036 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1711307567
transform 1 0 988 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1711307567
transform 1 0 860 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1711307567
transform 1 0 1028 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1711307567
transform 1 0 972 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1711307567
transform 1 0 748 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1711307567
transform 1 0 708 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1711307567
transform 1 0 724 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1711307567
transform 1 0 676 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1711307567
transform 1 0 516 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1711307567
transform 1 0 460 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1711307567
transform 1 0 596 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1711307567
transform 1 0 380 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1711307567
transform 1 0 220 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1711307567
transform 1 0 188 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1711307567
transform 1 0 340 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1711307567
transform 1 0 308 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1711307567
transform 1 0 220 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1711307567
transform 1 0 188 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1711307567
transform 1 0 316 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1711307567
transform 1 0 268 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1711307567
transform 1 0 2060 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1711307567
transform 1 0 1972 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1711307567
transform 1 0 2420 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1711307567
transform 1 0 2332 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1711307567
transform 1 0 1468 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1711307567
transform 1 0 1436 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1711307567
transform 1 0 1164 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1711307567
transform 1 0 1140 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1711307567
transform 1 0 948 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1711307567
transform 1 0 892 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1711307567
transform 1 0 844 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1711307567
transform 1 0 708 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1711307567
transform 1 0 572 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1711307567
transform 1 0 532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1711307567
transform 1 0 212 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1711307567
transform 1 0 212 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1711307567
transform 1 0 188 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1711307567
transform 1 0 188 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1711307567
transform 1 0 388 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1711307567
transform 1 0 356 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1711307567
transform 1 0 244 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1711307567
transform 1 0 204 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1711307567
transform 1 0 332 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1711307567
transform 1 0 196 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1711307567
transform 1 0 2548 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1711307567
transform 1 0 2500 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1711307567
transform 1 0 2676 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1711307567
transform 1 0 2644 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1711307567
transform 1 0 2628 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1711307567
transform 1 0 2684 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1711307567
transform 1 0 2652 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1711307567
transform 1 0 2644 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1711307567
transform 1 0 2620 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1711307567
transform 1 0 2556 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1711307567
transform 1 0 2644 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1711307567
transform 1 0 2604 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1711307567
transform 1 0 2500 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1711307567
transform 1 0 2476 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1711307567
transform 1 0 2436 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1711307567
transform 1 0 2436 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1711307567
transform 1 0 2684 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1711307567
transform 1 0 2604 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1711307567
transform 1 0 2452 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1711307567
transform 1 0 2420 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1711307567
transform 1 0 2700 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1711307567
transform 1 0 2644 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1711307567
transform 1 0 2612 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1711307567
transform 1 0 2460 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1711307567
transform 1 0 2372 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1711307567
transform 1 0 2660 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1711307567
transform 1 0 2532 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1711307567
transform 1 0 2284 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1711307567
transform 1 0 2596 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1711307567
transform 1 0 2524 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1711307567
transform 1 0 2492 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1711307567
transform 1 0 2388 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1711307567
transform 1 0 2348 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1711307567
transform 1 0 2252 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1711307567
transform 1 0 2708 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1711307567
transform 1 0 2540 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1711307567
transform 1 0 2460 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1711307567
transform 1 0 2284 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1711307567
transform 1 0 2756 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1711307567
transform 1 0 2572 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1711307567
transform 1 0 2572 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1711307567
transform 1 0 2524 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1711307567
transform 1 0 2484 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1711307567
transform 1 0 2356 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1711307567
transform 1 0 2284 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1711307567
transform 1 0 2756 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1711307567
transform 1 0 2628 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1711307567
transform 1 0 2620 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1711307567
transform 1 0 2596 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1711307567
transform 1 0 2756 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1711307567
transform 1 0 2644 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1711307567
transform 1 0 2380 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1711307567
transform 1 0 2332 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1711307567
transform 1 0 2308 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1711307567
transform 1 0 1876 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1711307567
transform 1 0 1852 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1711307567
transform 1 0 1780 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1711307567
transform 1 0 1780 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1711307567
transform 1 0 1668 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1711307567
transform 1 0 1644 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1711307567
transform 1 0 1628 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1711307567
transform 1 0 1588 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1711307567
transform 1 0 1588 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1711307567
transform 1 0 1556 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1711307567
transform 1 0 1188 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1711307567
transform 1 0 1156 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1711307567
transform 1 0 540 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1711307567
transform 1 0 532 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1711307567
transform 1 0 508 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1711307567
transform 1 0 492 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1711307567
transform 1 0 1028 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1711307567
transform 1 0 980 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1711307567
transform 1 0 820 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1711307567
transform 1 0 820 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1711307567
transform 1 0 764 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1711307567
transform 1 0 748 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1711307567
transform 1 0 660 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1711307567
transform 1 0 644 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1711307567
transform 1 0 524 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1711307567
transform 1 0 1492 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1711307567
transform 1 0 1428 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1711307567
transform 1 0 1924 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1711307567
transform 1 0 1868 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1711307567
transform 1 0 1644 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1711307567
transform 1 0 860 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1711307567
transform 1 0 860 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1711307567
transform 1 0 836 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1711307567
transform 1 0 2036 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1711307567
transform 1 0 1932 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1711307567
transform 1 0 1932 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1711307567
transform 1 0 1852 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1711307567
transform 1 0 1828 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1711307567
transform 1 0 1972 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1711307567
transform 1 0 1892 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1711307567
transform 1 0 1892 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1711307567
transform 1 0 1820 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1711307567
transform 1 0 1892 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1711307567
transform 1 0 1812 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1711307567
transform 1 0 1676 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1711307567
transform 1 0 996 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1711307567
transform 1 0 788 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1711307567
transform 1 0 956 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1711307567
transform 1 0 916 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1711307567
transform 1 0 1932 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1711307567
transform 1 0 1612 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1711307567
transform 1 0 1612 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1711307567
transform 1 0 1524 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1711307567
transform 1 0 1444 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1711307567
transform 1 0 1436 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1711307567
transform 1 0 836 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1711307567
transform 1 0 1676 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1711307567
transform 1 0 1412 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1711307567
transform 1 0 1076 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1711307567
transform 1 0 1076 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1711307567
transform 1 0 524 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1711307567
transform 1 0 1052 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1711307567
transform 1 0 1028 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1711307567
transform 1 0 860 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1711307567
transform 1 0 860 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1711307567
transform 1 0 772 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1711307567
transform 1 0 1900 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1711307567
transform 1 0 1788 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1711307567
transform 1 0 1748 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1711307567
transform 1 0 1252 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1711307567
transform 1 0 1516 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1711307567
transform 1 0 1436 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1711307567
transform 1 0 1388 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1711307567
transform 1 0 1388 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1711307567
transform 1 0 1340 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1711307567
transform 1 0 1308 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1711307567
transform 1 0 1916 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1711307567
transform 1 0 1844 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1711307567
transform 1 0 1508 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1711307567
transform 1 0 1316 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1711307567
transform 1 0 1228 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1711307567
transform 1 0 1604 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1711307567
transform 1 0 564 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1711307567
transform 1 0 380 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1711307567
transform 1 0 356 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1711307567
transform 1 0 316 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1711307567
transform 1 0 1660 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1711307567
transform 1 0 1620 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1711307567
transform 1 0 1332 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1711307567
transform 1 0 1132 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1711307567
transform 1 0 1604 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1711307567
transform 1 0 1572 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1711307567
transform 1 0 628 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1711307567
transform 1 0 628 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1711307567
transform 1 0 484 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1711307567
transform 1 0 1748 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1711307567
transform 1 0 1716 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1711307567
transform 1 0 1460 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1711307567
transform 1 0 1388 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1711307567
transform 1 0 1828 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1711307567
transform 1 0 1388 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1711307567
transform 1 0 988 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1711307567
transform 1 0 988 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1711307567
transform 1 0 540 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1711307567
transform 1 0 412 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1711307567
transform 1 0 412 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1711307567
transform 1 0 388 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1711307567
transform 1 0 572 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1711307567
transform 1 0 532 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1711307567
transform 1 0 484 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1711307567
transform 1 0 468 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1711307567
transform 1 0 1156 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1711307567
transform 1 0 1108 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1711307567
transform 1 0 900 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1711307567
transform 1 0 2028 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1711307567
transform 1 0 1748 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1711307567
transform 1 0 1412 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1711307567
transform 1 0 1388 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1711307567
transform 1 0 1084 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1711307567
transform 1 0 1356 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1711307567
transform 1 0 1148 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1711307567
transform 1 0 1060 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1711307567
transform 1 0 1692 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1711307567
transform 1 0 1588 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1711307567
transform 1 0 1236 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1711307567
transform 1 0 780 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1711307567
transform 1 0 524 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1711307567
transform 1 0 836 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1711307567
transform 1 0 748 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1711307567
transform 1 0 2116 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1711307567
transform 1 0 2044 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1711307567
transform 1 0 2036 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1711307567
transform 1 0 1988 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1711307567
transform 1 0 1396 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1711307567
transform 1 0 1396 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1711307567
transform 1 0 1252 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1711307567
transform 1 0 1044 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1711307567
transform 1 0 1004 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1711307567
transform 1 0 980 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1711307567
transform 1 0 1716 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1711307567
transform 1 0 1668 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1711307567
transform 1 0 812 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1711307567
transform 1 0 636 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1711307567
transform 1 0 532 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1711307567
transform 1 0 508 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1711307567
transform 1 0 1788 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1711307567
transform 1 0 1716 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1711307567
transform 1 0 1724 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1711307567
transform 1 0 1692 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1711307567
transform 1 0 1596 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1711307567
transform 1 0 1260 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1711307567
transform 1 0 1260 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1711307567
transform 1 0 1180 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1711307567
transform 1 0 732 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1711307567
transform 1 0 708 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1711307567
transform 1 0 588 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1711307567
transform 1 0 548 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1711307567
transform 1 0 1140 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1711307567
transform 1 0 988 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1711307567
transform 1 0 988 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1711307567
transform 1 0 820 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1711307567
transform 1 0 812 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1711307567
transform 1 0 764 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1711307567
transform 1 0 1980 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1711307567
transform 1 0 1876 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1711307567
transform 1 0 2332 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1711307567
transform 1 0 2268 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1711307567
transform 1 0 2228 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1711307567
transform 1 0 2388 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1711307567
transform 1 0 2292 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1711307567
transform 1 0 2220 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1711307567
transform 1 0 1108 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1711307567
transform 1 0 1028 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1711307567
transform 1 0 956 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1711307567
transform 1 0 1748 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1711307567
transform 1 0 1692 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1711307567
transform 1 0 2252 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1711307567
transform 1 0 2036 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1711307567
transform 1 0 1188 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1711307567
transform 1 0 820 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1711307567
transform 1 0 572 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1711307567
transform 1 0 2172 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1711307567
transform 1 0 2004 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1711307567
transform 1 0 2004 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1711307567
transform 1 0 1684 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1711307567
transform 1 0 1132 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1711307567
transform 1 0 612 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1711307567
transform 1 0 1900 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1711307567
transform 1 0 1804 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1711307567
transform 1 0 1796 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1711307567
transform 1 0 1220 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1711307567
transform 1 0 820 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1711307567
transform 1 0 1700 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1711307567
transform 1 0 1668 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1711307567
transform 1 0 2364 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1711307567
transform 1 0 2284 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1711307567
transform 1 0 2252 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1711307567
transform 1 0 2252 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1711307567
transform 1 0 2092 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1711307567
transform 1 0 1916 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1711307567
transform 1 0 1708 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1711307567
transform 1 0 844 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1711307567
transform 1 0 716 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1711307567
transform 1 0 1668 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1711307567
transform 1 0 1628 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1711307567
transform 1 0 1964 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1711307567
transform 1 0 1892 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1711307567
transform 1 0 1236 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1711307567
transform 1 0 1236 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1711307567
transform 1 0 1188 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1711307567
transform 1 0 852 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1711307567
transform 1 0 2276 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1711307567
transform 1 0 2036 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1711307567
transform 1 0 1228 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1711307567
transform 1 0 1228 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1711307567
transform 1 0 788 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1711307567
transform 1 0 596 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1711307567
transform 1 0 980 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1711307567
transform 1 0 892 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1711307567
transform 1 0 1612 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1711307567
transform 1 0 1596 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1711307567
transform 1 0 1492 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1711307567
transform 1 0 1476 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1711307567
transform 1 0 2076 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1711307567
transform 1 0 1676 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1711307567
transform 1 0 1084 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1711307567
transform 1 0 1084 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1711307567
transform 1 0 700 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1711307567
transform 1 0 2668 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1711307567
transform 1 0 2660 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1711307567
transform 1 0 2636 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1711307567
transform 1 0 2580 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1711307567
transform 1 0 2628 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1711307567
transform 1 0 2604 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1711307567
transform 1 0 2572 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1711307567
transform 1 0 2740 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1711307567
transform 1 0 2652 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1711307567
transform 1 0 2564 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1711307567
transform 1 0 2556 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1711307567
transform 1 0 2524 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1711307567
transform 1 0 196 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1711307567
transform 1 0 116 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1711307567
transform 1 0 1068 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1711307567
transform 1 0 1028 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1711307567
transform 1 0 972 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1711307567
transform 1 0 2708 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1711307567
transform 1 0 2644 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1711307567
transform 1 0 2644 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1711307567
transform 1 0 2604 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1711307567
transform 1 0 2524 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1711307567
transform 1 0 2468 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1711307567
transform 1 0 2316 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1711307567
transform 1 0 2284 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1711307567
transform 1 0 2324 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1711307567
transform 1 0 2292 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1711307567
transform 1 0 2316 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1711307567
transform 1 0 2284 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1711307567
transform 1 0 2580 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1711307567
transform 1 0 2428 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1711307567
transform 1 0 2548 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1711307567
transform 1 0 2428 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1711307567
transform 1 0 2468 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1711307567
transform 1 0 2436 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1711307567
transform 1 0 2540 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1711307567
transform 1 0 2516 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1711307567
transform 1 0 2516 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1711307567
transform 1 0 2468 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1711307567
transform 1 0 2580 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1711307567
transform 1 0 2532 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1711307567
transform 1 0 1620 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1711307567
transform 1 0 1268 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1711307567
transform 1 0 1580 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1711307567
transform 1 0 1508 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1711307567
transform 1 0 1204 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1711307567
transform 1 0 1780 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1711307567
transform 1 0 1716 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1711307567
transform 1 0 1980 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1711307567
transform 1 0 1964 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1711307567
transform 1 0 1900 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1711307567
transform 1 0 2012 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1711307567
transform 1 0 1884 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1711307567
transform 1 0 1860 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1711307567
transform 1 0 1828 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1711307567
transform 1 0 1852 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1711307567
transform 1 0 1716 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1711307567
transform 1 0 1716 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1711307567
transform 1 0 1660 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1711307567
transform 1 0 1652 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1711307567
transform 1 0 1540 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1711307567
transform 1 0 1484 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1711307567
transform 1 0 332 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1711307567
transform 1 0 308 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1711307567
transform 1 0 228 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1711307567
transform 1 0 220 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1711307567
transform 1 0 364 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1711307567
transform 1 0 220 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1711307567
transform 1 0 836 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1711307567
transform 1 0 676 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1711307567
transform 1 0 364 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1711307567
transform 1 0 308 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1711307567
transform 1 0 268 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1711307567
transform 1 0 484 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1711307567
transform 1 0 372 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1711307567
transform 1 0 332 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1711307567
transform 1 0 292 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1711307567
transform 1 0 420 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1711307567
transform 1 0 380 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1711307567
transform 1 0 364 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1711307567
transform 1 0 668 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1711307567
transform 1 0 572 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1711307567
transform 1 0 548 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1711307567
transform 1 0 604 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1711307567
transform 1 0 524 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1711307567
transform 1 0 508 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1711307567
transform 1 0 364 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1711307567
transform 1 0 684 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1711307567
transform 1 0 516 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1711307567
transform 1 0 1372 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1711307567
transform 1 0 796 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1711307567
transform 1 0 796 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1711307567
transform 1 0 772 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1711307567
transform 1 0 660 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1711307567
transform 1 0 1300 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1711307567
transform 1 0 828 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1711307567
transform 1 0 860 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1711307567
transform 1 0 732 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1711307567
transform 1 0 652 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1711307567
transform 1 0 572 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1711307567
transform 1 0 516 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1711307567
transform 1 0 724 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1711307567
transform 1 0 676 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1711307567
transform 1 0 636 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1711307567
transform 1 0 1628 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1711307567
transform 1 0 1388 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1711307567
transform 1 0 1028 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1711307567
transform 1 0 1004 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1711307567
transform 1 0 836 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1711307567
transform 1 0 508 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1711307567
transform 1 0 468 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1711307567
transform 1 0 396 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1711307567
transform 1 0 2180 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1711307567
transform 1 0 2140 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1711307567
transform 1 0 1412 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1711307567
transform 1 0 1116 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1711307567
transform 1 0 1492 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1711307567
transform 1 0 1004 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1711307567
transform 1 0 1004 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1711307567
transform 1 0 852 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1711307567
transform 1 0 852 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1711307567
transform 1 0 804 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1711307567
transform 1 0 1348 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1711307567
transform 1 0 1092 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1711307567
transform 1 0 1276 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1711307567
transform 1 0 1140 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1711307567
transform 1 0 1236 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1711307567
transform 1 0 1148 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1711307567
transform 1 0 988 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1711307567
transform 1 0 868 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1711307567
transform 1 0 1212 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1711307567
transform 1 0 1140 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1711307567
transform 1 0 1076 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1711307567
transform 1 0 996 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1711307567
transform 1 0 1100 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1711307567
transform 1 0 980 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1711307567
transform 1 0 980 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1711307567
transform 1 0 876 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1711307567
transform 1 0 804 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1711307567
transform 1 0 764 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1711307567
transform 1 0 1124 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1711307567
transform 1 0 1084 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1711307567
transform 1 0 956 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1711307567
transform 1 0 828 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1711307567
transform 1 0 1492 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1711307567
transform 1 0 1364 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1711307567
transform 1 0 1540 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1711307567
transform 1 0 1316 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1711307567
transform 1 0 1244 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1711307567
transform 1 0 1212 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1711307567
transform 1 0 1148 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1711307567
transform 1 0 1860 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1711307567
transform 1 0 1812 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1711307567
transform 1 0 1460 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1711307567
transform 1 0 1436 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1711307567
transform 1 0 1452 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1711307567
transform 1 0 1340 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1711307567
transform 1 0 1532 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1711307567
transform 1 0 1516 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1711307567
transform 1 0 1492 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1711307567
transform 1 0 1492 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1711307567
transform 1 0 1452 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1711307567
transform 1 0 1836 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1711307567
transform 1 0 1756 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1711307567
transform 1 0 1612 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1711307567
transform 1 0 1532 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1711307567
transform 1 0 2196 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1711307567
transform 1 0 2164 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1711307567
transform 1 0 2124 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1711307567
transform 1 0 1580 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1711307567
transform 1 0 1516 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1711307567
transform 1 0 1412 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1711307567
transform 1 0 1412 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1711307567
transform 1 0 1324 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1711307567
transform 1 0 2500 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1711307567
transform 1 0 2452 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1711307567
transform 1 0 1908 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1711307567
transform 1 0 1740 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1711307567
transform 1 0 1548 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1711307567
transform 1 0 1548 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1711307567
transform 1 0 1372 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1711307567
transform 1 0 1324 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1711307567
transform 1 0 2604 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1711307567
transform 1 0 2580 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1711307567
transform 1 0 1916 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1711307567
transform 1 0 1548 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1711307567
transform 1 0 2740 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1711307567
transform 1 0 2668 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1711307567
transform 1 0 2732 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1711307567
transform 1 0 2644 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1711307567
transform 1 0 2580 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1711307567
transform 1 0 2692 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1711307567
transform 1 0 2612 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1711307567
transform 1 0 2732 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1711307567
transform 1 0 2692 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1711307567
transform 1 0 2636 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1711307567
transform 1 0 2540 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1711307567
transform 1 0 2620 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1711307567
transform 1 0 2548 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1711307567
transform 1 0 2692 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1711307567
transform 1 0 2564 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1711307567
transform 1 0 2516 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1711307567
transform 1 0 2572 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1711307567
transform 1 0 2548 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1711307567
transform 1 0 2548 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1711307567
transform 1 0 2500 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1711307567
transform 1 0 2212 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1711307567
transform 1 0 2140 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1711307567
transform 1 0 2756 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1711307567
transform 1 0 2684 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1711307567
transform 1 0 2756 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1711307567
transform 1 0 2724 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1711307567
transform 1 0 2732 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1711307567
transform 1 0 2676 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1711307567
transform 1 0 2676 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1711307567
transform 1 0 2156 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1711307567
transform 1 0 2116 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1711307567
transform 1 0 2036 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1711307567
transform 1 0 2028 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1711307567
transform 1 0 2012 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1711307567
transform 1 0 1956 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1711307567
transform 1 0 1636 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1711307567
transform 1 0 1540 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1711307567
transform 1 0 1540 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1711307567
transform 1 0 1540 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1711307567
transform 1 0 1540 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1711307567
transform 1 0 1476 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1711307567
transform 1 0 1372 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1711307567
transform 1 0 1292 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1711307567
transform 1 0 1268 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1711307567
transform 1 0 1156 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1711307567
transform 1 0 2676 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1711307567
transform 1 0 932 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1711307567
transform 1 0 780 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1711307567
transform 1 0 636 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1711307567
transform 1 0 516 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1711307567
transform 1 0 388 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1711307567
transform 1 0 356 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1711307567
transform 1 0 348 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1711307567
transform 1 0 268 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1711307567
transform 1 0 148 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1711307567
transform 1 0 84 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1711307567
transform 1 0 2668 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1711307567
transform 1 0 2660 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1711307567
transform 1 0 2572 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1711307567
transform 1 0 2484 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1711307567
transform 1 0 2460 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1711307567
transform 1 0 2452 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1711307567
transform 1 0 2404 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1711307567
transform 1 0 2372 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1711307567
transform 1 0 2356 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1711307567
transform 1 0 2308 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1711307567
transform 1 0 2244 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1711307567
transform 1 0 2244 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1711307567
transform 1 0 2212 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1711307567
transform 1 0 2676 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1711307567
transform 1 0 2676 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1711307567
transform 1 0 2676 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1711307567
transform 1 0 2620 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1711307567
transform 1 0 2620 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1711307567
transform 1 0 2556 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1711307567
transform 1 0 2508 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1711307567
transform 1 0 2460 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1711307567
transform 1 0 2460 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1711307567
transform 1 0 2364 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1711307567
transform 1 0 2324 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1711307567
transform 1 0 2324 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1711307567
transform 1 0 2268 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1711307567
transform 1 0 2204 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1711307567
transform 1 0 2124 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1711307567
transform 1 0 2124 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1711307567
transform 1 0 2068 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1711307567
transform 1 0 1900 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1711307567
transform 1 0 1820 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1711307567
transform 1 0 1788 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1711307567
transform 1 0 1780 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1711307567
transform 1 0 1772 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1711307567
transform 1 0 1748 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1711307567
transform 1 0 1652 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1711307567
transform 1 0 1564 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1711307567
transform 1 0 1396 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1711307567
transform 1 0 1340 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1711307567
transform 1 0 1340 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1711307567
transform 1 0 1316 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1711307567
transform 1 0 1196 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1711307567
transform 1 0 1060 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1711307567
transform 1 0 860 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1711307567
transform 1 0 1484 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1711307567
transform 1 0 1436 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1711307567
transform 1 0 1356 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1711307567
transform 1 0 1356 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1711307567
transform 1 0 948 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1711307567
transform 1 0 684 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1711307567
transform 1 0 636 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1711307567
transform 1 0 564 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1711307567
transform 1 0 564 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1711307567
transform 1 0 516 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1711307567
transform 1 0 444 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1711307567
transform 1 0 244 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1711307567
transform 1 0 236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1711307567
transform 1 0 148 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1711307567
transform 1 0 140 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1711307567
transform 1 0 84 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1711307567
transform 1 0 84 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1711307567
transform 1 0 2444 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1711307567
transform 1 0 2348 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1711307567
transform 1 0 2252 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1711307567
transform 1 0 2196 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1711307567
transform 1 0 2108 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1711307567
transform 1 0 2084 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1711307567
transform 1 0 2020 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1711307567
transform 1 0 2020 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1711307567
transform 1 0 1988 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1711307567
transform 1 0 1820 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1711307567
transform 1 0 1716 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1711307567
transform 1 0 1708 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1711307567
transform 1 0 1612 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1711307567
transform 1 0 1572 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1711307567
transform 1 0 1508 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1711307567
transform 1 0 1428 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1711307567
transform 1 0 1356 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1711307567
transform 1 0 1316 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1711307567
transform 1 0 1228 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1711307567
transform 1 0 1156 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1711307567
transform 1 0 1156 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1711307567
transform 1 0 1060 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1711307567
transform 1 0 1020 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1711307567
transform 1 0 940 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1711307567
transform 1 0 852 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1711307567
transform 1 0 764 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1711307567
transform 1 0 676 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1711307567
transform 1 0 620 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1711307567
transform 1 0 596 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1711307567
transform 1 0 484 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1711307567
transform 1 0 380 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1711307567
transform 1 0 2556 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1711307567
transform 1 0 2476 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1711307567
transform 1 0 2476 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1711307567
transform 1 0 2428 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1711307567
transform 1 0 2412 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1711307567
transform 1 0 2372 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1711307567
transform 1 0 2324 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1711307567
transform 1 0 2292 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1711307567
transform 1 0 2204 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1711307567
transform 1 0 1476 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1711307567
transform 1 0 1476 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1711307567
transform 1 0 308 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1711307567
transform 1 0 308 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1711307567
transform 1 0 220 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1711307567
transform 1 0 132 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1711307567
transform 1 0 2028 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1711307567
transform 1 0 1532 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1711307567
transform 1 0 1516 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1711307567
transform 1 0 1460 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1711307567
transform 1 0 1524 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1711307567
transform 1 0 1492 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1711307567
transform 1 0 1420 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1711307567
transform 1 0 2548 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1711307567
transform 1 0 2452 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1711307567
transform 1 0 2396 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1711307567
transform 1 0 2380 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1711307567
transform 1 0 2372 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1711307567
transform 1 0 2356 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1711307567
transform 1 0 2340 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1711307567
transform 1 0 2300 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1711307567
transform 1 0 2300 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1711307567
transform 1 0 2284 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1711307567
transform 1 0 2284 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1711307567
transform 1 0 2228 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1711307567
transform 1 0 2228 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1711307567
transform 1 0 2180 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1711307567
transform 1 0 2180 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1711307567
transform 1 0 2140 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1711307567
transform 1 0 2092 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1711307567
transform 1 0 2092 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1711307567
transform 1 0 2012 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1711307567
transform 1 0 1772 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1711307567
transform 1 0 1772 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1711307567
transform 1 0 1660 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1711307567
transform 1 0 1660 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1711307567
transform 1 0 1444 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1711307567
transform 1 0 1188 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1711307567
transform 1 0 1180 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1711307567
transform 1 0 196 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1711307567
transform 1 0 188 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1711307567
transform 1 0 164 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1711307567
transform 1 0 2652 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1711307567
transform 1 0 2636 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1711307567
transform 1 0 2596 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1711307567
transform 1 0 2580 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1711307567
transform 1 0 2372 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1711307567
transform 1 0 2364 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1711307567
transform 1 0 2356 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1711307567
transform 1 0 2292 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1711307567
transform 1 0 2252 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1711307567
transform 1 0 2196 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1711307567
transform 1 0 2172 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1711307567
transform 1 0 2060 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1711307567
transform 1 0 2004 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1711307567
transform 1 0 2116 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1711307567
transform 1 0 2052 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1711307567
transform 1 0 1940 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1711307567
transform 1 0 1852 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1711307567
transform 1 0 1716 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1711307567
transform 1 0 1564 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1711307567
transform 1 0 1412 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1711307567
transform 1 0 1332 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1711307567
transform 1 0 1172 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1711307567
transform 1 0 1084 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1711307567
transform 1 0 1068 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1711307567
transform 1 0 1052 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1711307567
transform 1 0 2364 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1711307567
transform 1 0 772 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1711307567
transform 1 0 692 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1711307567
transform 1 0 604 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1711307567
transform 1 0 500 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1711307567
transform 1 0 396 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1711307567
transform 1 0 388 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1711307567
transform 1 0 388 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1711307567
transform 1 0 308 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1711307567
transform 1 0 172 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1711307567
transform 1 0 124 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1711307567
transform 1 0 1940 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1711307567
transform 1 0 1740 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1711307567
transform 1 0 1732 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1711307567
transform 1 0 1652 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1711307567
transform 1 0 1548 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1711307567
transform 1 0 1548 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1711307567
transform 1 0 1532 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1711307567
transform 1 0 1228 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1711307567
transform 1 0 1204 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1711307567
transform 1 0 1204 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1711307567
transform 1 0 1180 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1711307567
transform 1 0 1044 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1711307567
transform 1 0 924 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1711307567
transform 1 0 844 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1711307567
transform 1 0 644 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1711307567
transform 1 0 644 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1711307567
transform 1 0 468 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1711307567
transform 1 0 468 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1711307567
transform 1 0 428 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1711307567
transform 1 0 428 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1711307567
transform 1 0 396 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1711307567
transform 1 0 2300 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1711307567
transform 1 0 2284 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1711307567
transform 1 0 2236 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1711307567
transform 1 0 2236 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1711307567
transform 1 0 1892 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1711307567
transform 1 0 1884 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1711307567
transform 1 0 1612 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1711307567
transform 1 0 1356 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1711307567
transform 1 0 1164 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1711307567
transform 1 0 980 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1711307567
transform 1 0 804 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1711307567
transform 1 0 804 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1711307567
transform 1 0 708 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1711307567
transform 1 0 708 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1711307567
transform 1 0 636 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1711307567
transform 1 0 340 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1711307567
transform 1 0 2620 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1711307567
transform 1 0 2300 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1711307567
transform 1 0 2268 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1711307567
transform 1 0 2260 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1711307567
transform 1 0 2212 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1711307567
transform 1 0 2132 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1711307567
transform 1 0 2132 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1711307567
transform 1 0 2116 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1711307567
transform 1 0 2116 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1711307567
transform 1 0 2076 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1711307567
transform 1 0 2044 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1711307567
transform 1 0 2044 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1711307567
transform 1 0 2044 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1711307567
transform 1 0 1852 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1711307567
transform 1 0 1852 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1711307567
transform 1 0 1812 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1711307567
transform 1 0 1812 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1711307567
transform 1 0 1788 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1711307567
transform 1 0 1380 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1711307567
transform 1 0 1380 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1711307567
transform 1 0 1356 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1711307567
transform 1 0 1300 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1711307567
transform 1 0 1140 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1711307567
transform 1 0 1124 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1711307567
transform 1 0 1036 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1711307567
transform 1 0 916 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1711307567
transform 1 0 756 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1711307567
transform 1 0 668 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1711307567
transform 1 0 660 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1711307567
transform 1 0 652 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1711307567
transform 1 0 468 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1711307567
transform 1 0 452 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1711307567
transform 1 0 444 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1711307567
transform 1 0 388 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1711307567
transform 1 0 220 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1711307567
transform 1 0 220 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1711307567
transform 1 0 196 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1711307567
transform 1 0 196 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1711307567
transform 1 0 1932 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1711307567
transform 1 0 1876 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1711307567
transform 1 0 1828 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1711307567
transform 1 0 1828 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1711307567
transform 1 0 1660 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1711307567
transform 1 0 2044 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1711307567
transform 1 0 1924 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1711307567
transform 1 0 1852 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1711307567
transform 1 0 1772 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1711307567
transform 1 0 1676 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1711307567
transform 1 0 1580 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1711307567
transform 1 0 1572 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1711307567
transform 1 0 1420 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1711307567
transform 1 0 1380 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1711307567
transform 1 0 1212 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1711307567
transform 1 0 1204 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1711307567
transform 1 0 1140 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1711307567
transform 1 0 2308 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1711307567
transform 1 0 2012 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1711307567
transform 1 0 1988 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1711307567
transform 1 0 1012 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1711307567
transform 1 0 940 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1711307567
transform 1 0 860 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1711307567
transform 1 0 636 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1711307567
transform 1 0 2204 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1711307567
transform 1 0 1964 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1711307567
transform 1 0 420 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1711307567
transform 1 0 420 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1711307567
transform 1 0 420 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1711307567
transform 1 0 340 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1711307567
transform 1 0 324 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1711307567
transform 1 0 300 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1711307567
transform 1 0 220 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1711307567
transform 1 0 196 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1711307567
transform 1 0 140 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1711307567
transform 1 0 1940 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1711307567
transform 1 0 1844 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1711307567
transform 1 0 244 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1711307567
transform 1 0 2492 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1711307567
transform 1 0 2364 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1711307567
transform 1 0 2348 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1711307567
transform 1 0 2116 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1711307567
transform 1 0 2036 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1711307567
transform 1 0 1804 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1711307567
transform 1 0 1716 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1711307567
transform 1 0 2212 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1711307567
transform 1 0 2164 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1711307567
transform 1 0 2108 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1711307567
transform 1 0 1956 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1711307567
transform 1 0 1812 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1711307567
transform 1 0 1812 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1711307567
transform 1 0 1628 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1711307567
transform 1 0 1628 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1711307567
transform 1 0 1452 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1711307567
transform 1 0 1396 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1711307567
transform 1 0 1276 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1711307567
transform 1 0 1260 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1711307567
transform 1 0 684 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1711307567
transform 1 0 676 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1711307567
transform 1 0 612 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1711307567
transform 1 0 484 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1711307567
transform 1 0 484 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1711307567
transform 1 0 404 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1711307567
transform 1 0 404 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1711307567
transform 1 0 332 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1711307567
transform 1 0 316 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1711307567
transform 1 0 316 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1711307567
transform 1 0 292 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1711307567
transform 1 0 236 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1711307567
transform 1 0 236 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1711307567
transform 1 0 188 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1711307567
transform 1 0 2172 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1711307567
transform 1 0 2164 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1711307567
transform 1 0 2132 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1711307567
transform 1 0 2124 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1711307567
transform 1 0 2124 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1711307567
transform 1 0 2108 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1711307567
transform 1 0 2108 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1711307567
transform 1 0 2076 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1711307567
transform 1 0 2004 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1711307567
transform 1 0 1996 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1711307567
transform 1 0 1820 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1711307567
transform 1 0 1812 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1711307567
transform 1 0 1748 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1711307567
transform 1 0 1740 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1711307567
transform 1 0 1708 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1711307567
transform 1 0 1500 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1711307567
transform 1 0 1420 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1711307567
transform 1 0 1388 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1711307567
transform 1 0 1372 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1711307567
transform 1 0 1316 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1711307567
transform 1 0 1316 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1711307567
transform 1 0 1276 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1711307567
transform 1 0 1068 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1711307567
transform 1 0 1052 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1711307567
transform 1 0 1004 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1711307567
transform 1 0 996 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1711307567
transform 1 0 996 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1711307567
transform 1 0 996 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1711307567
transform 1 0 852 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1711307567
transform 1 0 764 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1711307567
transform 1 0 716 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1711307567
transform 1 0 684 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1711307567
transform 1 0 676 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1711307567
transform 1 0 588 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1711307567
transform 1 0 492 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1711307567
transform 1 0 492 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1711307567
transform 1 0 316 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1711307567
transform 1 0 268 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1711307567
transform 1 0 2060 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1711307567
transform 1 0 2028 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1711307567
transform 1 0 1996 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1711307567
transform 1 0 1924 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1711307567
transform 1 0 1916 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1711307567
transform 1 0 1836 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1711307567
transform 1 0 1636 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1711307567
transform 1 0 1564 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1711307567
transform 1 0 1020 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1711307567
transform 1 0 924 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1711307567
transform 1 0 476 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1711307567
transform 1 0 2012 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1711307567
transform 1 0 1996 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1711307567
transform 1 0 1972 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1711307567
transform 1 0 1940 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1711307567
transform 1 0 1932 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1711307567
transform 1 0 1884 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1711307567
transform 1 0 1812 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1711307567
transform 1 0 1804 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1711307567
transform 1 0 1732 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1711307567
transform 1 0 1596 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1711307567
transform 1 0 1548 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1711307567
transform 1 0 996 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1711307567
transform 1 0 900 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1711307567
transform 1 0 876 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1711307567
transform 1 0 444 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1711307567
transform 1 0 444 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1711307567
transform 1 0 388 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1711307567
transform 1 0 388 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1711307567
transform 1 0 300 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1711307567
transform 1 0 2444 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1711307567
transform 1 0 2228 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1711307567
transform 1 0 1988 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1711307567
transform 1 0 388 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1711307567
transform 1 0 1988 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1711307567
transform 1 0 1644 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1711307567
transform 1 0 1588 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1711307567
transform 1 0 1524 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1711307567
transform 1 0 1524 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1711307567
transform 1 0 1428 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1711307567
transform 1 0 1324 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1711307567
transform 1 0 1300 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1711307567
transform 1 0 1172 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1711307567
transform 1 0 1172 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1711307567
transform 1 0 1036 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1711307567
transform 1 0 924 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1711307567
transform 1 0 916 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1711307567
transform 1 0 780 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1711307567
transform 1 0 676 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1711307567
transform 1 0 564 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1711307567
transform 1 0 476 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1711307567
transform 1 0 372 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1711307567
transform 1 0 2292 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1711307567
transform 1 0 2220 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1711307567
transform 1 0 1596 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1711307567
transform 1 0 1436 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1711307567
transform 1 0 1276 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1711307567
transform 1 0 1244 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1711307567
transform 1 0 1116 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1711307567
transform 1 0 940 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1711307567
transform 1 0 836 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1711307567
transform 1 0 708 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1711307567
transform 1 0 636 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1711307567
transform 1 0 588 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1711307567
transform 1 0 2572 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1711307567
transform 1 0 2444 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1711307567
transform 1 0 2276 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1711307567
transform 1 0 2212 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1711307567
transform 1 0 2092 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1711307567
transform 1 0 2092 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1711307567
transform 1 0 1716 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1711307567
transform 1 0 1716 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1711307567
transform 1 0 1452 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1711307567
transform 1 0 1452 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1711307567
transform 1 0 444 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1711307567
transform 1 0 412 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1711307567
transform 1 0 412 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1711307567
transform 1 0 308 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1711307567
transform 1 0 212 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1711307567
transform 1 0 2620 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1711307567
transform 1 0 2548 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1711307567
transform 1 0 2540 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1711307567
transform 1 0 2492 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1711307567
transform 1 0 2308 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1711307567
transform 1 0 2212 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1711307567
transform 1 0 1996 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1711307567
transform 1 0 1964 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1711307567
transform 1 0 1948 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1711307567
transform 1 0 1924 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1711307567
transform 1 0 1876 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1711307567
transform 1 0 1876 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1711307567
transform 1 0 2124 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1711307567
transform 1 0 2068 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1711307567
transform 1 0 2060 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1711307567
transform 1 0 1980 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1711307567
transform 1 0 1908 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1711307567
transform 1 0 1836 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1711307567
transform 1 0 1836 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1711307567
transform 1 0 1820 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1711307567
transform 1 0 1820 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1711307567
transform 1 0 1300 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1711307567
transform 1 0 1300 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1711307567
transform 1 0 1228 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1711307567
transform 1 0 1228 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1711307567
transform 1 0 1012 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1711307567
transform 1 0 1012 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1711307567
transform 1 0 964 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1711307567
transform 1 0 748 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1711307567
transform 1 0 740 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1711307567
transform 1 0 732 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1711307567
transform 1 0 676 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1711307567
transform 1 0 676 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1711307567
transform 1 0 2284 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1711307567
transform 1 0 2260 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1711307567
transform 1 0 2260 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1711307567
transform 1 0 2148 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1711307567
transform 1 0 1900 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1711307567
transform 1 0 1572 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1711307567
transform 1 0 1452 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1711307567
transform 1 0 1452 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1711307567
transform 1 0 452 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1711307567
transform 1 0 388 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1711307567
transform 1 0 1020 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1711307567
transform 1 0 1004 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1711307567
transform 1 0 1572 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1711307567
transform 1 0 1540 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1711307567
transform 1 0 1028 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1711307567
transform 1 0 996 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1711307567
transform 1 0 1868 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1711307567
transform 1 0 1612 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1711307567
transform 1 0 1788 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1711307567
transform 1 0 348 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1711307567
transform 1 0 2188 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1711307567
transform 1 0 2116 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1711307567
transform 1 0 1780 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1711307567
transform 1 0 1708 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1711307567
transform 1 0 876 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1711307567
transform 1 0 724 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1711307567
transform 1 0 540 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1711307567
transform 1 0 788 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1711307567
transform 1 0 788 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1711307567
transform 1 0 748 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1711307567
transform 1 0 628 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1711307567
transform 1 0 540 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1711307567
transform 1 0 548 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1711307567
transform 1 0 364 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1711307567
transform 1 0 300 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1711307567
transform 1 0 692 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1711307567
transform 1 0 452 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1711307567
transform 1 0 1572 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1711307567
transform 1 0 1452 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1711307567
transform 1 0 1452 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1711307567
transform 1 0 772 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1711307567
transform 1 0 588 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1711307567
transform 1 0 1500 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1711307567
transform 1 0 1428 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1711307567
transform 1 0 804 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1711307567
transform 1 0 804 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1711307567
transform 1 0 580 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1711307567
transform 1 0 1900 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1711307567
transform 1 0 1796 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1711307567
transform 1 0 1172 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1711307567
transform 1 0 1156 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1711307567
transform 1 0 716 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1711307567
transform 1 0 388 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1711307567
transform 1 0 772 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1711307567
transform 1 0 716 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1711307567
transform 1 0 652 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1711307567
transform 1 0 604 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1711307567
transform 1 0 596 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1711307567
transform 1 0 1508 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1711307567
transform 1 0 1284 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1711307567
transform 1 0 1276 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1711307567
transform 1 0 1140 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1711307567
transform 1 0 1428 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1711307567
transform 1 0 1364 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1711307567
transform 1 0 1364 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1711307567
transform 1 0 1324 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1711307567
transform 1 0 1292 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1711307567
transform 1 0 1292 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1711307567
transform 1 0 1228 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1711307567
transform 1 0 2324 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1711307567
transform 1 0 2276 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1711307567
transform 1 0 2276 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1711307567
transform 1 0 1612 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1711307567
transform 1 0 1548 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1711307567
transform 1 0 1548 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1711307567
transform 1 0 1508 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1711307567
transform 1 0 1436 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1711307567
transform 1 0 1420 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1711307567
transform 1 0 1348 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1711307567
transform 1 0 1164 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1711307567
transform 1 0 1156 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1711307567
transform 1 0 884 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1711307567
transform 1 0 884 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1711307567
transform 1 0 884 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1711307567
transform 1 0 828 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1711307567
transform 1 0 828 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1711307567
transform 1 0 764 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1711307567
transform 1 0 484 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1711307567
transform 1 0 484 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1711307567
transform 1 0 476 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1711307567
transform 1 0 476 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1711307567
transform 1 0 428 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1711307567
transform 1 0 380 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1711307567
transform 1 0 340 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1711307567
transform 1 0 340 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1711307567
transform 1 0 340 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1711307567
transform 1 0 324 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1711307567
transform 1 0 292 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1711307567
transform 1 0 1356 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1711307567
transform 1 0 1076 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1711307567
transform 1 0 2220 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1711307567
transform 1 0 2180 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1711307567
transform 1 0 2108 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1711307567
transform 1 0 500 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1711307567
transform 1 0 420 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1711307567
transform 1 0 420 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1711307567
transform 1 0 356 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1711307567
transform 1 0 2276 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1711307567
transform 1 0 2220 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1711307567
transform 1 0 2204 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1711307567
transform 1 0 2164 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1711307567
transform 1 0 1980 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1711307567
transform 1 0 1756 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1711307567
transform 1 0 1380 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1711307567
transform 1 0 764 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1711307567
transform 1 0 548 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1711307567
transform 1 0 1940 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1711307567
transform 1 0 1844 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1711307567
transform 1 0 1236 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1711307567
transform 1 0 1228 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1711307567
transform 1 0 732 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1711307567
transform 1 0 420 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1711307567
transform 1 0 2284 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1711307567
transform 1 0 2260 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1711307567
transform 1 0 2052 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1711307567
transform 1 0 2036 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1711307567
transform 1 0 2036 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1711307567
transform 1 0 1684 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1711307567
transform 1 0 1564 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1711307567
transform 1 0 1516 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1711307567
transform 1 0 1444 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1711307567
transform 1 0 1380 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1711307567
transform 1 0 948 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1711307567
transform 1 0 948 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1711307567
transform 1 0 948 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1711307567
transform 1 0 948 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1711307567
transform 1 0 540 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1711307567
transform 1 0 500 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1711307567
transform 1 0 492 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1711307567
transform 1 0 348 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1711307567
transform 1 0 2556 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1711307567
transform 1 0 2052 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1711307567
transform 1 0 2044 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1711307567
transform 1 0 2020 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1711307567
transform 1 0 2020 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1711307567
transform 1 0 2004 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1711307567
transform 1 0 1180 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1711307567
transform 1 0 1164 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1711307567
transform 1 0 1164 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1711307567
transform 1 0 884 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1711307567
transform 1 0 804 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1711307567
transform 1 0 804 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1711307567
transform 1 0 788 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1711307567
transform 1 0 764 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1711307567
transform 1 0 764 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1711307567
transform 1 0 700 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1711307567
transform 1 0 692 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1711307567
transform 1 0 620 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1711307567
transform 1 0 620 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1711307567
transform 1 0 540 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1711307567
transform 1 0 540 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1711307567
transform 1 0 244 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1711307567
transform 1 0 2740 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1711307567
transform 1 0 2652 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1711307567
transform 1 0 2732 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1711307567
transform 1 0 2668 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1711307567
transform 1 0 2580 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1711307567
transform 1 0 2532 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1711307567
transform 1 0 2596 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1711307567
transform 1 0 2292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1711307567
transform 1 0 2580 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1711307567
transform 1 0 2508 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1711307567
transform 1 0 2524 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1711307567
transform 1 0 2412 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1711307567
transform 1 0 2516 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1711307567
transform 1 0 2452 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1711307567
transform 1 0 2564 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1711307567
transform 1 0 2468 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1711307567
transform 1 0 2020 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1711307567
transform 1 0 1996 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1711307567
transform 1 0 1876 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1711307567
transform 1 0 2444 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1711307567
transform 1 0 2404 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1711307567
transform 1 0 2220 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1711307567
transform 1 0 1964 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1711307567
transform 1 0 2468 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1711307567
transform 1 0 2236 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1711307567
transform 1 0 2356 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1711307567
transform 1 0 2204 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1711307567
transform 1 0 1740 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1711307567
transform 1 0 1740 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1711307567
transform 1 0 1700 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1711307567
transform 1 0 1700 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1711307567
transform 1 0 1748 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1711307567
transform 1 0 1540 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1711307567
transform 1 0 1524 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1711307567
transform 1 0 1508 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1711307567
transform 1 0 1084 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1711307567
transform 1 0 908 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1711307567
transform 1 0 1092 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1711307567
transform 1 0 1044 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1711307567
transform 1 0 516 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1711307567
transform 1 0 484 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1711307567
transform 1 0 436 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1711307567
transform 1 0 180 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1711307567
transform 1 0 388 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1711307567
transform 1 0 356 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1711307567
transform 1 0 316 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1711307567
transform 1 0 268 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1711307567
transform 1 0 1428 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1711307567
transform 1 0 1420 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1711307567
transform 1 0 1356 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1711307567
transform 1 0 1356 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1711307567
transform 1 0 1420 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1711307567
transform 1 0 1380 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1711307567
transform 1 0 1724 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1711307567
transform 1 0 1452 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1711307567
transform 1 0 1628 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1711307567
transform 1 0 1452 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1711307567
transform 1 0 1468 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1711307567
transform 1 0 1068 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1711307567
transform 1 0 1028 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1711307567
transform 1 0 572 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1711307567
transform 1 0 1228 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1711307567
transform 1 0 1124 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1711307567
transform 1 0 1724 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1711307567
transform 1 0 1668 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1711307567
transform 1 0 1604 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1711307567
transform 1 0 1628 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1711307567
transform 1 0 1124 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1711307567
transform 1 0 1124 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1711307567
transform 1 0 932 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1711307567
transform 1 0 932 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1711307567
transform 1 0 692 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1711307567
transform 1 0 612 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1711307567
transform 1 0 516 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1711307567
transform 1 0 572 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1711307567
transform 1 0 492 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1711307567
transform 1 0 460 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1711307567
transform 1 0 292 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1711307567
transform 1 0 540 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1711307567
transform 1 0 420 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1711307567
transform 1 0 412 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1711307567
transform 1 0 332 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1711307567
transform 1 0 332 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1711307567
transform 1 0 292 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1711307567
transform 1 0 572 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1711307567
transform 1 0 532 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1711307567
transform 1 0 476 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1711307567
transform 1 0 1508 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1711307567
transform 1 0 1084 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1711307567
transform 1 0 1084 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1711307567
transform 1 0 468 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1711307567
transform 1 0 476 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1711307567
transform 1 0 436 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1711307567
transform 1 0 428 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1711307567
transform 1 0 396 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1711307567
transform 1 0 1476 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1711307567
transform 1 0 1372 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1711307567
transform 1 0 1372 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1711307567
transform 1 0 1140 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1711307567
transform 1 0 548 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1711307567
transform 1 0 412 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1711307567
transform 1 0 316 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1711307567
transform 1 0 260 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1711307567
transform 1 0 1804 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1711307567
transform 1 0 1708 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1711307567
transform 1 0 1772 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1711307567
transform 1 0 1740 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1711307567
transform 1 0 2196 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1711307567
transform 1 0 2164 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1711307567
transform 1 0 2164 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1711307567
transform 1 0 1748 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1711307567
transform 1 0 1740 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1711307567
transform 1 0 1636 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1711307567
transform 1 0 1524 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1711307567
transform 1 0 1492 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1711307567
transform 1 0 1476 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1711307567
transform 1 0 1764 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1711307567
transform 1 0 1748 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1711307567
transform 1 0 2132 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1711307567
transform 1 0 1772 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1711307567
transform 1 0 1652 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1711307567
transform 1 0 1844 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1711307567
transform 1 0 1796 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1711307567
transform 1 0 1940 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1711307567
transform 1 0 1860 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1711307567
transform 1 0 2084 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1711307567
transform 1 0 1948 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1711307567
transform 1 0 2132 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1711307567
transform 1 0 1964 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1711307567
transform 1 0 1308 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1711307567
transform 1 0 1028 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1711307567
transform 1 0 1412 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1711307567
transform 1 0 1332 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1711307567
transform 1 0 1484 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1711307567
transform 1 0 1388 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1711307567
transform 1 0 1700 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1711307567
transform 1 0 1628 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1711307567
transform 1 0 1580 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1711307567
transform 1 0 1412 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1711307567
transform 1 0 1372 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1711307567
transform 1 0 1404 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1711307567
transform 1 0 1284 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1711307567
transform 1 0 1668 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1711307567
transform 1 0 1556 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1711307567
transform 1 0 1436 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1711307567
transform 1 0 1348 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1711307567
transform 1 0 1284 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1711307567
transform 1 0 1572 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1711307567
transform 1 0 1484 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1711307567
transform 1 0 1260 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1711307567
transform 1 0 1148 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1711307567
transform 1 0 1412 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1711307567
transform 1 0 1364 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1711307567
transform 1 0 1196 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1711307567
transform 1 0 996 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1711307567
transform 1 0 980 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1711307567
transform 1 0 980 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1711307567
transform 1 0 852 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1711307567
transform 1 0 812 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1711307567
transform 1 0 980 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1711307567
transform 1 0 812 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1711307567
transform 1 0 932 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1711307567
transform 1 0 724 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1711307567
transform 1 0 1052 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1711307567
transform 1 0 972 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1711307567
transform 1 0 1060 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1711307567
transform 1 0 1036 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1711307567
transform 1 0 1004 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1711307567
transform 1 0 1004 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1711307567
transform 1 0 724 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1711307567
transform 1 0 668 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1711307567
transform 1 0 1260 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1711307567
transform 1 0 1156 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1711307567
transform 1 0 1356 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1711307567
transform 1 0 860 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1711307567
transform 1 0 1388 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1711307567
transform 1 0 1316 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1711307567
transform 1 0 1356 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1711307567
transform 1 0 1268 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1711307567
transform 1 0 1364 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1711307567
transform 1 0 1188 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1711307567
transform 1 0 1132 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1711307567
transform 1 0 1668 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1711307567
transform 1 0 1596 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1711307567
transform 1 0 1532 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1711307567
transform 1 0 1380 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1711307567
transform 1 0 1380 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1711307567
transform 1 0 1340 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1711307567
transform 1 0 1332 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1711307567
transform 1 0 1588 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1711307567
transform 1 0 1548 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1711307567
transform 1 0 1396 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1711307567
transform 1 0 1468 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1711307567
transform 1 0 1228 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1711307567
transform 1 0 1188 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1711307567
transform 1 0 1172 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1711307567
transform 1 0 1172 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1711307567
transform 1 0 1172 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1711307567
transform 1 0 636 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1711307567
transform 1 0 572 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1711307567
transform 1 0 1164 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1711307567
transform 1 0 1052 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1711307567
transform 1 0 1676 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1711307567
transform 1 0 1604 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1711307567
transform 1 0 1444 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1711307567
transform 1 0 1284 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1711307567
transform 1 0 1308 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1711307567
transform 1 0 1148 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1711307567
transform 1 0 1148 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1711307567
transform 1 0 940 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1711307567
transform 1 0 1460 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1711307567
transform 1 0 1428 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1711307567
transform 1 0 1540 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1711307567
transform 1 0 1452 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1711307567
transform 1 0 2004 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1711307567
transform 1 0 1804 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1711307567
transform 1 0 1796 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1711307567
transform 1 0 1732 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1711307567
transform 1 0 1516 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1711307567
transform 1 0 1540 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1711307567
transform 1 0 572 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1711307567
transform 1 0 1132 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1711307567
transform 1 0 1092 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1711307567
transform 1 0 828 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1711307567
transform 1 0 820 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1711307567
transform 1 0 620 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1711307567
transform 1 0 556 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1711307567
transform 1 0 564 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1711307567
transform 1 0 524 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1711307567
transform 1 0 460 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1711307567
transform 1 0 460 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1711307567
transform 1 0 428 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1711307567
transform 1 0 1396 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1711307567
transform 1 0 1276 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1711307567
transform 1 0 1268 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1711307567
transform 1 0 1204 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1711307567
transform 1 0 1204 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1711307567
transform 1 0 1436 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1711307567
transform 1 0 1412 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1711307567
transform 1 0 1516 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1711307567
transform 1 0 1372 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1711307567
transform 1 0 1372 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1711307567
transform 1 0 1300 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1711307567
transform 1 0 1300 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1711307567
transform 1 0 1044 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1711307567
transform 1 0 1044 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1711307567
transform 1 0 1012 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1711307567
transform 1 0 1996 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1711307567
transform 1 0 1988 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1711307567
transform 1 0 1948 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1711307567
transform 1 0 1908 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1711307567
transform 1 0 1668 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1711307567
transform 1 0 1428 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1711307567
transform 1 0 1692 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1711307567
transform 1 0 1660 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1711307567
transform 1 0 1420 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1711307567
transform 1 0 804 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1711307567
transform 1 0 708 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1711307567
transform 1 0 932 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1711307567
transform 1 0 868 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1711307567
transform 1 0 980 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1711307567
transform 1 0 948 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1711307567
transform 1 0 940 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1711307567
transform 1 0 796 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1711307567
transform 1 0 644 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1711307567
transform 1 0 1044 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1711307567
transform 1 0 1020 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1711307567
transform 1 0 1436 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1711307567
transform 1 0 1332 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1711307567
transform 1 0 1244 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1711307567
transform 1 0 1020 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1711307567
transform 1 0 1044 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1711307567
transform 1 0 948 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1711307567
transform 1 0 948 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1711307567
transform 1 0 932 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1711307567
transform 1 0 1604 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1711307567
transform 1 0 868 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1711307567
transform 1 0 892 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1711307567
transform 1 0 844 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1711307567
transform 1 0 788 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1711307567
transform 1 0 372 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1711307567
transform 1 0 1988 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1711307567
transform 1 0 1940 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1711307567
transform 1 0 1820 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1711307567
transform 1 0 1732 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1711307567
transform 1 0 1732 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1711307567
transform 1 0 1652 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1711307567
transform 1 0 508 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1711307567
transform 1 0 508 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1711307567
transform 1 0 396 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1711307567
transform 1 0 340 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1711307567
transform 1 0 1828 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1711307567
transform 1 0 1596 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1711307567
transform 1 0 1620 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1711307567
transform 1 0 1620 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1711307567
transform 1 0 1612 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1711307567
transform 1 0 1604 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1711307567
transform 1 0 1556 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1711307567
transform 1 0 1524 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1711307567
transform 1 0 2028 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1711307567
transform 1 0 1812 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1711307567
transform 1 0 1804 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1711307567
transform 1 0 1708 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1711307567
transform 1 0 1556 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1711307567
transform 1 0 1868 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1711307567
transform 1 0 1852 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1711307567
transform 1 0 716 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1711307567
transform 1 0 604 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1711307567
transform 1 0 460 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1711307567
transform 1 0 764 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1711307567
transform 1 0 732 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1711307567
transform 1 0 732 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1711307567
transform 1 0 692 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1711307567
transform 1 0 1260 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1711307567
transform 1 0 772 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1711307567
transform 1 0 556 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1711307567
transform 1 0 412 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1711307567
transform 1 0 260 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1711307567
transform 1 0 260 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1711307567
transform 1 0 228 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1711307567
transform 1 0 228 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1711307567
transform 1 0 180 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1711307567
transform 1 0 804 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1711307567
transform 1 0 596 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1711307567
transform 1 0 484 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1711307567
transform 1 0 844 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1711307567
transform 1 0 668 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1711307567
transform 1 0 1292 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1711307567
transform 1 0 1052 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1711307567
transform 1 0 1284 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1711307567
transform 1 0 876 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1711307567
transform 1 0 940 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1711307567
transform 1 0 844 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1711307567
transform 1 0 860 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1711307567
transform 1 0 708 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1711307567
transform 1 0 628 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1711307567
transform 1 0 580 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1711307567
transform 1 0 676 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1711307567
transform 1 0 500 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1711307567
transform 1 0 332 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1711307567
transform 1 0 1220 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1711307567
transform 1 0 716 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1711307567
transform 1 0 508 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1711307567
transform 1 0 340 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1711307567
transform 1 0 300 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1711307567
transform 1 0 884 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1711307567
transform 1 0 580 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1711307567
transform 1 0 1644 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1711307567
transform 1 0 1420 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1711307567
transform 1 0 844 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1711307567
transform 1 0 1004 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1711307567
transform 1 0 908 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1711307567
transform 1 0 868 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1711307567
transform 1 0 964 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1711307567
transform 1 0 900 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1711307567
transform 1 0 884 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1711307567
transform 1 0 708 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1711307567
transform 1 0 660 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1711307567
transform 1 0 1564 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1711307567
transform 1 0 900 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1711307567
transform 1 0 908 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1711307567
transform 1 0 844 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1711307567
transform 1 0 1220 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1711307567
transform 1 0 948 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1711307567
transform 1 0 1332 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1711307567
transform 1 0 1212 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1711307567
transform 1 0 1252 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1711307567
transform 1 0 996 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1711307567
transform 1 0 996 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1711307567
transform 1 0 972 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1711307567
transform 1 0 956 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1711307567
transform 1 0 900 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1711307567
transform 1 0 772 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1711307567
transform 1 0 652 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1711307567
transform 1 0 604 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1711307567
transform 1 0 748 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1711307567
transform 1 0 460 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1711307567
transform 1 0 412 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1711307567
transform 1 0 396 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1711307567
transform 1 0 412 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1711307567
transform 1 0 292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1711307567
transform 1 0 276 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1711307567
transform 1 0 1828 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1711307567
transform 1 0 1556 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1711307567
transform 1 0 1572 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1711307567
transform 1 0 1532 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1711307567
transform 1 0 2068 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1711307567
transform 1 0 1884 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1711307567
transform 1 0 1836 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1711307567
transform 1 0 1836 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1711307567
transform 1 0 1772 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1711307567
transform 1 0 1996 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1711307567
transform 1 0 1916 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1711307567
transform 1 0 2068 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1711307567
transform 1 0 1948 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1711307567
transform 1 0 1340 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1711307567
transform 1 0 1276 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1711307567
transform 1 0 1276 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1711307567
transform 1 0 1244 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1711307567
transform 1 0 1468 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1711307567
transform 1 0 1348 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1711307567
transform 1 0 1228 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1711307567
transform 1 0 692 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1711307567
transform 1 0 692 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1711307567
transform 1 0 460 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1711307567
transform 1 0 436 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1711307567
transform 1 0 1340 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1711307567
transform 1 0 1316 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1711307567
transform 1 0 1508 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1711307567
transform 1 0 1372 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1711307567
transform 1 0 1788 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1711307567
transform 1 0 1628 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1711307567
transform 1 0 1628 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1711307567
transform 1 0 1468 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1711307567
transform 1 0 1492 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1711307567
transform 1 0 1380 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1711307567
transform 1 0 1380 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1711307567
transform 1 0 588 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1711307567
transform 1 0 580 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1711307567
transform 1 0 444 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1711307567
transform 1 0 1276 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1711307567
transform 1 0 1172 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1711307567
transform 1 0 1340 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1711307567
transform 1 0 1316 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1711307567
transform 1 0 1660 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1711307567
transform 1 0 1572 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1711307567
transform 1 0 1380 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1711307567
transform 1 0 788 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1711307567
transform 1 0 708 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1711307567
transform 1 0 708 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1711307567
transform 1 0 652 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1711307567
transform 1 0 1564 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1711307567
transform 1 0 1548 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1711307567
transform 1 0 1524 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1711307567
transform 1 0 1524 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1711307567
transform 1 0 1460 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1711307567
transform 1 0 1436 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1711307567
transform 1 0 1436 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1711307567
transform 1 0 1396 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1711307567
transform 1 0 1380 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1711307567
transform 1 0 1308 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1711307567
transform 1 0 2036 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1711307567
transform 1 0 1708 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1711307567
transform 1 0 1876 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1711307567
transform 1 0 1756 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1711307567
transform 1 0 1756 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1711307567
transform 1 0 1652 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1711307567
transform 1 0 1948 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1711307567
transform 1 0 1780 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1711307567
transform 1 0 1588 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1711307567
transform 1 0 1588 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1711307567
transform 1 0 1524 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1711307567
transform 1 0 1444 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1711307567
transform 1 0 1724 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1711307567
transform 1 0 1636 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1711307567
transform 1 0 2052 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1711307567
transform 1 0 1732 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1711307567
transform 1 0 212 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1711307567
transform 1 0 140 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1711307567
transform 1 0 276 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1711307567
transform 1 0 180 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1711307567
transform 1 0 260 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1711307567
transform 1 0 188 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1711307567
transform 1 0 532 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1711307567
transform 1 0 308 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1711307567
transform 1 0 268 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1711307567
transform 1 0 300 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1711307567
transform 1 0 212 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1711307567
transform 1 0 1948 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1711307567
transform 1 0 212 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1711307567
transform 1 0 188 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1711307567
transform 1 0 188 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1711307567
transform 1 0 188 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1711307567
transform 1 0 132 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1711307567
transform 1 0 244 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1711307567
transform 1 0 164 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1711307567
transform 1 0 228 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1711307567
transform 1 0 172 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1711307567
transform 1 0 252 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1711307567
transform 1 0 220 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1711307567
transform 1 0 548 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1711307567
transform 1 0 276 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1711307567
transform 1 0 172 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1711307567
transform 1 0 124 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1711307567
transform 1 0 180 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1711307567
transform 1 0 148 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1711307567
transform 1 0 212 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1711307567
transform 1 0 164 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1711307567
transform 1 0 308 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1711307567
transform 1 0 228 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1711307567
transform 1 0 188 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1711307567
transform 1 0 1108 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1711307567
transform 1 0 668 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1711307567
transform 1 0 668 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1711307567
transform 1 0 420 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1711307567
transform 1 0 316 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1711307567
transform 1 0 308 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1711307567
transform 1 0 276 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1711307567
transform 1 0 252 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1711307567
transform 1 0 548 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1711307567
transform 1 0 388 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1711307567
transform 1 0 276 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1711307567
transform 1 0 236 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1711307567
transform 1 0 236 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1711307567
transform 1 0 2420 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1711307567
transform 1 0 1788 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1711307567
transform 1 0 1948 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1711307567
transform 1 0 1740 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1711307567
transform 1 0 636 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1711307567
transform 1 0 380 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1711307567
transform 1 0 324 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1711307567
transform 1 0 332 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1711307567
transform 1 0 308 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1711307567
transform 1 0 2348 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1711307567
transform 1 0 1996 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1711307567
transform 1 0 1620 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1711307567
transform 1 0 972 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1711307567
transform 1 0 668 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1711307567
transform 1 0 500 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1711307567
transform 1 0 356 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1711307567
transform 1 0 2364 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1711307567
transform 1 0 1940 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1711307567
transform 1 0 660 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1711307567
transform 1 0 524 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1711307567
transform 1 0 1988 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1711307567
transform 1 0 1988 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1711307567
transform 1 0 1900 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1711307567
transform 1 0 1540 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1711307567
transform 1 0 1044 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1711307567
transform 1 0 660 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1711307567
transform 1 0 484 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1711307567
transform 1 0 396 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1711307567
transform 1 0 420 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1711307567
transform 1 0 420 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1711307567
transform 1 0 540 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1711307567
transform 1 0 476 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1711307567
transform 1 0 2084 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1711307567
transform 1 0 1988 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1711307567
transform 1 0 1572 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1711307567
transform 1 0 1124 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1711307567
transform 1 0 668 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1711307567
transform 1 0 700 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1711307567
transform 1 0 604 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1711307567
transform 1 0 876 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1711307567
transform 1 0 572 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1711307567
transform 1 0 572 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1711307567
transform 1 0 556 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1711307567
transform 1 0 540 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1711307567
transform 1 0 516 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1711307567
transform 1 0 484 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1711307567
transform 1 0 404 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1711307567
transform 1 0 2132 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1711307567
transform 1 0 2132 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1711307567
transform 1 0 2060 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1711307567
transform 1 0 1684 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1711307567
transform 1 0 1676 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1711307567
transform 1 0 1612 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1711307567
transform 1 0 1612 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1711307567
transform 1 0 1196 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1711307567
transform 1 0 1196 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1711307567
transform 1 0 1124 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1711307567
transform 1 0 644 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1711307567
transform 1 0 612 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1711307567
transform 1 0 532 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1711307567
transform 1 0 508 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1711307567
transform 1 0 500 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1711307567
transform 1 0 444 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1711307567
transform 1 0 580 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1711307567
transform 1 0 500 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1711307567
transform 1 0 764 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1711307567
transform 1 0 708 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1711307567
transform 1 0 500 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1711307567
transform 1 0 1844 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1711307567
transform 1 0 1676 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1711307567
transform 1 0 1668 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1711307567
transform 1 0 1580 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1711307567
transform 1 0 1484 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1711307567
transform 1 0 1460 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1711307567
transform 1 0 1460 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1711307567
transform 1 0 1164 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1711307567
transform 1 0 788 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1711307567
transform 1 0 756 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1711307567
transform 1 0 708 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1711307567
transform 1 0 612 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1711307567
transform 1 0 812 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1711307567
transform 1 0 732 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1711307567
transform 1 0 868 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1711307567
transform 1 0 732 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1711307567
transform 1 0 644 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1711307567
transform 1 0 700 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1711307567
transform 1 0 668 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1711307567
transform 1 0 788 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1711307567
transform 1 0 748 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1711307567
transform 1 0 900 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1711307567
transform 1 0 796 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1711307567
transform 1 0 796 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1711307567
transform 1 0 604 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1711307567
transform 1 0 708 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1711307567
transform 1 0 612 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1711307567
transform 1 0 652 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1711307567
transform 1 0 604 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1711307567
transform 1 0 1012 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1711307567
transform 1 0 932 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1711307567
transform 1 0 876 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1711307567
transform 1 0 860 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1711307567
transform 1 0 828 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1711307567
transform 1 0 1076 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1711307567
transform 1 0 1052 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1711307567
transform 1 0 1052 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1711307567
transform 1 0 892 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1711307567
transform 1 0 1996 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1711307567
transform 1 0 1124 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1711307567
transform 1 0 1116 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1711307567
transform 1 0 1060 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1711307567
transform 1 0 972 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1711307567
transform 1 0 1076 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1711307567
transform 1 0 1028 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1711307567
transform 1 0 1116 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1711307567
transform 1 0 1028 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1711307567
transform 1 0 1156 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1711307567
transform 1 0 1092 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1711307567
transform 1 0 1052 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1711307567
transform 1 0 988 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1711307567
transform 1 0 1140 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1711307567
transform 1 0 1100 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1711307567
transform 1 0 1180 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1711307567
transform 1 0 1108 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1711307567
transform 1 0 1196 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1711307567
transform 1 0 1148 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1711307567
transform 1 0 1228 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1711307567
transform 1 0 1164 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1711307567
transform 1 0 1068 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1711307567
transform 1 0 1148 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1711307567
transform 1 0 1012 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1711307567
transform 1 0 1492 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1711307567
transform 1 0 1212 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1711307567
transform 1 0 1212 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1711307567
transform 1 0 1164 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1711307567
transform 1 0 1172 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1711307567
transform 1 0 1124 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1711307567
transform 1 0 1276 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1711307567
transform 1 0 1236 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1711307567
transform 1 0 1204 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1711307567
transform 1 0 1172 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1711307567
transform 1 0 1140 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1711307567
transform 1 0 1004 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1711307567
transform 1 0 1204 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1711307567
transform 1 0 1188 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1711307567
transform 1 0 1188 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1711307567
transform 1 0 1116 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1711307567
transform 1 0 988 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1711307567
transform 1 0 1084 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1711307567
transform 1 0 940 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1711307567
transform 1 0 1020 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1711307567
transform 1 0 988 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1711307567
transform 1 0 1452 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1711307567
transform 1 0 1220 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1711307567
transform 1 0 1340 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1711307567
transform 1 0 1284 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1711307567
transform 1 0 1156 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1711307567
transform 1 0 1292 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1711307567
transform 1 0 1236 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1711307567
transform 1 0 1132 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1711307567
transform 1 0 1564 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1711307567
transform 1 0 1540 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1711307567
transform 1 0 1668 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1711307567
transform 1 0 1588 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1711307567
transform 1 0 1980 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1711307567
transform 1 0 1716 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1711307567
transform 1 0 1692 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1711307567
transform 1 0 1604 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1711307567
transform 1 0 1580 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1711307567
transform 1 0 1580 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1711307567
transform 1 0 1580 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1711307567
transform 1 0 1556 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1711307567
transform 1 0 1556 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1711307567
transform 1 0 2292 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1711307567
transform 1 0 2108 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1711307567
transform 1 0 2108 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1711307567
transform 1 0 2084 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1711307567
transform 1 0 1884 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1711307567
transform 1 0 1540 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1711307567
transform 1 0 1540 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1711307567
transform 1 0 1508 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1711307567
transform 1 0 1572 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1711307567
transform 1 0 1516 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1711307567
transform 1 0 1516 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1711307567
transform 1 0 1444 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1711307567
transform 1 0 2324 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1711307567
transform 1 0 2180 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1711307567
transform 1 0 1708 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1711307567
transform 1 0 1548 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1711307567
transform 1 0 1748 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1711307567
transform 1 0 1700 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1711307567
transform 1 0 1772 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1711307567
transform 1 0 1652 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1711307567
transform 1 0 2244 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1711307567
transform 1 0 2212 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1711307567
transform 1 0 2212 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1711307567
transform 1 0 2092 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1711307567
transform 1 0 1628 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1711307567
transform 1 0 1588 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1711307567
transform 1 0 1900 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1711307567
transform 1 0 1724 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1711307567
transform 1 0 1716 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1711307567
transform 1 0 1628 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1711307567
transform 1 0 1836 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1711307567
transform 1 0 1772 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1711307567
transform 1 0 1716 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1711307567
transform 1 0 2396 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1711307567
transform 1 0 2284 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1711307567
transform 1 0 1884 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1711307567
transform 1 0 1796 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1711307567
transform 1 0 1924 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1711307567
transform 1 0 1684 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1711307567
transform 1 0 1876 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1711307567
transform 1 0 1852 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1711307567
transform 1 0 2188 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1711307567
transform 1 0 2124 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1711307567
transform 1 0 2068 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1711307567
transform 1 0 1988 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1711307567
transform 1 0 2116 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1711307567
transform 1 0 1972 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1711307567
transform 1 0 1964 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1711307567
transform 1 0 1940 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1711307567
transform 1 0 2220 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1711307567
transform 1 0 2180 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1711307567
transform 1 0 1980 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1711307567
transform 1 0 1916 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1711307567
transform 1 0 2116 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1711307567
transform 1 0 2020 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1711307567
transform 1 0 1972 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1711307567
transform 1 0 2124 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1711307567
transform 1 0 2052 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1711307567
transform 1 0 2172 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1711307567
transform 1 0 2076 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1711307567
transform 1 0 2020 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1711307567
transform 1 0 1988 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1711307567
transform 1 0 1972 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1711307567
transform 1 0 1916 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1711307567
transform 1 0 1852 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1711307567
transform 1 0 1940 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1711307567
transform 1 0 1940 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1711307567
transform 1 0 1908 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1711307567
transform 1 0 1868 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1711307567
transform 1 0 1852 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1711307567
transform 1 0 1788 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1711307567
transform 1 0 1820 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1711307567
transform 1 0 1764 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1711307567
transform 1 0 1996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1711307567
transform 1 0 1900 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1711307567
transform 1 0 2196 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1711307567
transform 1 0 1980 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1711307567
transform 1 0 1852 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1711307567
transform 1 0 2012 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1711307567
transform 1 0 1972 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1711307567
transform 1 0 2036 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1711307567
transform 1 0 1964 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1711307567
transform 1 0 2060 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1711307567
transform 1 0 2028 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1711307567
transform 1 0 2228 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1711307567
transform 1 0 2204 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1711307567
transform 1 0 2148 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1711307567
transform 1 0 2148 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1711307567
transform 1 0 2148 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1711307567
transform 1 0 2140 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1711307567
transform 1 0 2084 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1711307567
transform 1 0 2084 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1711307567
transform 1 0 2028 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1711307567
transform 1 0 1972 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1711307567
transform 1 0 2212 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1711307567
transform 1 0 2084 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1711307567
transform 1 0 1844 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1711307567
transform 1 0 1620 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1711307567
transform 1 0 1556 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1711307567
transform 1 0 2236 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1711307567
transform 1 0 2140 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1711307567
transform 1 0 1908 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1711307567
transform 1 0 2300 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1711307567
transform 1 0 2276 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1711307567
transform 1 0 2228 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1711307567
transform 1 0 2156 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1711307567
transform 1 0 2308 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1711307567
transform 1 0 2268 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1711307567
transform 1 0 2220 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1711307567
transform 1 0 2180 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1711307567
transform 1 0 1884 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1711307567
transform 1 0 1580 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1711307567
transform 1 0 1524 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1711307567
transform 1 0 2076 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1711307567
transform 1 0 1980 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1711307567
transform 1 0 2196 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1711307567
transform 1 0 2148 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1711307567
transform 1 0 2084 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1711307567
transform 1 0 2108 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1711307567
transform 1 0 2060 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1711307567
transform 1 0 2108 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1711307567
transform 1 0 2076 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1711307567
transform 1 0 2716 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1711307567
transform 1 0 2684 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1711307567
transform 1 0 2660 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1711307567
transform 1 0 2628 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1711307567
transform 1 0 2556 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1711307567
transform 1 0 2540 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1711307567
transform 1 0 2532 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1711307567
transform 1 0 2724 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1711307567
transform 1 0 2708 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1711307567
transform 1 0 2676 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1711307567
transform 1 0 2676 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1711307567
transform 1 0 2572 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1711307567
transform 1 0 2588 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1711307567
transform 1 0 2524 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1711307567
transform 1 0 2740 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1711307567
transform 1 0 2708 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1711307567
transform 1 0 2676 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1711307567
transform 1 0 2676 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1711307567
transform 1 0 2660 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1711307567
transform 1 0 2644 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1711307567
transform 1 0 2636 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1711307567
transform 1 0 2604 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1711307567
transform 1 0 2732 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1711307567
transform 1 0 2724 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1711307567
transform 1 0 2724 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1711307567
transform 1 0 2676 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1711307567
transform 1 0 2676 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1711307567
transform 1 0 2668 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1711307567
transform 1 0 2660 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1711307567
transform 1 0 2604 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1711307567
transform 1 0 2580 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1711307567
transform 1 0 2668 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1711307567
transform 1 0 2540 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1711307567
transform 1 0 2708 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1711307567
transform 1 0 2596 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1711307567
transform 1 0 2652 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1711307567
transform 1 0 2604 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1711307567
transform 1 0 2588 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1711307567
transform 1 0 2540 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1711307567
transform 1 0 2708 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1711307567
transform 1 0 2572 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1711307567
transform 1 0 2724 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1711307567
transform 1 0 2612 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1711307567
transform 1 0 2412 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1711307567
transform 1 0 2308 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1711307567
transform 1 0 2212 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1711307567
transform 1 0 2148 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1711307567
transform 1 0 2044 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1711307567
transform 1 0 1948 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1711307567
transform 1 0 1980 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1711307567
transform 1 0 1812 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1711307567
transform 1 0 1868 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1711307567
transform 1 0 1844 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1711307567
transform 1 0 1804 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1711307567
transform 1 0 1740 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1711307567
transform 1 0 1676 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1711307567
transform 1 0 1596 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1711307567
transform 1 0 1028 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1711307567
transform 1 0 908 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1711307567
transform 1 0 1044 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1711307567
transform 1 0 972 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1711307567
transform 1 0 772 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1711307567
transform 1 0 684 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1711307567
transform 1 0 180 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1711307567
transform 1 0 132 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1711307567
transform 1 0 2308 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1711307567
transform 1 0 2252 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1711307567
transform 1 0 2244 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1711307567
transform 1 0 2188 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1711307567
transform 1 0 2156 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1711307567
transform 1 0 2076 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1711307567
transform 1 0 2004 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1711307567
transform 1 0 2308 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1711307567
transform 1 0 2268 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1711307567
transform 1 0 2204 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1711307567
transform 1 0 2164 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1711307567
transform 1 0 2476 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1711307567
transform 1 0 2140 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1711307567
transform 1 0 2172 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1711307567
transform 1 0 2132 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1711307567
transform 1 0 2084 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1711307567
transform 1 0 1956 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1711307567
transform 1 0 1884 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1711307567
transform 1 0 2172 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1711307567
transform 1 0 2132 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1711307567
transform 1 0 2076 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1711307567
transform 1 0 1964 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1711307567
transform 1 0 2132 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1711307567
transform 1 0 2060 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1711307567
transform 1 0 2132 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1711307567
transform 1 0 2052 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1711307567
transform 1 0 2140 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1711307567
transform 1 0 2084 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1711307567
transform 1 0 2132 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1711307567
transform 1 0 2068 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1711307567
transform 1 0 2036 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1711307567
transform 1 0 2020 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1711307567
transform 1 0 1980 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1711307567
transform 1 0 2116 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1711307567
transform 1 0 1948 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1711307567
transform 1 0 2012 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1711307567
transform 1 0 1916 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1711307567
transform 1 0 1908 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1711307567
transform 1 0 1812 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1711307567
transform 1 0 1916 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1711307567
transform 1 0 1844 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1711307567
transform 1 0 1820 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1711307567
transform 1 0 1780 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1711307567
transform 1 0 1692 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1711307567
transform 1 0 1492 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1711307567
transform 1 0 1940 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1711307567
transform 1 0 1820 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1711307567
transform 1 0 1708 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1711307567
transform 1 0 1636 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1711307567
transform 1 0 1972 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1711307567
transform 1 0 1892 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1711307567
transform 1 0 1860 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1711307567
transform 1 0 1788 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1711307567
transform 1 0 1684 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1711307567
transform 1 0 1548 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1711307567
transform 1 0 2420 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1711307567
transform 1 0 2364 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1711307567
transform 1 0 2348 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1711307567
transform 1 0 2348 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1711307567
transform 1 0 2268 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1711307567
transform 1 0 1732 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1711307567
transform 1 0 1580 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1711307567
transform 1 0 1828 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1711307567
transform 1 0 1660 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1711307567
transform 1 0 1756 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1711307567
transform 1 0 1644 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1711307567
transform 1 0 1644 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1711307567
transform 1 0 1500 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1711307567
transform 1 0 1388 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1711307567
transform 1 0 1908 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1711307567
transform 1 0 1652 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1711307567
transform 1 0 1772 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1711307567
transform 1 0 1540 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1711307567
transform 1 0 1836 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1711307567
transform 1 0 1468 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1711307567
transform 1 0 1692 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1711307567
transform 1 0 1564 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1711307567
transform 1 0 1500 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1711307567
transform 1 0 1468 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1711307567
transform 1 0 1468 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1711307567
transform 1 0 1396 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1711307567
transform 1 0 1364 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1711307567
transform 1 0 1316 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1711307567
transform 1 0 1244 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1711307567
transform 1 0 1244 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1711307567
transform 1 0 1188 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1711307567
transform 1 0 1180 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1711307567
transform 1 0 1084 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1711307567
transform 1 0 1428 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1711307567
transform 1 0 1140 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1711307567
transform 1 0 1140 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1711307567
transform 1 0 1092 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1711307567
transform 1 0 1004 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1711307567
transform 1 0 980 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1711307567
transform 1 0 940 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1711307567
transform 1 0 876 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1711307567
transform 1 0 780 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1711307567
transform 1 0 1748 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1711307567
transform 1 0 1612 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1711307567
transform 1 0 1460 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1711307567
transform 1 0 1596 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1711307567
transform 1 0 1572 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1711307567
transform 1 0 1420 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1711307567
transform 1 0 1276 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1711307567
transform 1 0 1188 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1711307567
transform 1 0 1180 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1711307567
transform 1 0 1164 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1711307567
transform 1 0 1300 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1711307567
transform 1 0 1236 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1711307567
transform 1 0 1260 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1711307567
transform 1 0 1156 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1711307567
transform 1 0 1164 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1711307567
transform 1 0 1036 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1711307567
transform 1 0 1204 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1711307567
transform 1 0 1156 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1711307567
transform 1 0 1452 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1711307567
transform 1 0 1340 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1711307567
transform 1 0 1332 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1711307567
transform 1 0 1020 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1711307567
transform 1 0 916 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1711307567
transform 1 0 964 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1711307567
transform 1 0 892 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1711307567
transform 1 0 892 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1711307567
transform 1 0 820 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1711307567
transform 1 0 1372 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1711307567
transform 1 0 1308 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1711307567
transform 1 0 1172 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1711307567
transform 1 0 1124 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1711307567
transform 1 0 1004 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1711307567
transform 1 0 916 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1711307567
transform 1 0 796 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1711307567
transform 1 0 668 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1711307567
transform 1 0 852 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1711307567
transform 1 0 756 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1711307567
transform 1 0 908 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1711307567
transform 1 0 844 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1711307567
transform 1 0 900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1711307567
transform 1 0 692 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1711307567
transform 1 0 940 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1711307567
transform 1 0 612 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1711307567
transform 1 0 1524 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1711307567
transform 1 0 948 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1711307567
transform 1 0 948 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1711307567
transform 1 0 700 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1711307567
transform 1 0 708 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1711307567
transform 1 0 532 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1711307567
transform 1 0 652 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1711307567
transform 1 0 580 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1711307567
transform 1 0 420 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1711307567
transform 1 0 300 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1711307567
transform 1 0 588 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1711307567
transform 1 0 452 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1711307567
transform 1 0 460 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1711307567
transform 1 0 372 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1711307567
transform 1 0 612 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1711307567
transform 1 0 468 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1711307567
transform 1 0 812 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1711307567
transform 1 0 524 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1711307567
transform 1 0 1316 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1711307567
transform 1 0 828 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1711307567
transform 1 0 332 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1711307567
transform 1 0 284 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1711307567
transform 1 0 444 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1711307567
transform 1 0 340 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1711307567
transform 1 0 572 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1711307567
transform 1 0 492 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1711307567
transform 1 0 436 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1711307567
transform 1 0 628 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1711307567
transform 1 0 564 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1711307567
transform 1 0 564 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1711307567
transform 1 0 484 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1711307567
transform 1 0 468 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1711307567
transform 1 0 292 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1711307567
transform 1 0 244 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1711307567
transform 1 0 452 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1711307567
transform 1 0 340 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1711307567
transform 1 0 412 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1711307567
transform 1 0 348 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1711307567
transform 1 0 548 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1711307567
transform 1 0 444 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1711307567
transform 1 0 396 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1711307567
transform 1 0 372 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1711307567
transform 1 0 548 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1711307567
transform 1 0 436 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1711307567
transform 1 0 788 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1711307567
transform 1 0 612 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1711307567
transform 1 0 588 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1711307567
transform 1 0 372 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1711307567
transform 1 0 2660 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1711307567
transform 1 0 2628 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1711307567
transform 1 0 2524 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1711307567
transform 1 0 2476 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1711307567
transform 1 0 2452 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1711307567
transform 1 0 2468 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1711307567
transform 1 0 2436 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1711307567
transform 1 0 2612 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1711307567
transform 1 0 2540 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1711307567
transform 1 0 2548 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1711307567
transform 1 0 2436 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1711307567
transform 1 0 2364 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1711307567
transform 1 0 1532 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1711307567
transform 1 0 2628 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1711307567
transform 1 0 2532 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1711307567
transform 1 0 2540 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1711307567
transform 1 0 2428 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1711307567
transform 1 0 1564 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1711307567
transform 1 0 1340 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1711307567
transform 1 0 2468 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1711307567
transform 1 0 2180 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1711307567
transform 1 0 1940 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1711307567
transform 1 0 308 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1711307567
transform 1 0 276 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1711307567
transform 1 0 1068 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1711307567
transform 1 0 1012 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1711307567
transform 1 0 2340 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1711307567
transform 1 0 2260 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1711307567
transform 1 0 2388 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1711307567
transform 1 0 2308 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1711307567
transform 1 0 2388 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1711307567
transform 1 0 2292 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1711307567
transform 1 0 2524 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1711307567
transform 1 0 2476 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1711307567
transform 1 0 2116 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1711307567
transform 1 0 2004 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1711307567
transform 1 0 1756 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1711307567
transform 1 0 1684 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1711307567
transform 1 0 1556 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1711307567
transform 1 0 1500 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1711307567
transform 1 0 1476 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1711307567
transform 1 0 1412 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1711307567
transform 1 0 1620 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1711307567
transform 1 0 1524 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1711307567
transform 1 0 892 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1711307567
transform 1 0 852 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1711307567
transform 1 0 484 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1711307567
transform 1 0 436 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1711307567
transform 1 0 244 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1711307567
transform 1 0 196 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1711307567
transform 1 0 364 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1711307567
transform 1 0 316 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1711307567
transform 1 0 252 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1711307567
transform 1 0 132 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1711307567
transform 1 0 228 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1711307567
transform 1 0 124 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1711307567
transform 1 0 236 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1711307567
transform 1 0 132 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1711307567
transform 1 0 444 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1711307567
transform 1 0 396 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1711307567
transform 1 0 2700 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1711307567
transform 1 0 2620 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1711307567
transform 1 0 2700 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1711307567
transform 1 0 2628 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1711307567
transform 1 0 2652 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1711307567
transform 1 0 2548 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1711307567
transform 1 0 2492 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1711307567
transform 1 0 2436 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1711307567
transform 1 0 2628 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1711307567
transform 1 0 2556 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1711307567
transform 1 0 2412 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1711307567
transform 1 0 2140 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1711307567
transform 1 0 2540 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1711307567
transform 1 0 2420 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1711307567
transform 1 0 2244 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1711307567
transform 1 0 1732 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1711307567
transform 1 0 1668 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1711307567
transform 1 0 1668 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1711307567
transform 1 0 1292 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1711307567
transform 1 0 2540 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1711307567
transform 1 0 2460 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1711307567
transform 1 0 2412 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1711307567
transform 1 0 2412 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1711307567
transform 1 0 2340 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1711307567
transform 1 0 1964 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1711307567
transform 1 0 1964 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1711307567
transform 1 0 1876 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1711307567
transform 1 0 1732 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1711307567
transform 1 0 1732 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1711307567
transform 1 0 1148 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1711307567
transform 1 0 1068 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1711307567
transform 1 0 996 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1711307567
transform 1 0 884 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1711307567
transform 1 0 1740 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1711307567
transform 1 0 1724 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1711307567
transform 1 0 1692 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1711307567
transform 1 0 1692 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1711307567
transform 1 0 1660 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1711307567
transform 1 0 1332 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1711307567
transform 1 0 2404 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1711307567
transform 1 0 2340 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1711307567
transform 1 0 2404 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1711307567
transform 1 0 2268 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1711307567
transform 1 0 380 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1711307567
transform 1 0 308 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1711307567
transform 1 0 292 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1711307567
transform 1 0 244 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1711307567
transform 1 0 228 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1711307567
transform 1 0 284 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1711307567
transform 1 0 260 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1711307567
transform 1 0 148 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1711307567
transform 1 0 300 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1711307567
transform 1 0 268 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1711307567
transform 1 0 268 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1711307567
transform 1 0 252 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1711307567
transform 1 0 228 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1711307567
transform 1 0 428 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1711307567
transform 1 0 324 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1711307567
transform 1 0 476 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1711307567
transform 1 0 356 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1711307567
transform 1 0 212 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1711307567
transform 1 0 508 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1711307567
transform 1 0 460 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1711307567
transform 1 0 396 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1711307567
transform 1 0 548 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1711307567
transform 1 0 500 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1711307567
transform 1 0 476 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1711307567
transform 1 0 476 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1711307567
transform 1 0 604 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1711307567
transform 1 0 548 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1711307567
transform 1 0 988 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1711307567
transform 1 0 900 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1711307567
transform 1 0 2636 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1711307567
transform 1 0 2316 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1711307567
transform 1 0 2316 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1711307567
transform 1 0 2220 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1711307567
transform 1 0 1060 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1711307567
transform 1 0 956 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1711307567
transform 1 0 924 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1711307567
transform 1 0 1172 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1711307567
transform 1 0 1148 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1711307567
transform 1 0 1548 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1711307567
transform 1 0 1444 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1711307567
transform 1 0 1444 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1711307567
transform 1 0 1076 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1711307567
transform 1 0 1076 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1711307567
transform 1 0 884 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1711307567
transform 1 0 1380 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1711307567
transform 1 0 1260 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1711307567
transform 1 0 1100 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1711307567
transform 1 0 1100 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1711307567
transform 1 0 828 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1711307567
transform 1 0 1484 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1711307567
transform 1 0 1388 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1711307567
transform 1 0 1204 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1711307567
transform 1 0 1204 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1711307567
transform 1 0 740 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1711307567
transform 1 0 1620 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1711307567
transform 1 0 1500 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1711307567
transform 1 0 1260 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1711307567
transform 1 0 1252 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1711307567
transform 1 0 1180 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1711307567
transform 1 0 1012 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1711307567
transform 1 0 1676 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1711307567
transform 1 0 1644 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1711307567
transform 1 0 1644 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1711307567
transform 1 0 1612 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1711307567
transform 1 0 1180 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1711307567
transform 1 0 1780 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1711307567
transform 1 0 1780 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1711307567
transform 1 0 1764 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1711307567
transform 1 0 1684 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1711307567
transform 1 0 1660 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1711307567
transform 1 0 1644 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1711307567
transform 1 0 1628 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1711307567
transform 1 0 1220 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1711307567
transform 1 0 2412 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1711307567
transform 1 0 1516 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1711307567
transform 1 0 2212 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1711307567
transform 1 0 2172 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1711307567
transform 1 0 2164 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1711307567
transform 1 0 2140 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1711307567
transform 1 0 2124 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1711307567
transform 1 0 2308 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1711307567
transform 1 0 2276 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1711307567
transform 1 0 2276 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1711307567
transform 1 0 2260 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1711307567
transform 1 0 2100 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1711307567
transform 1 0 2556 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1711307567
transform 1 0 2308 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1711307567
transform 1 0 2260 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1711307567
transform 1 0 2236 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2584
timestamp 1711307567
transform 1 0 2204 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1711307567
transform 1 0 2172 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1711307567
transform 1 0 2188 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1711307567
transform 1 0 2020 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1711307567
transform 1 0 2244 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1711307567
transform 1 0 2156 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1711307567
transform 1 0 2132 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1711307567
transform 1 0 1980 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1711307567
transform 1 0 1892 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1711307567
transform 1 0 2484 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1711307567
transform 1 0 2476 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1711307567
transform 1 0 2452 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1711307567
transform 1 0 2108 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1711307567
transform 1 0 2100 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1711307567
transform 1 0 1892 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2599
timestamp 1711307567
transform 1 0 1852 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1711307567
transform 1 0 1756 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1711307567
transform 1 0 2460 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1711307567
transform 1 0 2340 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1711307567
transform 1 0 2188 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1711307567
transform 1 0 1964 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1711307567
transform 1 0 1964 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1711307567
transform 1 0 1940 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1711307567
transform 1 0 1932 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1711307567
transform 1 0 1924 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1711307567
transform 1 0 1820 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1711307567
transform 1 0 2060 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1711307567
transform 1 0 1932 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1711307567
transform 1 0 1916 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1711307567
transform 1 0 1780 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1711307567
transform 1 0 1676 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1711307567
transform 1 0 1924 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1711307567
transform 1 0 1732 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1711307567
transform 1 0 1940 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1711307567
transform 1 0 1844 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1711307567
transform 1 0 1836 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1711307567
transform 1 0 1828 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1711307567
transform 1 0 1828 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1711307567
transform 1 0 1804 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1711307567
transform 1 0 1804 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1711307567
transform 1 0 1772 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1711307567
transform 1 0 1772 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1711307567
transform 1 0 1732 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1711307567
transform 1 0 1708 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1711307567
transform 1 0 1708 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1711307567
transform 1 0 1876 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1711307567
transform 1 0 1708 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1711307567
transform 1 0 1348 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1711307567
transform 1 0 1284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1711307567
transform 1 0 1260 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1711307567
transform 1 0 1196 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1711307567
transform 1 0 1196 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1711307567
transform 1 0 1140 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1711307567
transform 1 0 1212 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1711307567
transform 1 0 1148 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1711307567
transform 1 0 1284 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1711307567
transform 1 0 1284 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1711307567
transform 1 0 1252 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1711307567
transform 1 0 1044 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1711307567
transform 1 0 900 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1711307567
transform 1 0 700 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1711307567
transform 1 0 1220 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1711307567
transform 1 0 1180 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1711307567
transform 1 0 1116 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1711307567
transform 1 0 1100 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1711307567
transform 1 0 1076 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1711307567
transform 1 0 1060 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1711307567
transform 1 0 1052 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1711307567
transform 1 0 1052 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1711307567
transform 1 0 756 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1711307567
transform 1 0 668 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1711307567
transform 1 0 1116 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1711307567
transform 1 0 940 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1711307567
transform 1 0 828 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1711307567
transform 1 0 572 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1711307567
transform 1 0 1156 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1711307567
transform 1 0 932 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1711307567
transform 1 0 804 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1711307567
transform 1 0 620 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1711307567
transform 1 0 924 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1711307567
transform 1 0 732 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1711307567
transform 1 0 732 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1711307567
transform 1 0 444 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1711307567
transform 1 0 780 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1711307567
transform 1 0 780 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1711307567
transform 1 0 780 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1711307567
transform 1 0 724 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1711307567
transform 1 0 724 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1711307567
transform 1 0 684 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1711307567
transform 1 0 684 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1711307567
transform 1 0 532 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1711307567
transform 1 0 452 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1711307567
transform 1 0 868 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1711307567
transform 1 0 812 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1711307567
transform 1 0 596 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1711307567
transform 1 0 596 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1711307567
transform 1 0 852 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1711307567
transform 1 0 804 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1711307567
transform 1 0 724 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1711307567
transform 1 0 700 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1711307567
transform 1 0 628 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1711307567
transform 1 0 620 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1711307567
transform 1 0 540 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1711307567
transform 1 0 484 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1711307567
transform 1 0 468 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1711307567
transform 1 0 468 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1711307567
transform 1 0 436 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1711307567
transform 1 0 412 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1711307567
transform 1 0 412 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1711307567
transform 1 0 380 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1711307567
transform 1 0 372 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1711307567
transform 1 0 556 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1711307567
transform 1 0 500 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1711307567
transform 1 0 540 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1711307567
transform 1 0 524 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1711307567
transform 1 0 476 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1711307567
transform 1 0 468 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1711307567
transform 1 0 2692 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1711307567
transform 1 0 2676 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1711307567
transform 1 0 2604 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1711307567
transform 1 0 2500 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1711307567
transform 1 0 2356 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1711307567
transform 1 0 2356 0 1 585
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1711307567
transform 1 0 1400 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1711307567
transform 1 0 2216 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1711307567
transform 1 0 2120 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1711307567
transform 1 0 2040 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1711307567
transform 1 0 2128 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1711307567
transform 1 0 1544 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1711307567
transform 1 0 504 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1711307567
transform 1 0 328 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1711307567
transform 1 0 280 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1711307567
transform 1 0 296 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1711307567
transform 1 0 336 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1711307567
transform 1 0 2240 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1711307567
transform 1 0 2160 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1711307567
transform 1 0 1960 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1711307567
transform 1 0 1448 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1711307567
transform 1 0 432 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1711307567
transform 1 0 2600 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1711307567
transform 1 0 2248 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1711307567
transform 1 0 480 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1711307567
transform 1 0 1408 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1711307567
transform 1 0 832 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1711307567
transform 1 0 864 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1711307567
transform 1 0 648 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1711307567
transform 1 0 256 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1711307567
transform 1 0 216 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1711307567
transform 1 0 448 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1711307567
transform 1 0 576 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1711307567
transform 1 0 520 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1711307567
transform 1 0 456 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1711307567
transform 1 0 544 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1711307567
transform 1 0 800 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1711307567
transform 1 0 656 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1711307567
transform 1 0 720 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1711307567
transform 1 0 712 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1711307567
transform 1 0 528 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1711307567
transform 1 0 512 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1711307567
transform 1 0 600 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1711307567
transform 1 0 544 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1711307567
transform 1 0 912 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1711307567
transform 1 0 824 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1711307567
transform 1 0 1952 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1711307567
transform 1 0 768 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1711307567
transform 1 0 776 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1711307567
transform 1 0 1056 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1711307567
transform 1 0 760 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1711307567
transform 1 0 1152 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1711307567
transform 1 0 760 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1711307567
transform 1 0 1312 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1711307567
transform 1 0 1080 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1711307567
transform 1 0 976 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1711307567
transform 1 0 840 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1711307567
transform 1 0 824 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1711307567
transform 1 0 968 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1711307567
transform 1 0 1160 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1711307567
transform 1 0 1120 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1711307567
transform 1 0 1496 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1711307567
transform 1 0 1496 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1711307567
transform 1 0 1536 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1711307567
transform 1 0 1168 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1711307567
transform 1 0 1120 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1711307567
transform 1 0 2008 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1711307567
transform 1 0 1224 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1711307567
transform 1 0 1168 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1711307567
transform 1 0 1208 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1711307567
transform 1 0 1680 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1711307567
transform 1 0 1712 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1711307567
transform 1 0 1656 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1711307567
transform 1 0 1904 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1711307567
transform 1 0 1704 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1711307567
transform 1 0 1368 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1711307567
transform 1 0 1880 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1711307567
transform 1 0 1704 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1711307567
transform 1 0 1624 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1711307567
transform 1 0 1752 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1711307567
transform 1 0 1504 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1711307567
transform 1 0 1976 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1711307567
transform 1 0 1608 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1711307567
transform 1 0 1832 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1711307567
transform 1 0 1656 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1711307567
transform 1 0 1832 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1711307567
transform 1 0 1872 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1711307567
transform 1 0 1504 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1711307567
transform 1 0 1672 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1711307567
transform 1 0 1856 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1711307567
transform 1 0 2016 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1711307567
transform 1 0 1760 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1711307567
transform 1 0 2080 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1711307567
transform 1 0 2016 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_88
timestamp 1711307567
transform 1 0 1624 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_89
timestamp 1711307567
transform 1 0 1280 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1711307567
transform 1 0 2040 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_91
timestamp 1711307567
transform 1 0 2400 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_92
timestamp 1711307567
transform 1 0 2704 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1711307567
transform 1 0 2224 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_94
timestamp 1711307567
transform 1 0 2032 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_95
timestamp 1711307567
transform 1 0 2056 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1711307567
transform 1 0 2144 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_97
timestamp 1711307567
transform 1 0 2008 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_98
timestamp 1711307567
transform 1 0 1952 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1711307567
transform 1 0 1800 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_100
timestamp 1711307567
transform 1 0 1960 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_101
timestamp 1711307567
transform 1 0 1624 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1711307567
transform 1 0 1504 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_103
timestamp 1711307567
transform 1 0 1408 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1711307567
transform 1 0 1568 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1711307567
transform 1 0 1440 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_106
timestamp 1711307567
transform 1 0 1280 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_107
timestamp 1711307567
transform 1 0 1288 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_108
timestamp 1711307567
transform 1 0 1152 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_109
timestamp 1711307567
transform 1 0 1152 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_110
timestamp 1711307567
transform 1 0 1088 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_111
timestamp 1711307567
transform 1 0 1432 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_112
timestamp 1711307567
transform 1 0 1016 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1711307567
transform 1 0 664 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_114
timestamp 1711307567
transform 1 0 760 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_115
timestamp 1711307567
transform 1 0 888 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_116
timestamp 1711307567
transform 1 0 912 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_117
timestamp 1711307567
transform 1 0 464 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1711307567
transform 1 0 552 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_119
timestamp 1711307567
transform 1 0 296 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_120
timestamp 1711307567
transform 1 0 360 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1711307567
transform 1 0 296 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_122
timestamp 1711307567
transform 1 0 248 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1711307567
transform 1 0 344 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1711307567
transform 1 0 368 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1711307567
transform 1 0 2344 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_126
timestamp 1711307567
transform 1 0 2336 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_127
timestamp 1711307567
transform 1 0 744 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_128
timestamp 1711307567
transform 1 0 2448 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_129
timestamp 1711307567
transform 1 0 2432 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_130
timestamp 1711307567
transform 1 0 2208 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_131
timestamp 1711307567
transform 1 0 2184 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_132
timestamp 1711307567
transform 1 0 768 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_133
timestamp 1711307567
transform 1 0 1368 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_134
timestamp 1711307567
transform 1 0 2576 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_135
timestamp 1711307567
transform 1 0 2560 0 1 170
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1711307567
transform 1 0 1440 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1711307567
transform 1 0 1304 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1711307567
transform 1 0 896 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1711307567
transform 1 0 2104 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1711307567
transform 1 0 784 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1711307567
transform 1 0 760 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1711307567
transform 1 0 600 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1711307567
transform 1 0 1128 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1711307567
transform 1 0 992 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1711307567
transform 1 0 1200 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1711307567
transform 1 0 1784 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1711307567
transform 1 0 1976 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1711307567
transform 1 0 2032 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1711307567
transform 1 0 1856 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1711307567
transform 1 0 2392 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1711307567
transform 1 0 1960 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1711307567
transform 1 0 2264 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1711307567
transform 1 0 2344 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1711307567
transform 1 0 1816 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1711307567
transform 1 0 2024 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1711307567
transform 1 0 2296 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1711307567
transform 1 0 2368 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1711307567
transform 1 0 1856 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1711307567
transform 1 0 2000 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1711307567
transform 1 0 1824 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1711307567
transform 1 0 2320 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1711307567
transform 1 0 2280 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1711307567
transform 1 0 1920 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1711307567
transform 1 0 2216 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1711307567
transform 1 0 2568 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1711307567
transform 1 0 2552 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1711307567
transform 1 0 2536 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1711307567
transform 1 0 2632 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1711307567
transform 1 0 2192 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1711307567
transform 1 0 2208 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1711307567
transform 1 0 1848 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1711307567
transform 1 0 1504 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1711307567
transform 1 0 1704 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1711307567
transform 1 0 544 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1711307567
transform 1 0 344 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1711307567
transform 1 0 800 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1711307567
transform 1 0 1144 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1711307567
transform 1 0 992 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1711307567
transform 1 0 1704 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1711307567
transform 1 0 1912 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1711307567
transform 1 0 2432 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1711307567
transform 1 0 2480 0 -1 370
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1711307567
transform 1 0 2368 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1711307567
transform 1 0 2384 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1711307567
transform 1 0 360 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1711307567
transform 1 0 448 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1711307567
transform 1 0 736 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1711307567
transform 1 0 648 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1711307567
transform 1 0 632 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1711307567
transform 1 0 896 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1711307567
transform 1 0 1048 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1711307567
transform 1 0 1280 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1711307567
transform 1 0 1360 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1711307567
transform 1 0 1112 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1711307567
transform 1 0 1344 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1711307567
transform 1 0 1776 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1711307567
transform 1 0 1832 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1711307567
transform 1 0 2120 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1711307567
transform 1 0 2152 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1711307567
transform 1 0 1792 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1711307567
transform 1 0 2648 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1711307567
transform 1 0 2728 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1711307567
transform 1 0 2696 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1711307567
transform 1 0 1960 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1711307567
transform 1 0 2104 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1711307567
transform 1 0 2048 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1711307567
transform 1 0 1880 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1711307567
transform 1 0 1792 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1711307567
transform 1 0 1720 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1711307567
transform 1 0 1664 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1711307567
transform 1 0 1400 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1711307567
transform 1 0 1480 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1711307567
transform 1 0 1240 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1711307567
transform 1 0 976 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1711307567
transform 1 0 1032 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1711307567
transform 1 0 832 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1711307567
transform 1 0 568 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1711307567
transform 1 0 472 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1711307567
transform 1 0 288 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1711307567
transform 1 0 320 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1711307567
transform 1 0 688 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1711307567
transform 1 0 616 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1711307567
transform 1 0 960 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1711307567
transform 1 0 1144 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1711307567
transform 1 0 1336 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1711307567
transform 1 0 1872 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1711307567
transform 1 0 2192 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1711307567
transform 1 0 2216 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1711307567
transform 1 0 1592 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1711307567
transform 1 0 1360 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1711307567
transform 1 0 784 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1711307567
transform 1 0 240 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1711307567
transform 1 0 256 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1711307567
transform 1 0 288 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1711307567
transform 1 0 2608 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1711307567
transform 1 0 2600 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1711307567
transform 1 0 1448 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1711307567
transform 1 0 1368 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1711307567
transform 1 0 1416 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1711307567
transform 1 0 912 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1711307567
transform 1 0 680 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1711307567
transform 1 0 840 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1711307567
transform 1 0 1256 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1711307567
transform 1 0 1312 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1711307567
transform 1 0 336 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1711307567
transform 1 0 328 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1711307567
transform 1 0 288 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1711307567
transform 1 0 320 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1711307567
transform 1 0 1936 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1711307567
transform 1 0 504 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1711307567
transform 1 0 400 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1711307567
transform 1 0 504 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1711307567
transform 1 0 584 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1711307567
transform 1 0 1136 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1711307567
transform 1 0 760 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1711307567
transform 1 0 744 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1711307567
transform 1 0 616 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1711307567
transform 1 0 672 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1711307567
transform 1 0 720 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1711307567
transform 1 0 720 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1711307567
transform 1 0 608 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1711307567
transform 1 0 584 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1711307567
transform 1 0 552 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1711307567
transform 1 0 968 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1711307567
transform 1 0 848 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1711307567
transform 1 0 864 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1711307567
transform 1 0 1000 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1711307567
transform 1 0 1088 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1711307567
transform 1 0 952 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1711307567
transform 1 0 1024 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1711307567
transform 1 0 1256 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1711307567
transform 1 0 1216 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1711307567
transform 1 0 1072 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1711307567
transform 1 0 1336 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1711307567
transform 1 0 1272 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1711307567
transform 1 0 1272 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1711307567
transform 1 0 1504 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1711307567
transform 1 0 952 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1711307567
transform 1 0 1088 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1711307567
transform 1 0 1120 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1711307567
transform 1 0 936 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1711307567
transform 1 0 1320 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1711307567
transform 1 0 1288 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1711307567
transform 1 0 1136 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1711307567
transform 1 0 1424 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1711307567
transform 1 0 1520 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1711307567
transform 1 0 1480 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1711307567
transform 1 0 1480 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1711307567
transform 1 0 1456 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1711307567
transform 1 0 1368 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1711307567
transform 1 0 1752 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1711307567
transform 1 0 1552 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1711307567
transform 1 0 1704 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1711307567
transform 1 0 1696 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1711307567
transform 1 0 1560 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1711307567
transform 1 0 1352 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1711307567
transform 1 0 1856 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1711307567
transform 1 0 1768 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1711307567
transform 1 0 1768 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1711307567
transform 1 0 1600 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1711307567
transform 1 0 2096 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1711307567
transform 1 0 1952 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1711307567
transform 1 0 1912 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1711307567
transform 1 0 2176 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1711307567
transform 1 0 1968 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1711307567
transform 1 0 1992 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1711307567
transform 1 0 1816 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1711307567
transform 1 0 1656 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_126
timestamp 1711307567
transform 1 0 2120 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_127
timestamp 1711307567
transform 1 0 2192 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_128
timestamp 1711307567
transform 1 0 1656 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_129
timestamp 1711307567
transform 1 0 1712 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_130
timestamp 1711307567
transform 1 0 1952 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_131
timestamp 1711307567
transform 1 0 2208 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_132
timestamp 1711307567
transform 1 0 2624 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_133
timestamp 1711307567
transform 1 0 2360 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_134
timestamp 1711307567
transform 1 0 2168 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_135
timestamp 1711307567
transform 1 0 2200 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_136
timestamp 1711307567
transform 1 0 2720 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_137
timestamp 1711307567
transform 1 0 2608 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_138
timestamp 1711307567
transform 1 0 2280 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_139
timestamp 1711307567
transform 1 0 1888 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_140
timestamp 1711307567
transform 1 0 1584 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_141
timestamp 1711307567
transform 1 0 1632 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_142
timestamp 1711307567
transform 1 0 1608 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_143
timestamp 1711307567
transform 1 0 616 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_144
timestamp 1711307567
transform 1 0 592 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_145
timestamp 1711307567
transform 1 0 1656 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_146
timestamp 1711307567
transform 1 0 744 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_147
timestamp 1711307567
transform 1 0 488 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_148
timestamp 1711307567
transform 1 0 264 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_149
timestamp 1711307567
transform 1 0 1184 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_150
timestamp 1711307567
transform 1 0 1656 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_151
timestamp 1711307567
transform 1 0 2280 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_152
timestamp 1711307567
transform 1 0 312 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_153
timestamp 1711307567
transform 1 0 184 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_154
timestamp 1711307567
transform 1 0 104 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_155
timestamp 1711307567
transform 1 0 200 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_156
timestamp 1711307567
transform 1 0 240 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_157
timestamp 1711307567
transform 1 0 168 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_158
timestamp 1711307567
transform 1 0 528 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_159
timestamp 1711307567
transform 1 0 416 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_160
timestamp 1711307567
transform 1 0 776 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_161
timestamp 1711307567
transform 1 0 728 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_162
timestamp 1711307567
transform 1 0 624 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_163
timestamp 1711307567
transform 1 0 1048 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_164
timestamp 1711307567
transform 1 0 1040 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_165
timestamp 1711307567
transform 1 0 1088 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_166
timestamp 1711307567
transform 1 0 1128 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_167
timestamp 1711307567
transform 1 0 1216 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_168
timestamp 1711307567
transform 1 0 1576 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_169
timestamp 1711307567
transform 1 0 1368 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_170
timestamp 1711307567
transform 1 0 1432 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_171
timestamp 1711307567
transform 1 0 1720 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_172
timestamp 1711307567
transform 1 0 1872 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_173
timestamp 1711307567
transform 1 0 1840 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_174
timestamp 1711307567
transform 1 0 1936 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_175
timestamp 1711307567
transform 1 0 2000 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_176
timestamp 1711307567
transform 1 0 2064 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_177
timestamp 1711307567
transform 1 0 2656 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_178
timestamp 1711307567
transform 1 0 2632 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_179
timestamp 1711307567
transform 1 0 2488 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_180
timestamp 1711307567
transform 1 0 2264 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_181
timestamp 1711307567
transform 1 0 2464 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_182
timestamp 1711307567
transform 1 0 2576 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_183
timestamp 1711307567
transform 1 0 2304 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_184
timestamp 1711307567
transform 1 0 2272 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_185
timestamp 1711307567
transform 1 0 2400 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_186
timestamp 1711307567
transform 1 0 2600 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_187
timestamp 1711307567
transform 1 0 2104 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_188
timestamp 1711307567
transform 1 0 2368 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_189
timestamp 1711307567
transform 1 0 2664 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_190
timestamp 1711307567
transform 1 0 2720 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_191
timestamp 1711307567
transform 1 0 2608 0 -1 1770
box -8 -3 32 105
use NOR3X1  NOR3X1_0
timestamp 1711307567
transform 1 0 2232 0 -1 370
box -7 -3 68 105
use OAI21X1  OAI21X1_0
timestamp 1711307567
transform 1 0 2640 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1711307567
transform 1 0 1416 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1711307567
transform 1 0 1600 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1711307567
transform 1 0 640 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1711307567
transform 1 0 576 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1711307567
transform 1 0 1744 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1711307567
transform 1 0 1768 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1711307567
transform 1 0 1376 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1711307567
transform 1 0 1440 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1711307567
transform 1 0 952 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1711307567
transform 1 0 840 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1711307567
transform 1 0 1352 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1711307567
transform 1 0 1360 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1711307567
transform 1 0 1200 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1711307567
transform 1 0 1512 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1711307567
transform 1 0 1408 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1711307567
transform 1 0 952 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1711307567
transform 1 0 328 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1711307567
transform 1 0 1800 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1711307567
transform 1 0 720 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1711307567
transform 1 0 592 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1711307567
transform 1 0 688 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1711307567
transform 1 0 384 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1711307567
transform 1 0 1800 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1711307567
transform 1 0 1320 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1711307567
transform 1 0 1232 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1711307567
transform 1 0 1464 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1711307567
transform 1 0 1296 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1711307567
transform 1 0 176 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1711307567
transform 1 0 240 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1711307567
transform 1 0 272 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1711307567
transform 1 0 160 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1711307567
transform 1 0 208 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1711307567
transform 1 0 296 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1711307567
transform 1 0 208 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1711307567
transform 1 0 144 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1711307567
transform 1 0 184 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1711307567
transform 1 0 240 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1711307567
transform 1 0 448 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1711307567
transform 1 0 352 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1711307567
transform 1 0 632 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1711307567
transform 1 0 400 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1711307567
transform 1 0 656 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1711307567
transform 1 0 296 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1711307567
transform 1 0 632 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1711307567
transform 1 0 424 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1711307567
transform 1 0 536 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1711307567
transform 1 0 688 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1711307567
transform 1 0 704 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1711307567
transform 1 0 536 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1711307567
transform 1 0 904 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1711307567
transform 1 0 792 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1711307567
transform 1 0 1048 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1711307567
transform 1 0 1088 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1711307567
transform 1 0 1128 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1711307567
transform 1 0 912 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1711307567
transform 1 0 856 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1711307567
transform 1 0 1112 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1711307567
transform 1 0 1128 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1711307567
transform 1 0 1176 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1711307567
transform 1 0 920 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1711307567
transform 1 0 1208 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1711307567
transform 1 0 1488 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1711307567
transform 1 0 1480 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1711307567
transform 1 0 1552 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1711307567
transform 1 0 1552 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1711307567
transform 1 0 1408 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1711307567
transform 1 0 1568 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1711307567
transform 1 0 1632 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1711307567
transform 1 0 1504 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1711307567
transform 1 0 1600 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1711307567
transform 1 0 1584 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1711307567
transform 1 0 1672 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1711307567
transform 1 0 1744 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1711307567
transform 1 0 1928 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1711307567
transform 1 0 1992 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1711307567
transform 1 0 1872 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1711307567
transform 1 0 1984 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1711307567
transform 1 0 1984 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1711307567
transform 1 0 1904 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1711307567
transform 1 0 2000 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1711307567
transform 1 0 2200 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1711307567
transform 1 0 2160 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1711307567
transform 1 0 2160 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1711307567
transform 1 0 2104 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1711307567
transform 1 0 2224 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1711307567
transform 1 0 2168 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1711307567
transform 1 0 2216 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1711307567
transform 1 0 2144 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1711307567
transform 1 0 2064 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1711307567
transform 1 0 2032 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1711307567
transform 1 0 2048 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1711307567
transform 1 0 2176 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1711307567
transform 1 0 2688 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1711307567
transform 1 0 2640 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1711307567
transform 1 0 2496 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1711307567
transform 1 0 2496 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1711307567
transform 1 0 2560 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1711307567
transform 1 0 2568 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1711307567
transform 1 0 2560 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1711307567
transform 1 0 2592 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1711307567
transform 1 0 2280 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1711307567
transform 1 0 2272 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1711307567
transform 1 0 2456 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1711307567
transform 1 0 2144 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1711307567
transform 1 0 2088 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1711307567
transform 1 0 2104 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1711307567
transform 1 0 1784 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1711307567
transform 1 0 1864 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1711307567
transform 1 0 1720 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1711307567
transform 1 0 1592 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1711307567
transform 1 0 1472 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1711307567
transform 1 0 1472 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1711307567
transform 1 0 1448 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1711307567
transform 1 0 1384 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1711307567
transform 1 0 1592 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1711307567
transform 1 0 1536 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1711307567
transform 1 0 1464 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1711307567
transform 1 0 1520 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1711307567
transform 1 0 1296 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1711307567
transform 1 0 1320 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1711307567
transform 1 0 1224 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1711307567
transform 1 0 1280 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1711307567
transform 1 0 1136 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1711307567
transform 1 0 1216 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1711307567
transform 1 0 992 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1711307567
transform 1 0 1168 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1711307567
transform 1 0 1048 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1711307567
transform 1 0 1384 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1711307567
transform 1 0 1544 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1711307567
transform 1 0 1072 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1711307567
transform 1 0 960 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1711307567
transform 1 0 984 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1711307567
transform 1 0 664 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1711307567
transform 1 0 760 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1711307567
transform 1 0 744 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1711307567
transform 1 0 824 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1711307567
transform 1 0 856 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1711307567
transform 1 0 880 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1711307567
transform 1 0 864 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1711307567
transform 1 0 920 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1711307567
transform 1 0 456 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1711307567
transform 1 0 472 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1711307567
transform 1 0 576 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1711307567
transform 1 0 536 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1711307567
transform 1 0 216 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1711307567
transform 1 0 392 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1711307567
transform 1 0 336 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1711307567
transform 1 0 424 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1711307567
transform 1 0 664 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1711307567
transform 1 0 784 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1711307567
transform 1 0 232 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1711307567
transform 1 0 288 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1711307567
transform 1 0 192 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1711307567
transform 1 0 264 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1711307567
transform 1 0 208 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1711307567
transform 1 0 352 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1711307567
transform 1 0 416 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1711307567
transform 1 0 368 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1711307567
transform 1 0 2624 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1711307567
transform 1 0 2552 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1711307567
transform 1 0 2472 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1711307567
transform 1 0 2592 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_163
timestamp 1711307567
transform 1 0 2600 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_164
timestamp 1711307567
transform 1 0 1480 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_165
timestamp 1711307567
transform 1 0 2592 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_166
timestamp 1711307567
transform 1 0 2544 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_167
timestamp 1711307567
transform 1 0 2520 0 1 170
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1711307567
transform 1 0 1048 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1711307567
transform 1 0 544 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1711307567
transform 1 0 384 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1711307567
transform 1 0 1920 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1711307567
transform 1 0 1400 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1711307567
transform 1 0 1328 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1711307567
transform 1 0 1200 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1711307567
transform 1 0 776 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1711307567
transform 1 0 1032 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1711307567
transform 1 0 704 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1711307567
transform 1 0 864 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1711307567
transform 1 0 1200 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1711307567
transform 1 0 1904 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1711307567
transform 1 0 440 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1711307567
transform 1 0 736 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1711307567
transform 1 0 664 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1711307567
transform 1 0 688 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1711307567
transform 1 0 968 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1711307567
transform 1 0 896 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1711307567
transform 1 0 992 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1711307567
transform 1 0 1248 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1711307567
transform 1 0 1040 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1711307567
transform 1 0 1288 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1711307567
transform 1 0 1544 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1711307567
transform 1 0 1608 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1711307567
transform 1 0 1808 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1711307567
transform 1 0 2080 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1711307567
transform 1 0 2048 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1711307567
transform 1 0 1808 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1711307567
transform 1 0 1880 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1711307567
transform 1 0 1968 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1711307567
transform 1 0 2040 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1711307567
transform 1 0 2512 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1711307567
transform 1 0 2608 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1711307567
transform 1 0 2480 0 -1 170
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1711307567
transform 1 0 1272 0 -1 2370
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1711307567
transform 1 0 960 0 -1 2370
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1711307567
transform 1 0 176 0 -1 1970
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1711307567
transform 1 0 2464 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1711307567
transform 1 0 1024 0 1 570
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1711307567
transform 1 0 816 0 1 770
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1711307567
transform 1 0 2312 0 1 170
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1711307567
transform 1 0 2624 0 -1 370
box -8 -3 40 105
use OR2X2  OR2X2_0
timestamp 1711307567
transform 1 0 1752 0 -1 1770
box -7 -3 35 105
use OR2X2  OR2X2_1
timestamp 1711307567
transform 1 0 664 0 -1 1770
box -7 -3 35 105
use OR2X2  OR2X2_2
timestamp 1711307567
transform 1 0 2248 0 1 170
box -7 -3 35 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1711307567
transform 1 0 2808 0 1 2617
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1711307567
transform 1 0 2808 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1711307567
transform 1 0 24 0 1 2617
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1711307567
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1711307567
transform 1 0 2784 0 1 2593
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1711307567
transform 1 0 2784 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1711307567
transform 1 0 48 0 1 2593
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1711307567
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1711307567
transform 1 0 2808 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1711307567
transform 1 0 2808 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1711307567
transform 1 0 2808 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1711307567
transform 1 0 2808 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1711307567
transform 1 0 2808 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1711307567
transform 1 0 2808 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1711307567
transform 1 0 2808 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1711307567
transform 1 0 2808 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1711307567
transform 1 0 2808 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1711307567
transform 1 0 2808 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1711307567
transform 1 0 2808 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1711307567
transform 1 0 2808 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1711307567
transform 1 0 2808 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1711307567
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1711307567
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1711307567
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1711307567
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1711307567
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1711307567
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1711307567
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1711307567
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1711307567
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1711307567
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1711307567
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1711307567
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1711307567
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1711307567
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1711307567
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1711307567
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1711307567
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1711307567
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1711307567
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1711307567
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1711307567
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1711307567
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1711307567
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1711307567
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1711307567
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1711307567
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1711307567
transform 1 0 2784 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1711307567
transform 1 0 2784 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1711307567
transform 1 0 2784 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1711307567
transform 1 0 2784 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1711307567
transform 1 0 2784 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1711307567
transform 1 0 2784 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1711307567
transform 1 0 2784 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1711307567
transform 1 0 2784 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1711307567
transform 1 0 2784 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1711307567
transform 1 0 2784 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1711307567
transform 1 0 2784 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_50
timestamp 1711307567
transform 1 0 2784 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_51
timestamp 1711307567
transform 1 0 2784 0 1 2570
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1711307567
transform 1 0 2704 0 1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1711307567
transform 1 0 2104 0 -1 2570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1711307567
transform 1 0 2120 0 1 2370
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1711307567
transform 1 0 2552 0 1 2370
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1711307567
transform 1 0 2608 0 -1 2570
box -8 -3 64 105
<< labels >>
rlabel metal1 2708 605 2708 605 4 in_clka
rlabel electrodecontact s 1500 1125 1500 1125 4 in_clkb
rlabel electrodecontact s 2452 2135 2452 2135 4 in_restart
rlabel electrodecontact s 2708 1735 2708 1735 4 in_move[1]
rlabel electrodecontact s 2652 1735 2652 1735 4 in_move[0]
rlabel electrodecontact s 388 1125 388 1125 4 board_out[31]
rlabel metal1 300 1125 300 1125 4 board_out[30]
rlabel metal1 276 1525 276 1525 4 board_out[29]
rlabel electrodecontact s 260 1525 260 1525 4 board_out[28]
rlabel electrodecontact s 468 725 468 725 4 board_out[27]
rlabel metal1 484 725 484 725 4 board_out[26]
rlabel metal1 468 815 468 815 4 board_out[25]
rlabel electrodecontact s 484 925 484 925 4 board_out[24]
rlabel electrodecontact s 724 925 724 925 4 board_out[23]
rlabel metal1 628 1015 628 1015 4 board_out[22]
rlabel metal1 556 1125 556 1125 4 board_out[21]
rlabel metal1 908 925 908 925 4 board_out[20]
rlabel metal1 932 925 932 925 4 board_out[19]
rlabel metal1 964 815 964 815 4 board_out[18]
rlabel metal1 1188 925 1188 925 4 board_out[17]
rlabel electrodecontact s 1284 925 1284 925 4 board_out[16]
rlabel metal1 1100 815 1100 815 4 board_out[15]
rlabel metal1 1116 815 1116 815 4 board_out[14]
rlabel metal1 1236 725 1236 725 4 board_out[13]
rlabel metal1 1260 725 1260 725 4 board_out[12]
rlabel electrodecontact s 1668 525 1668 525 4 board_out[11]
rlabel metal1 1788 415 1788 415 4 board_out[10]
rlabel electrodecontact s 1708 815 1708 815 4 board_out[9]
rlabel metal1 1748 615 1748 615 4 board_out[8]
rlabel metal1 1948 1015 1948 1015 4 board_out[7]
rlabel electrodecontact s 2340 1325 2340 1325 4 board_out[6]
rlabel metal1 2484 1325 2484 1325 4 board_out[5]
rlabel metal1 2284 1215 2284 1215 4 board_out[4]
rlabel metal1 2004 1015 2004 1015 4 board_out[3]
rlabel electrodecontact s 2204 925 2204 925 4 board_out[2]
rlabel metal1 2324 815 2324 815 4 board_out[1]
rlabel metal1 2084 1015 2084 1015 4 board_out[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 24228.000 19575.000 24300.000 19575.000 
<< end >>
