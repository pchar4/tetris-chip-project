magic
tech scmos
timestamp 1713453518
<< m2contact >>
rect -2 -2 2 2
<< end >>
