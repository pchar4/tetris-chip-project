magic
tech scmos
timestamp 1713453518
<< metal1 >>
rect 14 3407 3506 3427
rect 38 3383 3482 3403
rect 38 3367 3482 3373
rect 1850 3343 1876 3346
rect 2194 3343 2204 3346
rect 2442 3343 2468 3346
rect 186 3326 189 3335
rect 244 3333 269 3336
rect 610 3326 613 3335
rect 652 3333 661 3336
rect 668 3333 685 3336
rect 1106 3333 1124 3336
rect 1188 3333 1196 3336
rect 1266 3326 1269 3335
rect 1292 3333 1316 3336
rect 1330 3333 1348 3336
rect 1378 3326 1381 3335
rect 1404 3333 1445 3336
rect 1650 3333 1708 3336
rect 1826 3326 1829 3335
rect 1834 3333 1925 3336
rect 2122 3333 2156 3336
rect 2178 3333 2212 3336
rect 2434 3333 2533 3336
rect 2570 3333 2588 3336
rect 2676 3333 2733 3336
rect 2756 3333 2789 3336
rect 2794 3333 2804 3336
rect 2818 3333 2860 3336
rect 3010 3333 3044 3336
rect 3068 3333 3100 3336
rect 3124 3333 3133 3336
rect 3170 3333 3180 3336
rect 3252 3333 3285 3336
rect 3314 3333 3324 3336
rect 108 3323 133 3326
rect 164 3323 189 3326
rect 196 3323 212 3326
rect 252 3323 269 3326
rect 404 3323 429 3326
rect 460 3323 469 3326
rect 540 3323 565 3326
rect 596 3323 613 3326
rect 620 3323 636 3326
rect 820 3323 845 3326
rect 948 3323 957 3326
rect 1044 3323 1069 3326
rect 1114 3323 1132 3326
rect 1154 3323 1172 3326
rect 1204 3323 1245 3326
rect 1252 3323 1269 3326
rect 1306 3323 1324 3326
rect 1370 3323 1381 3326
rect 1716 3323 1725 3326
rect 1770 3323 1812 3326
rect 1826 3323 1845 3326
rect 1892 3323 1901 3326
rect 1922 3323 1925 3333
rect 2530 3326 2533 3333
rect 2786 3326 2789 3333
rect 1970 3323 1996 3326
rect 2010 3323 2092 3326
rect 2164 3323 2205 3326
rect 2268 3323 2332 3326
rect 2364 3323 2428 3326
rect 2530 3323 2541 3326
rect 2562 3323 2596 3326
rect 2602 3323 2652 3326
rect 2714 3323 2732 3326
rect 2786 3323 2812 3326
rect 2826 3323 2852 3326
rect 2986 3323 3004 3326
rect 3082 3323 3108 3326
rect 3162 3323 3188 3326
rect 3258 3323 3284 3326
rect 3308 3323 3325 3326
rect 3346 3323 3356 3326
rect 1292 3313 1301 3316
rect 2012 3313 2029 3316
rect 2370 3303 2373 3323
rect 2604 3313 2645 3316
rect 2890 3313 2908 3316
rect 2938 3313 2956 3316
rect 2938 3303 2972 3306
rect 3194 3303 3212 3306
rect 14 3267 3506 3273
rect 3050 3233 3100 3236
rect 3154 3226 3157 3246
rect 3194 3233 3204 3236
rect 468 3223 509 3226
rect 1100 3223 1117 3226
rect 1220 3223 1245 3226
rect 1268 3223 1293 3226
rect 1340 3223 1349 3226
rect 1796 3223 1829 3226
rect 2516 3223 2565 3226
rect 2596 3223 2629 3226
rect 3074 3223 3084 3226
rect 3108 3223 3125 3226
rect 3140 3223 3157 3226
rect 3170 3223 3197 3226
rect 3274 3216 3277 3236
rect 204 3213 229 3216
rect 332 3213 357 3216
rect 388 3213 429 3216
rect 436 3213 452 3216
rect 548 3213 573 3216
rect 604 3213 629 3216
rect 636 3213 645 3216
rect 660 3213 677 3216
rect 780 3213 805 3216
rect 844 3213 853 3216
rect 882 3213 908 3216
rect 940 3213 965 3216
rect 1004 3213 1021 3216
rect 1050 3213 1084 3216
rect 1178 3213 1212 3216
rect 1260 3213 1309 3216
rect 1388 3213 1405 3216
rect 1460 3213 1509 3216
rect 1650 3213 1717 3216
rect 1724 3213 1765 3216
rect 1770 3213 1780 3216
rect 1892 3213 1909 3216
rect 1978 3213 2044 3216
rect 2076 3213 2085 3216
rect 2090 3213 2164 3216
rect 2188 3213 2261 3216
rect 2292 3213 2349 3216
rect 2354 3213 2372 3216
rect 2514 3213 2588 3216
rect 2594 3213 2644 3216
rect 2658 3213 2716 3216
rect 2786 3213 2836 3216
rect 2866 3213 2876 3216
rect 2906 3213 2940 3216
rect 2980 3213 3029 3216
rect 3114 3213 3132 3216
rect 3268 3213 3277 3216
rect 426 3205 429 3213
rect 626 3205 629 3213
rect 642 3195 645 3213
rect 1394 3206 1397 3213
rect 652 3203 685 3206
rect 810 3203 820 3206
rect 842 3203 852 3206
rect 906 3203 916 3206
rect 938 3203 980 3206
rect 1002 3203 1028 3206
rect 1042 3203 1076 3206
rect 1156 3203 1197 3206
rect 1218 3203 1252 3206
rect 1266 3203 1316 3206
rect 1340 3203 1365 3206
rect 1394 3203 1436 3206
rect 1506 3203 1524 3206
rect 1644 3203 1661 3206
rect 1714 3205 1717 3213
rect 2354 3206 2357 3213
rect 2786 3206 2789 3213
rect 1802 3203 1884 3206
rect 2018 3203 2052 3206
rect 2068 3203 2077 3206
rect 2186 3203 2268 3206
rect 2298 3203 2357 3206
rect 2370 3203 2380 3206
rect 2522 3203 2580 3206
rect 2594 3203 2636 3206
rect 2706 3203 2724 3206
rect 2740 3203 2789 3206
rect 2794 3203 2828 3206
rect 2858 3203 2868 3206
rect 2882 3203 2932 3206
rect 2946 3203 2972 3206
rect 3026 3196 3029 3213
rect 3036 3203 3069 3206
rect 3218 3203 3244 3206
rect 3290 3203 3308 3206
rect 3324 3203 3333 3206
rect 3362 3203 3380 3206
rect 1106 3193 1148 3196
rect 1810 3193 1876 3196
rect 1890 3193 1948 3196
rect 3010 3195 3029 3196
rect 3010 3193 3028 3195
rect 38 3167 3482 3173
rect 282 3143 300 3146
rect 1914 3136 1917 3146
rect 2202 3143 2220 3146
rect 2346 3143 2397 3146
rect 3162 3143 3196 3146
rect 308 3133 381 3136
rect 548 3133 589 3136
rect 626 3133 652 3136
rect 1082 3133 1100 3136
rect 1170 3133 1188 3136
rect 1220 3133 1229 3136
rect 1250 3133 1284 3136
rect 1324 3133 1333 3136
rect 1388 3133 1405 3136
rect 1426 3133 1444 3136
rect 1468 3133 1493 3136
rect 1498 3133 1516 3136
rect 1540 3133 1557 3136
rect 1562 3133 1596 3136
rect 1650 3133 1692 3136
rect 1796 3133 1876 3136
rect 1908 3133 1917 3136
rect 2068 3133 2093 3136
rect 2098 3133 2140 3136
rect 2164 3133 2189 3136
rect 2194 3133 2228 3136
rect 2394 3133 2404 3136
rect 2426 3133 2452 3136
rect 2540 3133 2549 3136
rect 2554 3133 2612 3136
rect 2636 3133 2677 3136
rect 2708 3133 2765 3136
rect 2796 3133 2829 3136
rect 2860 3133 2925 3136
rect 2954 3133 3020 3136
rect 3050 3133 3108 3136
rect 3122 3133 3132 3136
rect 3146 3133 3204 3136
rect 3226 3133 3237 3136
rect 116 3123 133 3126
rect 244 3123 260 3126
rect 476 3123 501 3126
rect 514 3123 524 3126
rect 618 3123 644 3126
rect 692 3123 733 3126
rect 772 3123 797 3126
rect 834 3123 876 3126
rect 948 3123 981 3126
rect 1020 3123 1037 3126
rect 1082 3123 1108 3126
rect 1196 3123 1205 3126
rect 1292 3123 1301 3126
rect 1354 3123 1372 3126
rect 1402 3123 1420 3126
rect 1442 3123 1452 3126
rect 1570 3123 1604 3126
rect 1626 3123 1685 3126
rect 1738 3123 1772 3126
rect 2138 3123 2148 3126
rect 2250 3123 2300 3126
rect 2332 3123 2389 3126
rect 2442 3123 2460 3126
rect 2466 3123 2524 3126
rect 2802 3123 2844 3126
rect 2954 3125 2957 3133
rect 3226 3126 3229 3133
rect 3124 3123 3133 3126
rect 3220 3123 3229 3126
rect 3274 3123 3284 3126
rect 3290 3123 3300 3126
rect 3428 3123 3445 3126
rect 514 3103 517 3123
rect 1402 3116 1405 3123
rect 620 3113 637 3116
rect 1324 3113 1349 3116
rect 1388 3113 1405 3116
rect 1468 3113 1493 3116
rect 1540 3113 1549 3116
rect 2004 3113 2053 3116
rect 2420 3113 2445 3116
rect 2636 3113 2645 3116
rect 14 3067 3506 3073
rect 1714 3033 1796 3036
rect 2658 3033 2748 3036
rect 604 3023 629 3026
rect 1068 3023 1109 3026
rect 1460 3023 1501 3026
rect 1596 3023 1629 3026
rect 1706 3023 1780 3026
rect 1804 3023 1853 3026
rect 2220 3023 2293 3026
rect 2476 3023 2525 3026
rect 2658 3023 2732 3026
rect 148 3013 204 3016
rect 218 3013 229 3016
rect 244 3013 261 3016
rect 388 3013 445 3016
rect 514 3013 524 3016
rect 610 3013 644 3016
rect 706 3013 756 3016
rect 788 3013 805 3016
rect 844 3013 877 3016
rect 916 3013 941 3016
rect 1034 3013 1045 3016
rect 1082 3013 1124 3016
rect 1156 3013 1197 3016
rect 1212 3013 1253 3016
rect 1268 3013 1293 3016
rect 1324 3013 1357 3016
rect 1388 3013 1437 3016
rect 1546 3013 1580 3016
rect 226 2995 229 3013
rect 236 3003 285 3006
rect 476 3003 501 3006
rect 506 3003 532 3006
rect 562 3003 580 3006
rect 706 3003 764 3006
rect 794 3003 820 3006
rect 986 3003 1012 3006
rect 1042 3005 1045 3013
rect 1354 3006 1357 3013
rect 1178 3003 1204 3006
rect 1266 3003 1300 3006
rect 1354 3003 1372 3006
rect 1386 3003 1436 3006
rect 1460 3003 1469 3006
rect 1538 3003 1572 3006
rect 1626 3003 1629 3023
rect 1634 3013 1676 3016
rect 2116 3013 2157 3016
rect 2290 3006 2293 3023
rect 2770 3016 2773 3056
rect 3194 3033 3220 3036
rect 3194 3026 3197 3033
rect 3108 3023 3125 3026
rect 3172 3023 3197 3026
rect 3228 3023 3253 3026
rect 3324 3023 3333 3026
rect 3250 3016 3253 3023
rect 2412 3013 2437 3016
rect 2482 3013 2540 3016
rect 2602 3013 2620 3016
rect 2652 3013 2725 3016
rect 2770 3013 2781 3016
rect 2794 3013 2844 3016
rect 2980 3013 3005 3016
rect 1642 3003 1668 3006
rect 1700 3003 1749 3006
rect 1810 3003 1860 3006
rect 1932 3003 1989 3006
rect 2010 3003 2092 3006
rect 2170 3003 2196 3006
rect 2220 3003 2285 3006
rect 2290 3003 2308 3006
rect 2354 3003 2404 3006
rect 2426 3003 2460 3006
rect 2474 3003 2532 3006
rect 2610 3003 2628 3006
rect 2778 3005 2781 3013
rect 2810 3003 2851 3006
rect 2914 3003 2956 3006
rect 1234 2993 1252 2996
rect 1388 2993 1429 2996
rect 1914 2993 1924 2996
rect 2378 2993 2396 2996
rect 3002 2995 3005 3013
rect 3058 3013 3069 3016
rect 3250 3013 3260 3016
rect 3284 3013 3293 3016
rect 3338 3013 3356 3016
rect 3380 3013 3389 3016
rect 3058 3006 3061 3013
rect 3012 3003 3061 3006
rect 3108 3003 3117 3006
rect 3146 3003 3156 3006
rect 3242 3003 3268 3006
rect 3282 2995 3285 3006
rect 3298 3003 3308 3006
rect 3378 3003 3388 3006
rect 2122 2983 2181 2986
rect 2810 2983 2837 2986
rect 38 2967 3482 2973
rect 2362 2953 2397 2956
rect 1322 2943 1348 2946
rect 2058 2943 2108 2946
rect 194 2926 197 2935
rect 252 2933 277 2936
rect 484 2933 525 2936
rect 594 2933 620 2936
rect 706 2933 716 2936
rect 1034 2933 1044 2936
rect 1100 2933 1133 2936
rect 116 2923 133 2926
rect 172 2923 197 2926
rect 204 2923 220 2926
rect 372 2923 381 2926
rect 442 2923 452 2926
rect 498 2923 540 2926
rect 698 2923 708 2926
rect 756 2923 789 2926
rect 828 2923 853 2926
rect 972 2923 997 2926
rect 1042 2923 1052 2926
rect 1138 2923 1141 2934
rect 1164 2933 1173 2936
rect 1204 2933 1245 2936
rect 1308 2933 1349 2936
rect 1362 2933 1380 2936
rect 1410 2933 1428 2936
rect 1452 2933 1485 2936
rect 1532 2933 1565 2936
rect 1636 2933 1669 2936
rect 1682 2933 1724 2936
rect 1740 2933 1797 2936
rect 1162 2923 1173 2926
rect 1234 2923 1260 2926
rect 1362 2925 1365 2933
rect 1842 2926 1845 2935
rect 1850 2933 1916 2936
rect 1986 2933 2020 2936
rect 2122 2933 2132 2936
rect 2146 2933 2220 2936
rect 2340 2933 2373 2936
rect 2450 2933 2476 2936
rect 2610 2933 2620 2936
rect 2636 2933 2653 2936
rect 2722 2933 2756 2936
rect 2780 2933 2813 2936
rect 2866 2933 2885 2936
rect 2922 2926 2925 2936
rect 2938 2933 2948 2936
rect 3114 2926 3117 2934
rect 3140 2933 3181 2936
rect 3210 2933 3220 2936
rect 3242 2933 3284 2936
rect 3332 2933 3365 2936
rect 3402 2933 3420 2936
rect 1402 2923 1436 2926
rect 1546 2923 1612 2926
rect 1650 2923 1716 2926
rect 1748 2923 1765 2926
rect 1842 2923 1861 2926
rect 1946 2923 2012 2926
rect 2044 2923 2053 2926
rect 2124 2923 2140 2926
rect 2170 2923 2212 2926
rect 2244 2923 2253 2926
rect 2258 2923 2316 2926
rect 644 2913 661 2916
rect 916 2913 933 2916
rect 658 2906 661 2913
rect 658 2903 677 2906
rect 1170 2893 1173 2923
rect 1452 2913 1469 2916
rect 1844 2913 1893 2916
rect 2162 2913 2189 2916
rect 2386 2913 2412 2916
rect 2418 2906 2421 2925
rect 2484 2923 2548 2926
rect 2602 2923 2612 2926
rect 2644 2923 2669 2926
rect 2810 2923 2828 2926
rect 2890 2923 2915 2926
rect 2922 2923 2956 2926
rect 3012 2923 3029 2926
rect 3100 2923 3117 2926
rect 3228 2923 3237 2926
rect 3292 2923 3301 2926
rect 3340 2923 3357 2926
rect 3362 2925 3365 2933
rect 3396 2923 3405 2926
rect 3410 2923 3428 2926
rect 2436 2913 2469 2916
rect 2492 2913 2533 2916
rect 2658 2913 2692 2916
rect 2780 2913 2797 2916
rect 3018 2913 3036 2916
rect 2410 2903 2421 2906
rect 2450 2903 2477 2906
rect 2666 2903 2708 2906
rect 1658 2893 1709 2896
rect 14 2867 3506 2873
rect 1442 2833 1468 2836
rect 2386 2833 2429 2836
rect 3130 2833 3172 2836
rect 860 2823 869 2826
rect 1340 2823 1357 2826
rect 116 2813 133 2816
rect 172 2813 213 2816
rect 220 2813 236 2816
rect 276 2813 301 2816
rect 404 2813 437 2816
rect 476 2813 485 2816
rect 538 2813 556 2816
rect 602 2813 628 2816
rect 666 2813 676 2816
rect 882 2813 916 2816
rect 956 2813 1029 2816
rect 1050 2813 1084 2816
rect 1116 2813 1173 2816
rect 1180 2813 1189 2816
rect 210 2805 213 2813
rect 268 2803 309 2806
rect 468 2803 508 2806
rect 524 2803 549 2806
rect 652 2803 661 2806
rect 810 2803 836 2806
rect 1052 2803 1069 2806
rect 1170 2805 1173 2813
rect 1186 2805 1189 2813
rect 1210 2813 1261 2816
rect 1282 2813 1324 2816
rect 1346 2813 1373 2816
rect 1380 2813 1405 2816
rect 1210 2805 1213 2813
rect 1442 2806 1445 2833
rect 1476 2823 1509 2826
rect 1676 2823 1685 2826
rect 1940 2823 1997 2826
rect 2082 2823 2109 2826
rect 2274 2823 2340 2826
rect 2364 2823 2373 2826
rect 2378 2823 2420 2826
rect 2444 2823 2453 2826
rect 2588 2823 2613 2826
rect 2618 2823 2645 2826
rect 3036 2823 3045 2826
rect 3124 2823 3156 2826
rect 2106 2816 2109 2823
rect 1490 2813 1524 2816
rect 1562 2813 1653 2816
rect 1740 2813 1797 2816
rect 1818 2813 1852 2816
rect 1866 2813 1932 2816
rect 2004 2813 2053 2816
rect 2060 2813 2101 2816
rect 2106 2813 2124 2816
rect 2268 2813 2333 2816
rect 1284 2803 1293 2806
rect 1298 2803 1316 2806
rect 1354 2803 1372 2806
rect 1412 2803 1445 2806
rect 1498 2803 1516 2806
rect 1540 2803 1573 2806
rect 1674 2803 1732 2806
rect 1794 2805 1797 2813
rect 1810 2803 1844 2806
rect 1946 2803 1996 2806
rect 2010 2803 2052 2806
rect 2114 2803 2132 2806
rect 2162 2803 2244 2806
rect 1386 2793 1404 2796
rect 2450 2793 2453 2823
rect 2498 2813 2508 2816
rect 2546 2813 2580 2816
rect 2602 2813 2652 2816
rect 2666 2813 2684 2816
rect 2724 2813 2749 2816
rect 2756 2813 2773 2816
rect 2876 2813 2885 2816
rect 2898 2813 2908 2816
rect 3028 2813 3037 2816
rect 3090 2813 3101 2816
rect 3212 2813 3237 2816
rect 3244 2813 3269 2816
rect 3300 2813 3317 2816
rect 3324 2813 3341 2816
rect 2498 2783 2501 2813
rect 2506 2803 2516 2806
rect 2532 2803 2565 2806
rect 2594 2803 2644 2806
rect 2698 2803 2716 2806
rect 2722 2803 2748 2806
rect 2780 2803 2797 2806
rect 2836 2803 2853 2806
rect 2930 2803 2940 2806
rect 3034 2803 3068 2806
rect 3098 2805 3101 2813
rect 3124 2803 3149 2806
rect 3258 2803 3268 2806
rect 3306 2803 3316 2806
rect 3330 2803 3356 2806
rect 3386 2803 3396 2806
rect 3420 2803 3429 2806
rect 3436 2803 3445 2806
rect 2850 2796 2853 2803
rect 2786 2793 2805 2796
rect 3426 2795 3429 2803
rect 38 2767 3482 2773
rect 522 2743 532 2746
rect 834 2736 837 2756
rect 2570 2743 2612 2746
rect 2746 2736 2749 2756
rect 3228 2743 3237 2746
rect 250 2726 253 2734
rect 308 2733 357 2736
rect 466 2733 492 2736
rect 516 2733 533 2736
rect 546 2733 588 2736
rect 618 2733 628 2736
rect 634 2733 684 2736
rect 700 2733 725 2736
rect 730 2733 748 2736
rect 778 2733 804 2736
rect 828 2733 837 2736
rect 850 2733 860 2736
rect 882 2733 892 2736
rect 1042 2733 1068 2736
rect 140 2723 165 2726
rect 196 2723 253 2726
rect 260 2723 276 2726
rect 452 2723 485 2726
rect 500 2723 509 2726
rect 546 2725 549 2733
rect 1098 2726 1101 2734
rect 1178 2733 1204 2736
rect 1226 2734 1244 2736
rect 1226 2733 1245 2734
rect 1268 2733 1293 2736
rect 1298 2733 1316 2736
rect 1386 2733 1420 2736
rect 1458 2733 1532 2736
rect 1546 2733 1588 2736
rect 1602 2733 1628 2736
rect 1642 2733 1693 2736
rect 1836 2733 1853 2736
rect 1874 2733 1892 2736
rect 1922 2733 1988 2736
rect 2170 2733 2212 2736
rect 2306 2733 2332 2736
rect 2348 2733 2405 2736
rect 2452 2733 2509 2736
rect 2514 2733 2540 2736
rect 2620 2733 2645 2736
rect 2650 2733 2660 2736
rect 2738 2733 2749 2736
rect 2826 2733 2837 2736
rect 2882 2733 2908 2736
rect 2978 2733 2996 2736
rect 3018 2733 3036 2736
rect 3124 2733 3149 2736
rect 3186 2733 3212 2736
rect 3274 2733 3284 2736
rect 3306 2733 3332 2736
rect 3346 2733 3364 2736
rect 3386 2733 3412 2736
rect 1242 2726 1245 2733
rect 714 2723 740 2726
rect 834 2723 852 2726
rect 884 2723 893 2726
rect 980 2723 1005 2726
rect 1036 2723 1045 2726
rect 1050 2723 1076 2726
rect 1090 2723 1101 2726
rect 1108 2723 1149 2726
rect 1164 2723 1189 2726
rect 1212 2723 1245 2726
rect 1252 2723 1261 2726
rect 1298 2716 1301 2733
rect 1642 2726 1645 2733
rect 1306 2723 1356 2726
rect 1394 2723 1428 2726
rect 1500 2723 1533 2726
rect 1540 2723 1581 2726
rect 1596 2723 1629 2726
rect 1636 2723 1645 2726
rect 1650 2723 1716 2726
rect 1882 2723 1900 2726
rect 1930 2723 1980 2726
rect 2026 2723 2084 2726
rect 2098 2723 2140 2726
rect 2172 2723 2181 2726
rect 2220 2723 2245 2726
rect 2258 2723 2324 2726
rect 2356 2723 2373 2726
rect 2402 2723 2428 2726
rect 2460 2723 2485 2726
rect 2490 2723 2532 2726
rect 828 2713 837 2716
rect 1172 2713 1205 2716
rect 1220 2713 1237 2716
rect 1298 2713 1309 2716
rect 1836 2713 1885 2716
rect 1916 2713 1965 2716
rect 2092 2713 2125 2716
rect 2178 2703 2181 2723
rect 2242 2703 2245 2723
rect 2260 2713 2285 2716
rect 2490 2706 2493 2723
rect 2690 2713 2708 2716
rect 2466 2703 2493 2706
rect 2746 2703 2780 2706
rect 2826 2703 2829 2733
rect 2882 2726 2885 2733
rect 3018 2726 3021 2733
rect 2868 2723 2885 2726
rect 2890 2723 2900 2726
rect 2970 2723 3021 2726
rect 3068 2723 3077 2726
rect 3090 2723 3100 2726
rect 2964 2713 2973 2716
rect 3090 2713 3093 2723
rect 3138 2703 3141 2726
rect 3186 2716 3189 2733
rect 3346 2726 3349 2733
rect 3228 2723 3261 2726
rect 3282 2723 3292 2726
rect 3340 2723 3349 2726
rect 3180 2713 3189 2716
rect 3154 2703 3172 2706
rect 14 2667 3506 2673
rect 2882 2643 2901 2646
rect 2090 2633 2132 2636
rect 2538 2633 2588 2636
rect 1084 2623 1093 2626
rect 1380 2623 1397 2626
rect 1540 2623 1549 2626
rect 1612 2623 1653 2626
rect 1740 2623 1757 2626
rect 1810 2623 1829 2626
rect 1852 2623 1893 2626
rect 2076 2623 2101 2626
rect 2116 2623 2125 2626
rect 2140 2623 2149 2626
rect 2554 2623 2572 2626
rect 2596 2623 2605 2626
rect 1810 2616 1813 2623
rect 124 2613 149 2616
rect 180 2613 205 2616
rect 210 2613 228 2616
rect 234 2613 244 2616
rect 260 2613 284 2616
rect 298 2613 309 2616
rect 404 2613 413 2616
rect 460 2613 477 2616
rect 516 2613 525 2616
rect 266 2603 276 2606
rect 306 2595 309 2613
rect 538 2606 541 2614
rect 570 2606 573 2614
rect 316 2603 365 2606
rect 514 2603 541 2606
rect 562 2603 573 2606
rect 594 2606 597 2614
rect 772 2613 781 2616
rect 810 2613 828 2616
rect 940 2613 965 2616
rect 1002 2613 1036 2616
rect 1140 2613 1173 2616
rect 1210 2613 1252 2616
rect 1274 2613 1292 2616
rect 1316 2613 1364 2616
rect 1420 2613 1469 2616
rect 1532 2613 1541 2616
rect 1554 2613 1596 2616
rect 1684 2613 1717 2616
rect 1722 2613 1797 2616
rect 1804 2613 1813 2616
rect 1818 2613 1844 2616
rect 2026 2613 2068 2616
rect 1794 2606 1797 2613
rect 594 2603 636 2606
rect 730 2603 748 2606
rect 770 2603 780 2606
rect 804 2603 821 2606
rect 1018 2603 1028 2606
rect 1084 2603 1125 2606
rect 1162 2603 1172 2606
rect 1268 2603 1285 2606
rect 1290 2603 1300 2606
rect 1330 2603 1356 2606
rect 1380 2603 1389 2606
rect 1402 2603 1412 2606
rect 1458 2603 1468 2606
rect 1492 2603 1517 2606
rect 1538 2603 1588 2606
rect 1612 2603 1668 2606
rect 1706 2603 1724 2606
rect 1754 2605 1797 2606
rect 1754 2603 1796 2605
rect 1850 2603 1916 2606
rect 1986 2603 1996 2606
rect 2026 2603 2060 2606
rect 2146 2603 2149 2623
rect 2882 2616 2885 2643
rect 2898 2633 2925 2636
rect 2890 2623 2901 2626
rect 2906 2623 2916 2626
rect 2220 2613 2229 2616
rect 2268 2613 2277 2616
rect 2316 2613 2341 2616
rect 2402 2613 2444 2616
rect 2490 2613 2524 2616
rect 2610 2613 2660 2616
rect 2666 2613 2676 2616
rect 2794 2613 2813 2616
rect 2844 2613 2861 2616
rect 2868 2613 2877 2616
rect 2882 2613 2893 2616
rect 2490 2606 2493 2613
rect 2874 2606 2877 2613
rect 2898 2606 2901 2623
rect 2922 2615 2925 2633
rect 3228 2623 3245 2626
rect 3282 2616 3285 2625
rect 2964 2613 2973 2616
rect 2986 2613 3012 2616
rect 3036 2613 3045 2616
rect 3138 2613 3188 2616
rect 3234 2613 3276 2616
rect 3282 2613 3293 2616
rect 3300 2613 3317 2616
rect 3410 2613 3428 2616
rect 2186 2603 2204 2606
rect 2226 2603 2253 2606
rect 2260 2603 2308 2606
rect 2372 2603 2389 2606
rect 2468 2603 2501 2606
rect 2506 2603 2516 2606
rect 2626 2603 2652 2606
rect 2692 2603 2709 2606
rect 2716 2603 2749 2606
rect 2754 2603 2772 2606
rect 2810 2603 2828 2606
rect 2874 2603 2901 2606
rect 1316 2593 1325 2596
rect 2220 2593 2245 2596
rect 2250 2595 2253 2603
rect 2844 2593 2853 2596
rect 2946 2595 2949 2606
rect 2956 2603 2965 2606
rect 2970 2603 3004 2606
rect 3122 2603 3180 2606
rect 3250 2603 3268 2606
rect 3282 2603 3292 2606
rect 3370 2603 3396 2606
rect 38 2567 3482 2573
rect 202 2526 205 2534
rect 260 2533 301 2536
rect 514 2533 524 2536
rect 554 2533 564 2536
rect 690 2526 693 2546
rect 116 2523 141 2526
rect 172 2523 205 2526
rect 212 2523 228 2526
rect 348 2523 357 2526
rect 404 2523 421 2526
rect 626 2523 660 2526
rect 684 2523 693 2526
rect 706 2525 709 2556
rect 730 2543 764 2546
rect 1090 2543 1116 2546
rect 1138 2543 1157 2546
rect 1268 2543 1277 2546
rect 2338 2543 2389 2546
rect 2722 2543 2741 2546
rect 2786 2543 2797 2546
rect 1154 2536 1157 2543
rect 730 2533 772 2536
rect 1076 2533 1117 2536
rect 1124 2533 1149 2536
rect 1154 2533 1164 2536
rect 1196 2533 1213 2536
rect 1218 2533 1252 2536
rect 1308 2533 1341 2536
rect 1370 2533 1380 2536
rect 1442 2533 1484 2536
rect 1522 2533 1572 2536
rect 1596 2533 1629 2536
rect 1634 2526 1637 2534
rect 1660 2533 1701 2536
rect 1706 2526 1709 2534
rect 1722 2533 1764 2536
rect 1786 2533 1820 2536
rect 1858 2533 1884 2536
rect 1978 2533 1996 2536
rect 2228 2533 2301 2536
rect 2324 2533 2341 2536
rect 1978 2526 1981 2533
rect 2378 2526 2381 2536
rect 2546 2533 2572 2536
rect 2602 2533 2644 2536
rect 2714 2533 2756 2536
rect 786 2523 796 2526
rect 828 2523 837 2526
rect 924 2523 949 2526
rect 986 2523 1028 2526
rect 1050 2523 1060 2526
rect 1132 2523 1157 2526
rect 1268 2523 1292 2526
rect 1356 2523 1365 2526
rect 1378 2523 1412 2526
rect 1516 2523 1573 2526
rect 1594 2523 1637 2526
rect 1658 2523 1709 2526
rect 1716 2523 1749 2526
rect 1780 2523 1813 2526
rect 1844 2523 1885 2526
rect 1940 2523 1981 2526
rect 2020 2523 2061 2526
rect 2092 2523 2125 2526
rect 2170 2523 2204 2526
rect 2236 2523 2277 2526
rect 2282 2523 2300 2526
rect 2332 2523 2381 2526
rect 2596 2523 2613 2526
rect 2652 2523 2677 2526
rect 2780 2523 2789 2526
rect 2794 2516 2797 2543
rect 3026 2533 3060 2536
rect 3242 2533 3276 2536
rect 604 2513 653 2516
rect 690 2513 700 2516
rect 724 2513 741 2516
rect 1660 2513 1693 2516
rect 2354 2513 2404 2516
rect 2708 2513 2741 2516
rect 2786 2513 2797 2516
rect 2818 2506 2821 2525
rect 2876 2523 2893 2526
rect 2940 2523 2957 2526
rect 3004 2523 3013 2526
rect 3068 2523 3093 2526
rect 3098 2523 3108 2526
rect 3132 2523 3165 2526
rect 3242 2516 3245 2533
rect 3410 2526 3413 2534
rect 3428 2533 3453 2536
rect 3250 2523 3284 2526
rect 3370 2523 3396 2526
rect 3410 2523 3421 2526
rect 3436 2523 3453 2526
rect 2884 2513 2893 2516
rect 3140 2513 3197 2516
rect 3242 2513 3253 2516
rect 578 2503 596 2506
rect 2346 2503 2420 2506
rect 2442 2503 2484 2506
rect 2690 2503 2700 2506
rect 2794 2503 2821 2506
rect 3194 2503 3197 2513
rect 14 2467 3506 2473
rect 1338 2433 1380 2436
rect 2562 2433 2588 2436
rect 434 2423 461 2426
rect 668 2423 677 2426
rect 1202 2423 1220 2426
rect 1244 2423 1293 2426
rect 1346 2423 1364 2426
rect 1388 2423 1397 2426
rect 2196 2423 2213 2426
rect 2538 2423 2572 2426
rect 2596 2423 2645 2426
rect 3082 2423 3117 2426
rect 3420 2423 3429 2426
rect 434 2416 437 2423
rect 3114 2416 3117 2423
rect 204 2413 245 2416
rect 340 2413 389 2416
rect 428 2413 437 2416
rect 442 2413 476 2416
rect 612 2413 637 2416
rect 642 2413 652 2416
rect 794 2413 828 2416
rect 860 2413 869 2416
rect 972 2413 997 2416
rect 1050 2413 1076 2416
rect 1138 2413 1180 2416
rect 1186 2413 1196 2416
rect 1258 2413 1308 2416
rect 1394 2413 1444 2416
rect 1532 2413 1565 2416
rect 1618 2413 1628 2416
rect 1708 2413 1741 2416
rect 1772 2413 1813 2416
rect 1844 2413 1869 2416
rect 196 2403 245 2406
rect 394 2403 404 2406
rect 458 2403 468 2406
rect 546 2403 572 2406
rect 596 2403 604 2406
rect 618 2403 644 2406
rect 668 2403 693 2406
rect 698 2403 716 2406
rect 746 2403 764 2406
rect 780 2403 789 2406
rect 802 2403 836 2406
rect 858 2403 868 2406
rect 1042 2403 1068 2406
rect 1124 2403 1157 2406
rect 1274 2403 1300 2406
rect 1468 2403 1493 2406
rect 1572 2403 1613 2406
rect 1658 2403 1700 2406
rect 1738 2403 1748 2406
rect 1836 2403 1853 2406
rect 1866 2403 1869 2413
rect 1930 2413 1956 2416
rect 2028 2413 2069 2416
rect 2108 2413 2117 2416
rect 2122 2413 2180 2416
rect 2236 2413 2261 2416
rect 2324 2413 2341 2416
rect 2378 2413 2412 2416
rect 2738 2413 2764 2416
rect 2788 2413 2797 2416
rect 2804 2413 2829 2416
rect 2884 2413 2909 2416
rect 2914 2413 2924 2416
rect 2930 2413 2948 2416
rect 2970 2413 2996 2416
rect 3068 2413 3109 2416
rect 3114 2413 3132 2416
rect 3178 2413 3237 2416
rect 3290 2413 3308 2416
rect 3330 2413 3373 2416
rect 3380 2413 3397 2416
rect 1930 2406 1933 2413
rect 2066 2406 2069 2413
rect 3106 2406 3109 2413
rect 1884 2403 1933 2406
rect 1980 2403 1997 2406
rect 2002 2403 2020 2406
rect 2066 2403 2084 2406
rect 2300 2403 2316 2406
rect 2362 2403 2404 2406
rect 2436 2403 2453 2406
rect 2498 2403 2516 2406
rect 2660 2403 2676 2406
rect 2700 2403 2757 2406
rect 2810 2403 2876 2406
rect 2954 2403 3004 2406
rect 3026 2403 3060 2406
rect 3106 2403 3140 2406
rect 3156 2403 3197 2406
rect 3362 2403 3372 2406
rect 3394 2405 3397 2413
rect 1538 2393 1564 2396
rect 1818 2393 1828 2396
rect 1850 2393 1876 2396
rect 2242 2393 2292 2396
rect 2532 2393 2541 2396
rect 2626 2393 2652 2396
rect 38 2367 3482 2373
rect 2354 2353 2389 2356
rect 1202 2343 1236 2346
rect 1948 2343 1965 2346
rect 2354 2336 2357 2353
rect 2386 2343 2396 2346
rect 2642 2336 2645 2356
rect 2786 2343 2820 2346
rect 186 2326 189 2335
rect 228 2333 245 2336
rect 378 2326 381 2335
rect 436 2333 461 2336
rect 698 2333 740 2336
rect 764 2333 773 2336
rect 858 2333 868 2336
rect 1010 2333 1044 2336
rect 1100 2333 1141 2336
rect 1146 2333 1156 2336
rect 1244 2333 1269 2336
rect 1378 2333 1388 2336
rect 1146 2326 1149 2333
rect 1426 2326 1429 2335
rect 1506 2333 1556 2336
rect 1570 2333 1604 2336
rect 1642 2333 1700 2336
rect 1724 2333 1773 2336
rect 1812 2333 1861 2336
rect 1866 2326 1869 2335
rect 1882 2333 1932 2336
rect 2004 2333 2053 2336
rect 2058 2333 2068 2336
rect 2092 2333 2101 2336
rect 2186 2333 2204 2336
rect 2228 2333 2237 2336
rect 2298 2333 2308 2336
rect 2324 2333 2357 2336
rect 2362 2333 2404 2336
rect 2410 2333 2437 2336
rect 2538 2333 2556 2336
rect 2570 2333 2612 2336
rect 2634 2333 2645 2336
rect 2674 2333 2692 2336
rect 2828 2333 2876 2336
rect 2900 2333 2941 2336
rect 3090 2333 3148 2336
rect 3172 2333 3197 2336
rect 3226 2333 3260 2336
rect 3290 2333 3300 2336
rect 3338 2333 3404 2336
rect 116 2323 141 2326
rect 172 2323 189 2326
rect 196 2323 212 2326
rect 292 2323 317 2326
rect 348 2323 381 2326
rect 388 2323 404 2326
rect 508 2323 517 2326
rect 570 2323 580 2326
rect 612 2323 621 2326
rect 658 2323 668 2326
rect 762 2323 772 2326
rect 810 2323 828 2326
rect 860 2323 869 2326
rect 948 2323 973 2326
rect 1026 2323 1052 2326
rect 1074 2323 1084 2326
rect 1130 2323 1149 2326
rect 1180 2323 1189 2326
rect 1266 2323 1276 2326
rect 1346 2323 1364 2326
rect 1396 2323 1429 2326
rect 1450 2323 1484 2326
rect 1500 2323 1549 2326
rect 1564 2323 1605 2326
rect 1650 2323 1708 2326
rect 1722 2323 1796 2326
rect 1850 2323 1869 2326
rect 1876 2323 1901 2326
rect 1914 2323 1924 2326
rect 2050 2323 2053 2333
rect 2090 2323 2148 2326
rect 2154 2323 2212 2326
rect 2282 2323 2300 2326
rect 2410 2325 2413 2333
rect 2418 2323 2452 2326
rect 2564 2323 2597 2326
rect 2634 2325 2637 2333
rect 3290 2326 3293 2333
rect 2642 2323 2684 2326
rect 2836 2323 2877 2326
rect 2964 2323 3005 2326
rect 3012 2323 3029 2326
rect 3034 2323 3060 2326
rect 3092 2323 3141 2326
rect 3202 2323 3261 2326
rect 3268 2323 3293 2326
rect 3308 2323 3317 2326
rect 3332 2323 3389 2326
rect 3428 2323 3437 2326
rect 228 2313 253 2316
rect 1100 2313 1109 2316
rect 1724 2313 1749 2316
rect 1812 2313 1837 2316
rect 2228 2313 2293 2316
rect 2780 2313 2789 2316
rect 3220 2313 3229 2316
rect 14 2267 3506 2273
rect 650 2233 701 2236
rect 2906 2233 2956 2236
rect 3090 2233 3148 2236
rect 650 2223 692 2226
rect 172 2213 213 2216
rect 220 2213 236 2216
rect 276 2213 285 2216
rect 404 2213 437 2216
rect 210 2205 213 2213
rect 442 2206 445 2214
rect 522 2213 572 2216
rect 650 2213 653 2223
rect 698 2215 701 2233
rect 1204 2223 1213 2226
rect 1346 2223 1364 2226
rect 1388 2223 1397 2226
rect 1458 2216 1461 2225
rect 1564 2223 1573 2226
rect 1660 2223 1701 2226
rect 1740 2223 1773 2226
rect 1812 2223 1861 2226
rect 746 2213 772 2216
rect 804 2213 813 2216
rect 892 2213 917 2216
rect 954 2213 996 2216
rect 1042 2213 1100 2216
rect 1138 2213 1188 2216
rect 1234 2206 1237 2214
rect 1260 2213 1309 2216
rect 1426 2213 1444 2216
rect 1458 2213 1469 2216
rect 1484 2213 1533 2216
rect 1556 2213 1565 2216
rect 1466 2206 1469 2213
rect 268 2203 301 2206
rect 410 2203 445 2206
rect 610 2203 620 2206
rect 636 2203 685 2206
rect 722 2203 732 2206
rect 1044 2203 1077 2206
rect 1082 2203 1092 2206
rect 1204 2203 1237 2206
rect 1266 2203 1308 2206
rect 1332 2203 1341 2206
rect 1418 2203 1436 2206
rect 1466 2203 1476 2206
rect 1482 2203 1548 2206
rect 1570 2205 1573 2223
rect 2250 2216 2253 2225
rect 2708 2223 2717 2226
rect 2914 2223 2940 2226
rect 3090 2223 3132 2226
rect 3156 2223 3165 2226
rect 1580 2213 1637 2216
rect 1634 2205 1637 2213
rect 1658 2213 1717 2216
rect 1810 2213 1868 2216
rect 1956 2213 1973 2216
rect 2060 2213 2093 2216
rect 2122 2213 2132 2216
rect 2202 2213 2236 2216
rect 2250 2213 2300 2216
rect 2410 2213 2444 2216
rect 2490 2213 2540 2216
rect 2572 2213 2621 2216
rect 2674 2213 2700 2216
rect 2738 2213 2772 2216
rect 2820 2213 2853 2216
rect 2900 2213 2933 2216
rect 3028 2213 3061 2216
rect 1658 2205 1661 2213
rect 2090 2206 2093 2213
rect 1666 2203 1716 2206
rect 1740 2203 1773 2206
rect 1890 2203 1932 2206
rect 1948 2203 1965 2206
rect 2010 2203 2036 2206
rect 2090 2203 2140 2206
rect 2156 2203 2221 2206
rect 2252 2203 2277 2206
rect 2298 2203 2308 2206
rect 2324 2203 2341 2206
rect 2354 2203 2380 2206
rect 2468 2203 2548 2206
rect 2570 2203 2636 2206
rect 2660 2203 2685 2206
rect 2730 2203 2764 2206
rect 2788 2203 2797 2206
rect 2866 2203 2876 2206
rect 2970 2203 3004 2206
rect 3058 2205 3061 2213
rect 3162 2206 3165 2223
rect 3306 2216 3309 2225
rect 3170 2213 3196 2216
rect 3220 2213 3261 2216
rect 3266 2213 3284 2216
rect 3306 2213 3317 2216
rect 3324 2213 3341 2216
rect 3346 2213 3364 2216
rect 3266 2206 3269 2213
rect 3084 2203 3117 2206
rect 3162 2203 3204 2206
rect 3258 2203 3269 2206
rect 3330 2203 3372 2206
rect 3220 2193 3229 2196
rect 38 2167 3482 2173
rect 1626 2143 1660 2146
rect 2058 2143 2068 2146
rect 2514 2143 2533 2146
rect 3034 2143 3068 2146
rect 3154 2143 3181 2146
rect 3212 2143 3229 2146
rect 3154 2136 3157 2143
rect 218 2126 221 2135
rect 276 2133 317 2136
rect 468 2133 477 2136
rect 522 2133 532 2136
rect 642 2133 692 2136
rect 818 2133 828 2136
rect 1074 2133 1084 2136
rect 1108 2133 1125 2136
rect 1170 2133 1196 2136
rect 1212 2133 1229 2136
rect 124 2123 149 2126
rect 180 2123 221 2126
rect 228 2123 244 2126
rect 412 2123 437 2126
rect 506 2123 549 2126
rect 562 2123 580 2126
rect 690 2123 700 2126
rect 714 2123 725 2126
rect 754 2123 788 2126
rect 916 2123 941 2126
rect 1066 2123 1092 2126
rect 1140 2123 1149 2126
rect 1170 2123 1173 2133
rect 1220 2123 1237 2126
rect 1276 2123 1293 2126
rect 714 2115 717 2123
rect 1298 2116 1301 2135
rect 1346 2133 1364 2136
rect 1458 2133 1476 2136
rect 1538 2133 1572 2136
rect 1594 2133 1604 2136
rect 1634 2126 1637 2136
rect 1668 2133 1693 2136
rect 1700 2133 1717 2136
rect 1722 2133 1772 2136
rect 1796 2133 1837 2136
rect 1860 2133 1869 2136
rect 1986 2133 2028 2136
rect 2034 2133 2076 2136
rect 2082 2133 2133 2136
rect 2172 2133 2221 2136
rect 2236 2133 2269 2136
rect 2346 2133 2364 2136
rect 2402 2133 2452 2136
rect 2466 2133 2476 2136
rect 2500 2133 2509 2136
rect 2580 2133 2597 2136
rect 2602 2133 2612 2136
rect 2634 2133 2652 2136
rect 2802 2133 2812 2136
rect 2836 2133 2853 2136
rect 2906 2133 2924 2136
rect 2938 2133 2956 2136
rect 2994 2133 3004 2136
rect 3076 2133 3116 2136
rect 3140 2133 3157 2136
rect 3258 2133 3308 2136
rect 3362 2133 3404 2136
rect 1372 2123 1389 2126
rect 1394 2123 1412 2126
rect 1484 2123 1501 2126
rect 1148 2113 1181 2116
rect 1284 2113 1301 2116
rect 1394 2113 1397 2123
rect 1490 2113 1508 2116
rect 1514 2106 1517 2125
rect 1580 2123 1605 2126
rect 1612 2123 1637 2126
rect 1676 2123 1685 2126
rect 1730 2123 1780 2126
rect 2036 2123 2045 2126
rect 2082 2125 2085 2133
rect 2266 2127 2269 2133
rect 2090 2123 2148 2126
rect 2266 2124 2284 2127
rect 2338 2123 2356 2126
rect 2460 2123 2484 2126
rect 2498 2123 2556 2126
rect 2602 2123 2620 2126
rect 2626 2123 2660 2126
rect 2682 2123 2700 2126
rect 2714 2123 2748 2126
rect 2778 2123 2820 2126
rect 1532 2113 1573 2116
rect 1796 2113 1837 2116
rect 1964 2113 1973 2116
rect 2276 2113 2285 2116
rect 2300 2113 2317 2116
rect 2500 2113 2517 2116
rect 1506 2103 1517 2106
rect 1946 2103 1956 2106
rect 2274 2103 2292 2106
rect 2602 2093 2605 2123
rect 2714 2103 2717 2123
rect 2764 2113 2773 2116
rect 2850 2106 2853 2133
rect 3362 2126 3365 2133
rect 2932 2123 2957 2126
rect 2978 2123 2996 2126
rect 3084 2123 3101 2126
rect 3106 2123 3124 2126
rect 3162 2123 3188 2126
rect 3212 2123 3245 2126
rect 3252 2123 3285 2126
rect 3316 2123 3325 2126
rect 3340 2123 3365 2126
rect 3386 2123 3396 2126
rect 3106 2116 3109 2123
rect 3090 2113 3109 2116
rect 2850 2103 2892 2106
rect 14 2067 3506 2073
rect 1346 2053 1389 2056
rect 602 2026 605 2036
rect 588 2023 605 2026
rect 754 2033 780 2036
rect 754 2016 757 2033
rect 764 2023 773 2026
rect 1052 2023 1069 2026
rect 1234 2016 1237 2036
rect 1714 2033 1764 2036
rect 2050 2033 2068 2036
rect 2626 2033 2661 2036
rect 3130 2033 3188 2036
rect 1420 2023 1429 2026
rect 1634 2016 1637 2026
rect 1722 2023 1748 2026
rect 1772 2023 1821 2026
rect 1844 2023 1853 2026
rect 1996 2023 2005 2026
rect 2010 2023 2052 2026
rect 2076 2023 2085 2026
rect 2282 2023 2301 2026
rect 2386 2023 2444 2026
rect 2554 2023 2589 2026
rect 2002 2016 2005 2023
rect 124 2013 149 2016
rect 180 2013 221 2016
rect 228 2013 244 2016
rect 258 2013 269 2016
rect 404 2013 437 2016
rect 218 2005 221 2013
rect 266 1995 269 2013
rect 442 2006 445 2014
rect 516 2013 572 2016
rect 602 2013 620 2016
rect 658 2013 676 2016
rect 740 2013 757 2016
rect 836 2013 845 2016
rect 852 2013 885 2016
rect 932 2013 957 2016
rect 1002 2013 1036 2016
rect 418 2003 445 2006
rect 474 2003 492 2006
rect 530 2003 564 2006
rect 594 2003 612 2006
rect 642 2003 668 2006
rect 692 2003 701 2006
rect 706 2003 716 2006
rect 794 2003 812 2006
rect 834 2003 844 2006
rect 1010 2003 1028 2006
rect 1090 1996 1093 2014
rect 1116 2013 1165 2016
rect 1196 2013 1237 2016
rect 1282 2013 1309 2016
rect 1098 2003 1133 2006
rect 1138 2003 1164 2006
rect 1210 2003 1252 2006
rect 1268 2003 1293 2006
rect 1306 2005 1309 2013
rect 1346 2013 1404 2016
rect 1442 2013 1468 2016
rect 1506 2013 1524 2016
rect 1562 2013 1604 2016
rect 1634 2013 1668 2016
rect 1836 2013 1893 2016
rect 1970 2013 1980 2016
rect 2002 2013 2029 2016
rect 2042 2013 2060 2016
rect 2148 2013 2157 2016
rect 2164 2013 2189 2016
rect 1346 2003 1349 2013
rect 2042 2006 2045 2013
rect 2234 2006 2237 2014
rect 2268 2013 2309 2016
rect 2330 2013 2348 2016
rect 2380 2013 2437 2016
rect 2482 2013 2516 2016
rect 2554 2006 2557 2023
rect 2562 2013 2596 2016
rect 2658 2015 2661 2033
rect 2676 2023 2693 2026
rect 2716 2023 2757 2026
rect 3116 2023 3172 2026
rect 3268 2023 3285 2026
rect 2682 2013 2708 2016
rect 2780 2013 2789 2016
rect 2804 2013 2821 2016
rect 2858 2013 2868 2016
rect 2900 2013 2956 2016
rect 2988 2013 2997 2016
rect 3060 2013 3077 2016
rect 3082 2013 3100 2016
rect 3114 2013 3165 2016
rect 3260 2013 3293 2016
rect 3332 2013 3373 2016
rect 3290 2006 3293 2013
rect 1498 2003 1532 2006
rect 1570 2003 1596 2006
rect 1634 2003 1660 2006
rect 1692 2003 1725 2006
rect 1786 2003 1828 2006
rect 1916 2003 1965 2006
rect 1996 2003 2045 2006
rect 2090 2003 2140 2006
rect 2186 2003 2237 2006
rect 2260 2003 2285 2006
rect 2346 2003 2356 2006
rect 2540 2003 2557 2006
rect 2570 2003 2588 2006
rect 2682 2003 2700 2006
rect 2714 2003 2772 2006
rect 2796 2003 2853 2006
rect 2906 2003 2964 2006
rect 2980 2003 3045 2006
rect 3052 2003 3092 2006
rect 3116 2003 3165 2006
rect 3242 2003 3252 2006
rect 3290 2003 3308 2006
rect 3324 2003 3341 2006
rect 3362 2003 3372 2006
rect 3396 2003 3405 2006
rect 1130 1996 1133 2003
rect 2282 1996 2285 2003
rect 1090 1993 1100 1996
rect 1130 1993 1149 1996
rect 2282 1993 2341 1996
rect 2722 1993 2764 1996
rect 2850 1983 2853 2003
rect 2994 1993 3044 1996
rect 3162 1993 3165 2003
rect 3402 1995 3405 2003
rect 38 1967 3482 1973
rect 610 1943 620 1946
rect 1210 1943 1252 1946
rect 1290 1943 1348 1946
rect 210 1926 213 1934
rect 268 1933 285 1936
rect 410 1933 428 1936
rect 628 1933 645 1936
rect 650 1933 660 1936
rect 682 1933 724 1936
rect 746 1933 764 1936
rect 836 1933 852 1936
rect 868 1933 893 1936
rect 1116 1933 1165 1936
rect 1170 1926 1173 1934
rect 1266 1933 1276 1936
rect 1338 1933 1356 1936
rect 116 1923 141 1926
rect 172 1923 213 1926
rect 220 1923 236 1926
rect 396 1923 405 1926
rect 458 1923 485 1926
rect 540 1923 557 1926
rect 596 1923 621 1926
rect 636 1923 645 1926
rect 684 1923 709 1926
rect 876 1923 901 1926
rect 940 1923 965 1926
rect 996 1923 1005 1926
rect 1018 1923 1052 1926
rect 1122 1923 1173 1926
rect 1180 1923 1197 1926
rect 1204 1923 1245 1926
rect 1268 1923 1277 1926
rect 1364 1923 1373 1926
rect 1380 1923 1445 1926
rect 1490 1923 1493 1946
rect 2114 1943 2125 1946
rect 1556 1933 1581 1936
rect 1602 1933 1628 1936
rect 1650 1933 1700 1936
rect 1714 1933 1764 1936
rect 1794 1933 1836 1936
rect 1860 1933 1925 1936
rect 1932 1933 1956 1936
rect 2018 1933 2036 1936
rect 2052 1933 2117 1936
rect 2018 1926 2021 1933
rect 2122 1926 2125 1943
rect 2130 1933 2140 1936
rect 2156 1933 2205 1936
rect 2242 1933 2252 1936
rect 2314 1933 2324 1936
rect 2348 1933 2357 1936
rect 2394 1926 2397 1934
rect 2498 1933 2509 1936
rect 2532 1933 2565 1936
rect 2682 1933 2692 1936
rect 2850 1933 2876 1936
rect 2900 1933 2941 1936
rect 3034 1933 3076 1936
rect 3098 1933 3148 1936
rect 3194 1933 3204 1936
rect 3290 1933 3300 1936
rect 3338 1933 3404 1936
rect 1554 1923 1629 1926
rect 1636 1923 1701 1926
rect 1708 1923 1757 1926
rect 1788 1923 1837 1926
rect 1964 1923 2021 1926
rect 2060 1923 2101 1926
rect 2122 1923 2132 1926
rect 2260 1923 2332 1926
rect 2346 1923 2397 1926
rect 2418 1923 2436 1926
rect 482 1916 485 1923
rect 2498 1916 2501 1933
rect 2682 1923 2700 1926
rect 2714 1923 2748 1926
rect 2754 1923 2764 1926
rect 2978 1923 3020 1926
rect 3114 1923 3140 1926
rect 3164 1923 3205 1926
rect 3212 1923 3229 1926
rect 3308 1923 3325 1926
rect 3332 1923 3357 1926
rect 3386 1923 3396 1926
rect 2730 1916 2733 1923
rect 482 1913 500 1916
rect 1484 1913 1525 1916
rect 1716 1913 1749 1916
rect 1860 1913 1909 1916
rect 2268 1913 2317 1916
rect 2444 1913 2501 1916
rect 2546 1913 2581 1916
rect 2602 1913 2644 1916
rect 2708 1913 2733 1916
rect 2772 1913 2820 1916
rect 2844 1913 2853 1916
rect 2900 1913 2948 1916
rect 3028 1913 3061 1916
rect 3220 1913 3229 1916
rect 498 1903 516 1906
rect 2546 1903 2588 1906
rect 2642 1903 2660 1906
rect 2794 1903 2836 1906
rect 2906 1903 2964 1906
rect 2610 1883 2637 1886
rect 14 1867 3506 1873
rect 2186 1853 2229 1856
rect 498 1833 516 1836
rect 1290 1833 1309 1836
rect 3394 1833 3421 1836
rect 372 1823 397 1826
rect 524 1823 549 1826
rect 1180 1823 1205 1826
rect 1268 1823 1285 1826
rect 1290 1816 1293 1833
rect 164 1813 205 1816
rect 244 1813 261 1816
rect 300 1813 333 1816
rect 340 1813 356 1816
rect 386 1813 404 1816
rect 436 1813 453 1816
rect 538 1813 564 1816
rect 156 1803 197 1806
rect 330 1805 333 1813
rect 586 1806 589 1814
rect 618 1806 621 1814
rect 732 1813 757 1816
rect 868 1813 892 1816
rect 924 1813 941 1816
rect 980 1813 1005 1816
rect 1036 1813 1045 1816
rect 1050 1813 1076 1816
rect 1090 1813 1101 1816
rect 1132 1813 1149 1816
rect 1212 1813 1229 1816
rect 1234 1813 1260 1816
rect 1266 1813 1293 1816
rect 1306 1815 1309 1833
rect 1324 1823 1333 1826
rect 1660 1823 1669 1826
rect 1860 1823 1909 1826
rect 2018 1823 2029 1826
rect 2084 1823 2141 1826
rect 554 1803 572 1806
rect 586 1803 597 1806
rect 618 1803 668 1806
rect 698 1803 708 1806
rect 724 1803 733 1806
rect 1058 1803 1068 1806
rect 1098 1805 1101 1813
rect 1330 1806 1333 1823
rect 1378 1813 1395 1816
rect 1524 1813 1565 1816
rect 1602 1813 1644 1816
rect 1716 1813 1765 1816
rect 1780 1813 1837 1816
rect 1948 1813 1965 1816
rect 1130 1803 1156 1806
rect 1180 1803 1197 1806
rect 1330 1803 1340 1806
rect 1370 1803 1388 1806
rect 1468 1803 1501 1806
rect 1522 1803 1564 1806
rect 1626 1803 1636 1806
rect 1660 1803 1701 1806
rect 1834 1805 1837 1813
rect 2018 1806 2021 1823
rect 2378 1816 2381 1824
rect 2580 1823 2605 1826
rect 2930 1823 2964 1826
rect 3092 1823 3101 1826
rect 3370 1823 3412 1826
rect 3098 1816 3101 1823
rect 2026 1813 2068 1816
rect 2180 1813 2197 1816
rect 2252 1813 2293 1816
rect 2308 1813 2349 1816
rect 2378 1813 2397 1816
rect 2452 1813 2493 1816
rect 1860 1803 1932 1806
rect 2012 1803 2021 1806
rect 2034 1803 2060 1806
rect 2084 1803 2093 1806
rect 2114 1803 2156 1806
rect 2172 1803 2205 1806
rect 620 1793 629 1796
rect 1442 1793 1460 1796
rect 1524 1793 1557 1796
rect 1874 1793 1924 1796
rect 2290 1795 2293 1813
rect 2394 1796 2397 1813
rect 2498 1806 2501 1815
rect 2538 1813 2572 1816
rect 2578 1813 2628 1816
rect 2666 1813 2700 1816
rect 2714 1813 2733 1816
rect 2740 1813 2757 1816
rect 2868 1813 2893 1816
rect 3004 1813 3013 1816
rect 3050 1813 3076 1816
rect 3098 1813 3108 1816
rect 3180 1813 3197 1816
rect 3221 1813 3229 1816
rect 3234 1813 3277 1816
rect 3292 1813 3325 1816
rect 3364 1813 3405 1816
rect 3418 1815 3421 1833
rect 3436 1823 3493 1826
rect 2402 1803 2444 1806
rect 2466 1803 2501 1806
rect 2530 1803 2564 1806
rect 2610 1803 2636 1806
rect 2674 1803 2692 1806
rect 2714 1803 2732 1806
rect 2780 1803 2837 1806
rect 2866 1803 2892 1806
rect 2916 1803 2941 1806
rect 3124 1803 3165 1806
rect 3172 1803 3181 1806
rect 3258 1803 3284 1806
rect 3314 1803 3340 1806
rect 2394 1793 2405 1796
rect 2938 1793 2941 1803
rect 3130 1793 3164 1796
rect 2602 1783 2621 1786
rect 38 1767 3482 1773
rect 3490 1756 3493 1823
rect 282 1743 308 1746
rect 474 1743 500 1746
rect 210 1726 213 1734
rect 356 1733 381 1736
rect 538 1733 548 1736
rect 650 1733 660 1736
rect 676 1733 693 1736
rect 818 1733 829 1736
rect 860 1733 876 1736
rect 898 1733 908 1736
rect 826 1726 829 1733
rect 922 1726 925 1746
rect 1410 1743 1444 1746
rect 1050 1733 1068 1736
rect 1108 1733 1125 1736
rect 1146 1733 1196 1736
rect 1226 1733 1236 1736
rect 1482 1733 1492 1736
rect 1530 1733 1556 1736
rect 1594 1726 1597 1756
rect 3434 1753 3493 1756
rect 1706 1736 1709 1746
rect 1650 1733 1684 1736
rect 1706 1733 1732 1736
rect 1754 1733 1804 1736
rect 1828 1733 1869 1736
rect 1922 1726 1925 1745
rect 1946 1743 1973 1746
rect 1970 1736 1973 1743
rect 2178 1743 2205 1746
rect 2210 1743 2228 1746
rect 2914 1743 2924 1746
rect 2178 1736 2181 1743
rect 1932 1733 1965 1736
rect 1970 1733 1988 1736
rect 2012 1733 2029 1736
rect 2034 1733 2068 1736
rect 2098 1733 2148 1736
rect 2164 1733 2181 1736
rect 2194 1733 2236 1736
rect 2258 1733 2284 1736
rect 2402 1733 2420 1736
rect 2436 1733 2485 1736
rect 2514 1733 2556 1736
rect 2618 1733 2652 1736
rect 2842 1733 2876 1736
rect 2932 1733 2949 1736
rect 2098 1726 2101 1733
rect 124 1723 149 1726
rect 180 1723 213 1726
rect 220 1723 236 1726
rect 364 1723 405 1726
rect 540 1723 556 1726
rect 596 1723 613 1726
rect 684 1723 717 1726
rect 812 1723 821 1726
rect 826 1723 844 1726
rect 900 1723 909 1726
rect 916 1723 925 1726
rect 980 1723 1005 1726
rect 1036 1723 1045 1726
rect 1066 1723 1076 1726
rect 1082 1723 1092 1726
rect 1106 1723 1133 1726
rect 1148 1723 1197 1726
rect 1354 1723 1380 1726
rect 1460 1723 1493 1726
rect 1546 1723 1564 1726
rect 1570 1723 1597 1726
rect 444 1713 453 1716
rect 468 1713 485 1716
rect 1252 1713 1285 1716
rect 1594 1713 1612 1716
rect 1618 1706 1621 1725
rect 1740 1723 1805 1726
rect 1884 1723 1925 1726
rect 1940 1723 1989 1726
rect 2092 1723 2101 1726
rect 2122 1723 2140 1726
rect 2292 1723 2356 1726
rect 2378 1723 2412 1726
rect 2444 1723 2469 1726
rect 2516 1723 2549 1726
rect 2554 1723 2564 1726
rect 1636 1713 1669 1716
rect 1748 1713 1765 1716
rect 1828 1713 1869 1716
rect 1892 1713 1901 1716
rect 2300 1713 2325 1716
rect 2378 1713 2381 1723
rect 2578 1706 2581 1725
rect 2690 1723 2700 1726
rect 2722 1723 2772 1726
rect 2778 1723 2788 1726
rect 2946 1716 2949 1733
rect 3010 1733 3044 1736
rect 3060 1733 3101 1736
rect 3204 1733 3229 1736
rect 3234 1733 3260 1736
rect 3282 1733 3300 1736
rect 3394 1733 3413 1736
rect 3010 1716 3013 1733
rect 2676 1713 2685 1716
rect 2946 1713 2956 1716
rect 2980 1713 3013 1716
rect 3018 1723 3036 1726
rect 3068 1723 3085 1726
rect 3116 1723 3141 1726
rect 3018 1706 3021 1723
rect 3124 1713 3157 1716
rect 3226 1713 3229 1733
rect 3268 1723 3301 1726
rect 3308 1723 3325 1726
rect 3338 1723 3364 1726
rect 3394 1725 3397 1733
rect 3402 1723 3428 1726
rect 3276 1713 3285 1716
rect 442 1703 460 1706
rect 1154 1703 1197 1706
rect 1610 1703 1621 1706
rect 2570 1703 2581 1706
rect 2954 1703 2972 1706
rect 2986 1703 3021 1706
rect 14 1667 3506 1673
rect 3066 1643 3093 1646
rect 3226 1643 3245 1646
rect 506 1633 532 1636
rect 1266 1633 1300 1636
rect 1970 1633 2004 1636
rect 2466 1633 2508 1636
rect 3114 1626 3117 1636
rect 3130 1633 3140 1636
rect 356 1623 365 1626
rect 498 1623 516 1626
rect 1028 1623 1061 1626
rect 1250 1623 1284 1626
rect 1548 1623 1557 1626
rect 1804 1623 1845 1626
rect 1978 1623 1988 1626
rect 2340 1623 2373 1626
rect 2482 1623 2492 1626
rect 2724 1623 2741 1626
rect 2948 1623 2957 1626
rect 3114 1623 3124 1626
rect 3148 1623 3189 1626
rect 1978 1616 1981 1623
rect 228 1613 253 1616
rect 284 1613 317 1616
rect 324 1613 340 1616
rect 578 1613 588 1616
rect 644 1613 653 1616
rect 666 1613 676 1616
rect 956 1613 981 1616
rect 986 1613 996 1616
rect 1002 1613 1012 1616
rect 1066 1613 1076 1616
rect 1116 1613 1125 1616
rect 1138 1613 1156 1616
rect 1338 1613 1405 1616
rect 1458 1613 1468 1616
rect 1492 1613 1532 1616
rect 1546 1613 1588 1616
rect 1668 1613 1685 1616
rect 1692 1613 1741 1616
rect 1756 1613 1781 1616
rect 1858 1613 1868 1616
rect 1964 1613 1981 1616
rect 2076 1613 2085 1616
rect 2090 1613 2108 1616
rect 2140 1613 2173 1616
rect 2300 1613 2324 1616
rect 2452 1613 2469 1616
rect 2596 1613 2637 1616
rect 2652 1613 2661 1616
rect 2684 1613 2701 1616
rect 2722 1613 2772 1616
rect 2804 1613 2829 1616
rect 2844 1613 2877 1616
rect 2978 1613 2996 1616
rect 3020 1613 3045 1616
rect 3052 1613 3069 1616
rect 3074 1613 3108 1616
rect 314 1605 317 1613
rect 410 1603 444 1606
rect 484 1603 509 1606
rect 570 1603 580 1606
rect 636 1603 677 1606
rect 916 1603 925 1606
rect 954 1603 988 1606
rect 1042 1603 1068 1606
rect 1092 1603 1101 1606
rect 1108 1603 1125 1606
rect 1154 1603 1164 1606
rect 1180 1603 1205 1606
rect 1210 1603 1220 1606
rect 1330 1603 1364 1606
rect 1402 1605 1405 1613
rect 2090 1606 2093 1613
rect 1436 1603 1461 1606
rect 1490 1603 1524 1606
rect 1548 1603 1573 1606
rect 1626 1603 1660 1606
rect 1706 1603 1748 1606
rect 1770 1603 1780 1606
rect 1804 1603 1869 1606
rect 1922 1603 1940 1606
rect 2026 1603 2060 1606
rect 2082 1603 2093 1606
rect 2098 1603 2116 1606
rect 2132 1603 2188 1606
rect 2250 1603 2292 1606
rect 2386 1603 2396 1606
rect 2572 1603 2581 1606
rect 2594 1603 2644 1606
rect 2676 1603 2700 1606
rect 2724 1603 2757 1606
rect 2796 1603 2805 1606
rect 2018 1593 2052 1596
rect 2578 1595 2581 1603
rect 2658 1593 2668 1596
rect 2754 1583 2757 1603
rect 2826 1595 2829 1613
rect 3186 1606 3189 1623
rect 3226 1616 3229 1643
rect 3221 1613 3229 1616
rect 3234 1606 3237 1636
rect 3282 1623 3293 1626
rect 3290 1616 3293 1623
rect 3242 1613 3285 1616
rect 3290 1613 3308 1616
rect 3314 1613 3340 1616
rect 2836 1603 2884 1606
rect 2914 1603 2924 1606
rect 2962 1603 3004 1606
rect 3186 1603 3204 1606
rect 3234 1603 3252 1606
rect 3322 1603 3348 1606
rect 3402 1603 3412 1606
rect 3220 1593 3229 1596
rect 38 1567 3482 1573
rect 1170 1553 1181 1556
rect 178 1543 196 1546
rect 370 1536 373 1546
rect 122 1533 132 1536
rect 204 1533 253 1536
rect 354 1533 389 1536
rect 412 1533 421 1536
rect 140 1523 156 1526
rect 212 1523 245 1526
rect 348 1523 381 1526
rect 386 1525 389 1533
rect 554 1526 557 1534
rect 586 1533 604 1536
rect 634 1526 637 1534
rect 730 1533 740 1536
rect 1002 1533 1028 1536
rect 1170 1526 1173 1553
rect 2098 1546 2101 1556
rect 1212 1543 1237 1546
rect 1442 1543 1476 1546
rect 1802 1543 1812 1546
rect 2090 1543 2101 1546
rect 1178 1533 1196 1536
rect 1234 1533 1252 1536
rect 1276 1533 1293 1536
rect 1322 1533 1364 1536
rect 1386 1526 1389 1534
rect 1402 1533 1420 1536
rect 1484 1533 1517 1536
rect 1562 1533 1588 1536
rect 1610 1533 1652 1536
rect 1674 1533 1684 1536
rect 1698 1533 1756 1536
rect 1780 1533 1820 1536
rect 1930 1533 1940 1536
rect 1986 1533 2004 1536
rect 506 1523 557 1526
rect 626 1523 637 1526
rect 738 1523 748 1526
rect 802 1523 812 1526
rect 932 1523 957 1526
rect 994 1523 1036 1526
rect 1148 1523 1173 1526
rect 1212 1523 1253 1526
rect 1298 1523 1316 1526
rect 1346 1523 1372 1526
rect 1386 1523 1421 1526
rect 1428 1523 1477 1526
rect 1596 1523 1653 1526
rect 1660 1523 1685 1526
rect 1692 1523 1757 1526
rect 1836 1523 1877 1526
rect 1906 1523 1948 1526
rect 1962 1523 1996 1526
rect 2028 1523 2037 1526
rect 2090 1525 2093 1543
rect 2146 1526 2149 1546
rect 2740 1543 2757 1546
rect 2154 1533 2163 1536
rect 2188 1533 2205 1536
rect 2268 1533 2301 1536
rect 2330 1533 2365 1536
rect 2298 1526 2301 1533
rect 2098 1523 2132 1526
rect 2146 1523 2172 1526
rect 2186 1523 2243 1526
rect 2298 1523 2357 1526
rect 2362 1525 2365 1533
rect 2394 1533 2405 1536
rect 2474 1533 2508 1536
rect 2554 1533 2572 1536
rect 2594 1533 2604 1536
rect 2826 1533 2836 1536
rect 2858 1533 2900 1536
rect 2922 1533 2957 1536
rect 3106 1533 3132 1536
rect 3146 1533 3180 1536
rect 3234 1533 3252 1536
rect 3282 1533 3324 1536
rect 2394 1526 2397 1533
rect 2394 1525 2429 1526
rect 2396 1523 2429 1525
rect 2490 1523 2500 1526
rect 2546 1523 2580 1526
rect 2612 1523 2621 1526
rect 2634 1523 2684 1526
rect 2740 1523 2757 1526
rect 2834 1523 2844 1526
rect 2850 1523 2892 1526
rect 2922 1525 2925 1533
rect 3002 1526 3020 1527
rect 2954 1523 2972 1526
rect 2994 1524 3020 1526
rect 2994 1523 3005 1524
rect 3106 1523 3173 1526
rect 3188 1523 3237 1526
rect 3276 1523 3293 1526
rect 3298 1523 3316 1526
rect 3348 1523 3357 1526
rect 3362 1523 3388 1526
rect 3410 1523 3420 1526
rect 172 1513 181 1516
rect 506 1515 509 1523
rect 580 1513 597 1516
rect 666 1513 700 1516
rect 802 1513 805 1523
rect 2490 1516 2493 1523
rect 3298 1516 3301 1523
rect 1084 1513 1109 1516
rect 1388 1513 1413 1516
rect 1436 1513 1445 1516
rect 1514 1513 1524 1516
rect 1548 1513 1557 1516
rect 1780 1513 1797 1516
rect 1956 1513 1973 1516
rect 2098 1513 2117 1516
rect 2140 1513 2157 1516
rect 2188 1513 2237 1516
rect 2418 1513 2444 1516
rect 2468 1513 2493 1516
rect 2634 1513 2661 1516
rect 2692 1513 2709 1516
rect 2762 1513 2788 1516
rect 2812 1513 2821 1516
rect 3196 1513 3205 1516
rect 3282 1513 3301 1516
rect 706 1503 716 1506
rect 1498 1503 1540 1506
rect 2154 1493 2157 1513
rect 2402 1503 2460 1506
rect 2754 1503 2804 1506
rect 2986 1503 3028 1506
rect 1154 1483 1181 1486
rect 14 1467 3506 1473
rect 2434 1443 2445 1446
rect 394 1423 405 1426
rect 402 1416 405 1423
rect 522 1423 533 1426
rect 522 1416 525 1423
rect 172 1413 197 1416
rect 204 1413 220 1416
rect 234 1413 245 1416
rect 260 1413 293 1416
rect 388 1413 397 1416
rect 402 1413 412 1416
rect 492 1413 525 1416
rect 586 1416 589 1425
rect 676 1423 685 1426
rect 1460 1423 1469 1426
rect 1700 1423 1709 1426
rect 1780 1423 1813 1426
rect 1844 1423 1893 1426
rect 1988 1423 2029 1426
rect 2260 1423 2277 1426
rect 586 1413 604 1416
rect 644 1413 653 1416
rect 194 1405 197 1413
rect 242 1395 245 1413
rect 714 1406 717 1414
rect 722 1413 732 1416
rect 738 1413 764 1416
rect 892 1413 917 1416
rect 962 1413 996 1416
rect 1090 1413 1100 1416
rect 1146 1413 1164 1416
rect 1178 1413 1229 1416
rect 1260 1413 1277 1416
rect 1380 1413 1413 1416
rect 1418 1413 1444 1416
rect 252 1403 293 1406
rect 498 1403 532 1406
rect 626 1403 636 1406
rect 714 1403 724 1406
rect 820 1403 837 1406
rect 970 1403 988 1406
rect 1044 1403 1085 1406
rect 1146 1403 1149 1413
rect 1466 1406 1469 1423
rect 1492 1413 1533 1416
rect 1538 1413 1556 1416
rect 1668 1413 1685 1416
rect 1692 1413 1757 1416
rect 1802 1413 1821 1416
rect 1866 1413 1900 1416
rect 1962 1413 1980 1416
rect 1986 1413 2036 1416
rect 2068 1413 2077 1416
rect 2154 1413 2164 1416
rect 2252 1413 2261 1416
rect 2333 1413 2365 1416
rect 2378 1413 2388 1416
rect 2412 1413 2421 1416
rect 1194 1403 1212 1406
rect 1226 1403 1236 1406
rect 1266 1403 1308 1406
rect 1322 1403 1332 1406
rect 1354 1403 1372 1406
rect 1466 1403 1525 1406
rect 1610 1403 1660 1406
rect 1674 1403 1684 1406
rect 1754 1405 1757 1413
rect 1780 1403 1813 1406
rect 1818 1405 1821 1413
rect 1844 1403 1853 1406
rect 1874 1403 1908 1406
rect 1946 1403 1972 1406
rect 2018 1403 2044 1406
rect 2074 1403 2108 1406
rect 2130 1403 2172 1406
rect 2188 1403 2229 1406
rect 2234 1403 2243 1406
rect 2258 1403 2261 1413
rect 2298 1406 2301 1413
rect 2290 1403 2301 1406
rect 2324 1403 2333 1406
rect 2338 1403 2396 1406
rect 2410 1403 2420 1406
rect 690 1393 700 1396
rect 2434 1386 2437 1443
rect 2442 1433 2492 1436
rect 3058 1433 3076 1436
rect 2442 1423 2476 1426
rect 2506 1423 2540 1426
rect 2684 1423 2725 1426
rect 3042 1423 3060 1426
rect 3084 1423 3093 1426
rect 2442 1393 2445 1423
rect 2506 1413 2525 1416
rect 2628 1413 2661 1416
rect 2690 1413 2740 1416
rect 2756 1413 2789 1416
rect 2828 1413 2861 1416
rect 2930 1413 2948 1416
rect 2980 1413 2989 1416
rect 3036 1413 3053 1416
rect 3162 1413 3188 1416
rect 3234 1413 3261 1416
rect 3268 1413 3277 1416
rect 3348 1413 3365 1416
rect 3396 1413 3405 1416
rect 2570 1403 2604 1406
rect 2658 1405 2661 1413
rect 2684 1403 2725 1406
rect 2810 1403 2820 1406
rect 2978 1403 3028 1406
rect 3162 1403 3180 1406
rect 3204 1403 3245 1406
rect 3258 1405 3261 1413
rect 3274 1405 3277 1413
rect 3300 1403 3325 1406
rect 3330 1403 3340 1406
rect 3412 1403 3429 1406
rect 3322 1396 3325 1403
rect 3322 1393 3332 1396
rect 3362 1393 3372 1396
rect 2434 1383 2469 1386
rect 38 1367 3482 1373
rect 194 1326 197 1335
rect 242 1326 245 1345
rect 1164 1343 1181 1346
rect 1594 1343 1604 1346
rect 2154 1343 2172 1346
rect 2450 1336 2453 1356
rect 3106 1353 3141 1356
rect 2748 1343 2757 1346
rect 3290 1343 3332 1346
rect 252 1333 277 1336
rect 386 1333 405 1336
rect 172 1323 197 1326
rect 204 1323 220 1326
rect 234 1323 245 1326
rect 316 1323 325 1326
rect 372 1323 397 1326
rect 402 1325 405 1333
rect 434 1333 445 1336
rect 468 1333 508 1336
rect 586 1333 612 1336
rect 434 1325 437 1333
rect 476 1323 509 1326
rect 634 1323 637 1335
rect 668 1333 677 1336
rect 844 1333 860 1336
rect 876 1333 909 1336
rect 1018 1333 1036 1336
rect 1058 1326 1061 1335
rect 1098 1333 1148 1336
rect 1170 1333 1195 1336
rect 1234 1333 1292 1336
rect 1308 1333 1317 1336
rect 1322 1333 1356 1336
rect 1388 1333 1421 1336
rect 1426 1333 1436 1336
rect 1460 1333 1477 1336
rect 1506 1333 1516 1336
rect 1554 1333 1580 1336
rect 1612 1333 1637 1336
rect 1642 1333 1660 1336
rect 1698 1333 1732 1336
rect 1756 1333 1813 1336
rect 1986 1333 1996 1336
rect 2018 1333 2052 1336
rect 2074 1333 2116 1336
rect 2138 1333 2180 1336
rect 2338 1333 2404 1336
rect 2426 1333 2453 1336
rect 2490 1333 2508 1336
rect 2602 1333 2612 1336
rect 2714 1333 2732 1336
rect 2818 1333 2868 1336
rect 2890 1333 2932 1336
rect 2948 1333 2957 1336
rect 3050 1333 3084 1336
rect 3114 1333 3156 1336
rect 3172 1333 3181 1336
rect 3186 1333 3260 1336
rect 3340 1333 3365 1336
rect 3370 1333 3388 1336
rect 810 1323 828 1326
rect 884 1323 909 1326
rect 948 1323 965 1326
rect 1026 1323 1044 1326
rect 1058 1323 1069 1326
rect 1114 1323 1140 1326
rect 1164 1323 1173 1326
rect 1186 1323 1203 1326
rect 1258 1323 1284 1326
rect 1316 1323 1333 1326
rect 1394 1323 1444 1326
rect 1458 1323 1484 1326
rect 1540 1323 1557 1326
rect 1562 1323 1588 1326
rect 1620 1323 1629 1326
rect 1650 1323 1668 1326
rect 1698 1323 1740 1326
rect 1802 1323 1812 1326
rect 1844 1323 1869 1326
rect 668 1313 677 1316
rect 1092 1313 1133 1316
rect 1170 1306 1173 1323
rect 1554 1316 1557 1323
rect 1554 1313 1573 1316
rect 1756 1313 1797 1316
rect 1914 1306 1917 1325
rect 1962 1323 1988 1326
rect 2034 1323 2060 1326
rect 2098 1323 2108 1326
rect 2202 1323 2236 1326
rect 2268 1323 2277 1326
rect 2290 1323 2308 1326
rect 2340 1323 2365 1326
rect 2386 1323 2396 1326
rect 2428 1323 2437 1326
rect 2442 1323 2468 1326
rect 2474 1323 2516 1326
rect 2434 1316 2437 1323
rect 1932 1313 1941 1316
rect 2068 1313 2101 1316
rect 2434 1313 2445 1316
rect 2476 1313 2501 1316
rect 2538 1313 2572 1316
rect 2578 1306 2581 1325
rect 2620 1323 2629 1326
rect 2714 1316 2717 1333
rect 3114 1326 3117 1333
rect 2748 1323 2789 1326
rect 2796 1323 2805 1326
rect 2956 1323 2989 1326
rect 3092 1323 3117 1326
rect 3122 1323 3148 1326
rect 3180 1323 3213 1326
rect 3234 1323 3252 1326
rect 3284 1323 3301 1326
rect 3410 1323 3420 1326
rect 2692 1313 2717 1316
rect 2802 1313 2805 1323
rect 2970 1313 3012 1316
rect 3036 1313 3069 1316
rect 3100 1313 3109 1316
rect 1170 1303 1181 1306
rect 1906 1303 1917 1306
rect 1938 1303 1981 1306
rect 2562 1303 2581 1306
rect 2634 1303 2684 1306
rect 3010 1303 3028 1306
rect 14 1267 3506 1273
rect 602 1233 620 1236
rect 1634 1233 1660 1236
rect 2194 1233 2220 1236
rect 2386 1233 2405 1236
rect 3298 1233 3340 1236
rect 586 1223 613 1226
rect 1244 1223 1285 1226
rect 1602 1223 1653 1226
rect 1796 1223 1821 1226
rect 1844 1223 1885 1226
rect 2044 1223 2077 1226
rect 2386 1223 2396 1226
rect 586 1216 589 1223
rect 124 1213 149 1216
rect 180 1213 221 1216
rect 228 1213 244 1216
rect 412 1213 453 1216
rect 466 1213 476 1216
rect 482 1213 500 1216
rect 506 1213 540 1216
rect 572 1213 589 1216
rect 788 1213 805 1216
rect 852 1213 877 1216
rect 972 1213 989 1216
rect 1042 1213 1068 1216
rect 1100 1213 1149 1216
rect 1210 1213 1228 1216
rect 1330 1213 1365 1216
rect 1372 1213 1389 1216
rect 1396 1213 1437 1216
rect 1460 1213 1477 1216
rect 1482 1213 1492 1216
rect 1516 1213 1541 1216
rect 1596 1213 1637 1216
rect 1708 1213 1773 1216
rect 1794 1213 1836 1216
rect 1908 1213 1917 1216
rect 1922 1213 1940 1216
rect 2082 1213 2092 1216
rect 2130 1213 2165 1216
rect 2268 1213 2285 1216
rect 2290 1213 2316 1216
rect 2348 1213 2365 1216
rect 2402 1215 2405 1233
rect 2476 1223 2509 1226
rect 2596 1223 2605 1226
rect 2692 1223 2701 1226
rect 2876 1223 2885 1226
rect 2932 1223 2941 1226
rect 3122 1223 3133 1226
rect 3228 1223 3237 1226
rect 3258 1223 3277 1226
rect 3348 1223 3373 1226
rect 2482 1213 2524 1216
rect 2660 1213 2669 1216
rect 2698 1213 2701 1223
rect 3130 1216 3133 1223
rect 3258 1216 3261 1223
rect 3378 1216 3381 1246
rect 2746 1213 2764 1216
rect 2924 1213 2933 1216
rect 3004 1213 3013 1216
rect 3018 1213 3052 1216
rect 3100 1213 3125 1216
rect 3130 1213 3140 1216
rect 3170 1213 3261 1216
rect 3266 1213 3277 1216
rect 3378 1213 3396 1216
rect 218 1205 221 1213
rect 276 1203 309 1206
rect 426 1203 452 1206
rect 506 1183 509 1213
rect 538 1203 548 1206
rect 564 1203 589 1206
rect 780 1203 797 1206
rect 1042 1203 1060 1206
rect 1138 1203 1148 1206
rect 1180 1203 1220 1206
rect 1244 1203 1277 1206
rect 1282 1203 1300 1206
rect 1362 1205 1365 1213
rect 1378 1203 1388 1206
rect 1452 1203 1461 1206
rect 1564 1203 1581 1206
rect 1588 1203 1629 1206
rect 1674 1203 1700 1206
rect 1762 1203 1772 1206
rect 1796 1203 1805 1206
rect 1858 1203 1884 1206
rect 1964 1203 1981 1206
rect 2010 1203 2020 1206
rect 2044 1203 2053 1206
rect 2116 1203 2157 1206
rect 2162 1205 2165 1213
rect 2234 1203 2260 1206
rect 2274 1203 2301 1206
rect 2482 1203 2516 1206
rect 2540 1203 2549 1206
rect 2562 1203 2572 1206
rect 2642 1203 2652 1206
rect 2714 1203 2756 1206
rect 2810 1203 2820 1206
rect 2874 1203 2916 1206
rect 2930 1203 2933 1213
rect 3018 1206 3021 1213
rect 3130 1206 3133 1213
rect 3170 1206 3173 1213
rect 3002 1203 3021 1206
rect 3034 1203 3044 1206
rect 3066 1203 3092 1206
rect 3106 1203 3133 1206
rect 3162 1203 3173 1206
rect 3178 1203 3212 1206
rect 3274 1205 3277 1213
rect 3362 1203 3388 1206
rect 3412 1203 3421 1206
rect 586 1183 589 1203
rect 794 1193 797 1203
rect 1282 1196 1285 1203
rect 1274 1193 1285 1196
rect 1410 1193 1444 1196
rect 1522 1193 1556 1196
rect 2602 1193 2644 1196
rect 3004 1193 3013 1196
rect 2706 1183 2741 1186
rect 38 1167 3482 1173
rect 2458 1153 2485 1156
rect 378 1133 396 1136
rect 412 1133 429 1136
rect 442 1133 452 1136
rect 474 1127 477 1134
rect 556 1133 589 1136
rect 618 1133 636 1136
rect 788 1133 797 1136
rect 1026 1133 1060 1136
rect 1116 1133 1157 1136
rect 1178 1133 1196 1136
rect 1266 1133 1292 1136
rect 1314 1133 1348 1136
rect 1380 1133 1429 1136
rect 1468 1133 1485 1136
rect 1546 1133 1564 1136
rect 124 1123 149 1126
rect 180 1123 197 1126
rect 236 1123 245 1126
rect 292 1123 317 1126
rect 372 1123 381 1126
rect 434 1123 460 1126
rect 474 1124 492 1127
rect 1586 1126 1589 1134
rect 1594 1133 1604 1136
rect 1626 1133 1652 1136
rect 666 1123 700 1126
rect 746 1123 756 1126
rect 802 1123 812 1126
rect 876 1123 901 1126
rect 946 1123 972 1126
rect 994 1123 1004 1126
rect 1026 1123 1068 1126
rect 1082 1123 1100 1126
rect 1114 1123 1156 1126
rect 1180 1123 1197 1126
rect 1204 1123 1213 1126
rect 1218 1123 1244 1126
rect 1300 1123 1341 1126
rect 1356 1123 1373 1126
rect 1388 1123 1413 1126
rect 1426 1123 1444 1126
rect 1538 1123 1572 1126
rect 1586 1123 1605 1126
rect 1660 1123 1669 1126
rect 1674 1116 1677 1134
rect 1690 1133 1724 1136
rect 1738 1133 1756 1136
rect 1770 1133 1796 1136
rect 1884 1133 1901 1136
rect 1954 1133 1964 1136
rect 1988 1133 2013 1136
rect 2042 1126 2045 1134
rect 2050 1133 2084 1136
rect 2098 1133 2108 1136
rect 2122 1133 2172 1136
rect 2298 1133 2333 1136
rect 2356 1133 2373 1136
rect 2378 1133 2388 1136
rect 2458 1133 2500 1136
rect 2522 1133 2564 1136
rect 2370 1126 2373 1133
rect 2586 1126 2589 1134
rect 2610 1133 2620 1136
rect 2634 1133 2652 1136
rect 2682 1133 2700 1136
rect 2722 1133 2772 1136
rect 2786 1133 2804 1136
rect 2818 1133 2876 1136
rect 2892 1133 2901 1136
rect 2930 1133 2973 1136
rect 3050 1133 3060 1136
rect 3076 1133 3085 1136
rect 3122 1133 3140 1136
rect 3218 1133 3284 1136
rect 3322 1133 3332 1136
rect 3362 1133 3388 1136
rect 1684 1123 1717 1126
rect 1732 1123 1757 1126
rect 1764 1123 1789 1126
rect 1794 1123 1804 1126
rect 1818 1123 1860 1126
rect 1922 1123 1932 1126
rect 2042 1123 2069 1126
rect 2154 1123 2164 1126
rect 2196 1123 2205 1126
rect 2258 1123 2276 1126
rect 2282 1123 2330 1126
rect 2370 1123 2396 1126
rect 2524 1123 2557 1126
rect 2572 1123 2589 1126
rect 2596 1123 2621 1126
rect 2628 1123 2653 1126
rect 2660 1123 2692 1126
rect 2780 1123 2805 1126
rect 2812 1123 2861 1126
rect 2900 1123 2909 1126
rect 2924 1123 2965 1126
rect 2970 1125 2973 1133
rect 3004 1123 3013 1126
rect 3042 1123 3052 1126
rect 3090 1123 3148 1126
rect 3234 1123 3276 1126
rect 3340 1123 3396 1126
rect 3402 1123 3412 1126
rect 508 1113 525 1116
rect 1308 1113 1349 1116
rect 1588 1113 1597 1116
rect 1668 1113 1677 1116
rect 1820 1113 1853 1116
rect 1948 1113 1957 1116
rect 1988 1113 2013 1116
rect 2260 1113 2269 1116
rect 2284 1113 2301 1116
rect 2404 1113 2421 1116
rect 2426 1106 2429 1115
rect 2820 1113 2853 1116
rect 2906 1113 2909 1123
rect 3156 1113 3181 1116
rect 3212 1113 3221 1116
rect 3420 1113 3429 1116
rect 490 1103 500 1106
rect 2418 1103 2429 1106
rect 2730 1093 2757 1096
rect 14 1067 3506 1073
rect 2338 1033 2372 1036
rect 2762 1026 2765 1056
rect 2850 1033 2860 1036
rect 276 1023 301 1026
rect 386 1016 389 1026
rect 540 1023 549 1026
rect 674 1016 677 1025
rect 1028 1023 1045 1026
rect 1244 1023 1253 1026
rect 1940 1023 1973 1026
rect 2322 1023 2356 1026
rect 2444 1023 2477 1026
rect 2748 1023 2765 1026
rect 2828 1023 2844 1026
rect 3044 1023 3053 1026
rect 3332 1023 3365 1026
rect 108 1013 117 1016
rect 220 1013 229 1016
rect 114 995 117 1013
rect 124 1003 133 1006
rect 130 993 133 1003
rect 226 995 229 1013
rect 346 1006 349 1014
rect 380 1013 389 1016
rect 434 1006 437 1014
rect 468 1013 477 1016
rect 532 1013 541 1016
rect 556 1013 573 1016
rect 578 1013 588 1016
rect 634 1013 660 1016
rect 674 1013 685 1016
rect 706 1013 748 1016
rect 788 1013 797 1016
rect 876 1013 901 1016
rect 938 1013 972 1016
rect 986 1013 997 1016
rect 1026 1013 1068 1016
rect 1148 1013 1157 1016
rect 682 1006 685 1013
rect 994 1006 997 1013
rect 1162 1006 1165 1014
rect 1188 1013 1197 1016
rect 1258 1013 1269 1016
rect 1356 1013 1373 1016
rect 1380 1013 1437 1016
rect 1460 1013 1475 1016
rect 1652 1013 1669 1016
rect 1676 1013 1717 1016
rect 1796 1013 1812 1016
rect 1834 1013 1884 1016
rect 1898 1013 1924 1016
rect 1970 1013 1988 1016
rect 2028 1013 2061 1016
rect 1258 1006 1261 1013
rect 1434 1007 1437 1013
rect 298 1003 316 1006
rect 338 1003 349 1006
rect 378 1003 428 1006
rect 434 1003 445 1006
rect 466 1003 476 1006
rect 682 1003 692 1006
rect 722 1003 740 1006
rect 786 1003 796 1006
rect 994 1003 1004 1006
rect 1028 1003 1053 1006
rect 1140 1003 1165 1006
rect 1210 1003 1220 1006
rect 1244 1003 1261 1006
rect 1292 1003 1317 1006
rect 1338 1003 1348 1006
rect 1362 1003 1372 1006
rect 1602 1003 1644 1006
rect 1658 1003 1668 1006
rect 1682 1003 1716 1006
rect 1740 1003 1757 1006
rect 1762 1003 1780 1006
rect 1834 1003 1876 1006
rect 1898 1005 1901 1013
rect 2066 1006 2069 1014
rect 2172 1013 2196 1016
rect 2268 1013 2277 1016
rect 2316 1013 2349 1016
rect 2426 1013 2436 1016
rect 2492 1013 2501 1016
rect 2746 1013 2788 1016
rect 2820 1013 2837 1016
rect 2972 1013 2989 1016
rect 3010 1013 3036 1016
rect 3164 1013 3189 1016
rect 3234 1013 3268 1016
rect 3346 1013 3380 1016
rect 2026 1003 2069 1006
rect 2098 1003 2108 1006
rect 2178 1003 2188 1006
rect 2282 1003 2292 1006
rect 2308 1003 2317 1006
rect 2418 1003 2428 1006
rect 2458 1003 2484 1006
rect 2524 1003 2533 1006
rect 2540 1003 2557 1006
rect 2708 1003 2724 1006
rect 2794 1003 2812 1006
rect 2898 1003 2924 1006
rect 2938 1003 2948 1006
rect 2970 1003 3028 1006
rect 3042 1003 3076 1006
rect 3156 1003 3188 1006
rect 3218 1003 3276 1006
rect 3298 1003 3308 1006
rect 3386 1003 3396 1006
rect 386 993 420 996
rect 490 993 517 996
rect 1188 993 1213 996
rect 3092 993 3125 996
rect 3292 993 3301 996
rect 38 967 3482 973
rect 1474 953 1493 956
rect 444 943 453 946
rect 682 943 725 946
rect 330 933 340 936
rect 394 933 428 936
rect 458 933 468 936
rect 530 926 533 934
rect 562 926 565 934
rect 666 933 676 936
rect 116 923 141 926
rect 236 923 261 926
rect 314 923 332 926
rect 356 923 365 926
rect 490 923 533 926
rect 554 923 565 926
rect 682 925 685 943
rect 690 933 732 936
rect 746 933 756 936
rect 770 933 780 936
rect 884 933 893 936
rect 914 926 917 946
rect 1898 936 1901 945
rect 2738 936 2741 946
rect 3004 943 3021 946
rect 930 933 940 936
rect 954 933 996 936
rect 1052 933 1069 936
rect 1082 933 1100 936
rect 1122 926 1125 934
rect 1194 933 1204 936
rect 1228 933 1237 936
rect 1290 933 1308 936
rect 1330 933 1340 936
rect 1370 933 1380 936
rect 1410 926 1413 934
rect 1436 933 1444 936
rect 1498 926 1501 934
rect 1530 933 1540 936
rect 1554 926 1557 934
rect 1578 933 1604 936
rect 1618 933 1636 936
rect 1706 926 1709 934
rect 1732 933 1757 936
rect 1796 933 1805 936
rect 1810 933 1820 936
rect 1844 933 1861 936
rect 1892 933 1901 936
rect 1930 933 1948 936
rect 1994 933 2028 936
rect 2034 933 2052 936
rect 2098 933 2108 936
rect 2132 933 2141 936
rect 2202 933 2212 936
rect 2226 933 2236 936
rect 2314 933 2332 936
rect 2348 933 2389 936
rect 2420 933 2429 936
rect 2434 933 2444 936
rect 2226 926 2229 933
rect 2530 926 2533 936
rect 2554 933 2572 936
rect 2666 933 2684 936
rect 2738 934 2780 936
rect 2738 933 2781 934
rect 2802 933 2812 936
rect 706 923 740 926
rect 754 923 764 926
rect 804 923 829 926
rect 892 923 901 926
rect 908 923 941 926
rect 1018 923 1036 926
rect 1114 923 1125 926
rect 1164 923 1173 926
rect 1194 923 1212 926
rect 1236 923 1245 926
rect 1276 923 1301 926
rect 1316 923 1341 926
rect 1348 923 1357 926
rect 1388 923 1413 926
rect 1468 923 1501 926
rect 1530 923 1557 926
rect 1564 923 1597 926
rect 1612 923 1637 926
rect 1644 923 1653 926
rect 1668 923 1709 926
rect 1730 923 1772 926
rect 1818 923 1828 926
rect 1850 923 1876 926
rect 1922 923 1956 926
rect 1970 923 1988 926
rect 2036 923 2053 926
rect 2090 923 2116 926
rect 2220 923 2229 926
rect 2250 923 2276 926
rect 2356 923 2396 926
rect 2428 923 2437 926
rect 2530 923 2548 926
rect 2596 923 2605 926
rect 492 913 501 916
rect 610 913 636 916
rect 1114 915 1117 923
rect 1402 903 1405 923
rect 1530 916 1533 923
rect 1524 913 1533 916
rect 1732 913 1749 916
rect 1844 913 1853 916
rect 1970 915 1973 923
rect 2434 916 2437 923
rect 2434 913 2445 916
rect 2602 913 2620 916
rect 2626 906 2629 925
rect 2666 916 2669 933
rect 2700 923 2709 926
rect 2716 923 2741 926
rect 2778 916 2781 933
rect 2836 923 2877 926
rect 2644 913 2669 916
rect 2770 913 2781 916
rect 2850 913 2884 916
rect 2618 903 2629 906
rect 2730 903 2749 906
rect 2730 893 2733 903
rect 2770 896 2773 913
rect 2842 903 2900 906
rect 2914 903 2917 934
rect 3058 926 3061 934
rect 3090 933 3124 936
rect 3146 933 3164 936
rect 3178 933 3212 936
rect 3226 933 3260 936
rect 3290 926 3293 934
rect 2924 923 2933 926
rect 2938 923 2980 926
rect 3004 923 3013 926
rect 3052 923 3061 926
rect 3082 923 3132 926
rect 3162 923 3172 926
rect 3186 923 3220 926
rect 3284 923 3293 926
rect 3306 923 3348 926
rect 3354 923 3364 926
rect 3378 923 3412 926
rect 2932 913 2973 916
rect 3140 913 3157 916
rect 3180 913 3213 916
rect 3228 913 3261 916
rect 2746 893 2773 896
rect 14 867 3506 873
rect 1186 853 1205 856
rect 1130 833 1141 836
rect 108 813 125 816
rect 252 813 285 816
rect 324 813 340 816
rect 492 813 525 816
rect 562 813 573 816
rect 716 813 725 816
rect 772 813 797 816
rect 834 813 860 816
rect 932 813 957 816
rect 1002 813 1020 816
rect 1092 813 1109 816
rect 1114 813 1124 816
rect 1138 815 1141 833
rect 1186 813 1197 816
rect 100 803 157 806
rect 300 803 309 806
rect 364 803 389 806
rect 498 803 524 806
rect 562 805 565 813
rect 596 803 613 806
rect 876 803 885 806
rect 1194 796 1197 813
rect 1202 806 1205 853
rect 1578 833 1613 836
rect 2682 833 2724 836
rect 2818 833 2860 836
rect 3346 833 3404 836
rect 1226 816 1229 825
rect 1314 816 1317 826
rect 1586 823 1604 826
rect 1226 813 1237 816
rect 1250 806 1253 814
rect 1274 813 1317 816
rect 1426 806 1429 816
rect 1434 813 1452 816
rect 1482 806 1485 816
rect 1202 803 1212 806
rect 1250 803 1276 806
rect 1332 803 1341 806
rect 1370 803 1396 806
rect 1412 803 1429 806
rect 1476 803 1485 806
rect 1490 806 1493 816
rect 1538 813 1548 816
rect 1572 813 1597 816
rect 1610 815 1613 833
rect 1860 823 1885 826
rect 1980 823 1997 826
rect 2098 823 2109 826
rect 2676 823 2701 826
rect 2804 823 2837 826
rect 3036 823 3045 826
rect 3132 823 3197 826
rect 3236 823 3269 826
rect 3370 823 3388 826
rect 1634 813 1644 816
rect 1708 813 1717 816
rect 1732 813 1749 816
rect 1756 813 1805 816
rect 1834 813 1844 816
rect 1940 813 1964 816
rect 2042 813 2053 816
rect 2092 813 2101 816
rect 2050 806 2053 813
rect 2106 806 2109 823
rect 3266 816 3269 823
rect 2164 813 2181 816
rect 2186 813 2204 816
rect 2210 813 2228 816
rect 2234 813 2244 816
rect 2250 813 2276 816
rect 2402 813 2412 816
rect 2588 813 2629 816
rect 2644 813 2653 816
rect 2770 813 2780 816
rect 2882 813 2900 816
rect 1490 803 1499 806
rect 1660 803 1693 806
rect 1738 803 1748 806
rect 1762 803 1804 806
rect 2002 803 2020 806
rect 2050 803 2084 806
rect 2106 803 2116 806
rect 2130 803 2140 806
rect 2162 803 2196 806
rect 2210 803 2220 806
rect 2300 803 2325 806
rect 2378 803 2420 806
rect 2506 803 2516 806
rect 1186 793 1197 796
rect 1298 793 1324 796
rect 2626 795 2629 813
rect 2930 806 2933 814
rect 2938 813 2964 816
rect 2970 813 3004 816
rect 3018 813 3028 816
rect 3042 813 3100 816
rect 3186 813 3204 816
rect 3218 813 3228 816
rect 3266 813 3292 816
rect 3330 813 3340 816
rect 3428 813 3445 816
rect 2636 803 2652 806
rect 2738 803 2748 806
rect 2930 803 2941 806
rect 2946 803 2956 806
rect 3010 803 3020 806
rect 3106 803 3116 806
rect 3146 803 3196 806
rect 2938 796 2941 803
rect 2938 793 2949 796
rect 38 767 3482 773
rect 1218 743 1228 746
rect 1242 743 1276 746
rect 1996 743 2021 746
rect 244 733 252 736
rect 402 733 436 736
rect 468 733 476 736
rect 500 733 533 736
rect 594 733 604 736
rect 724 733 749 736
rect 1010 733 1020 736
rect 1178 733 1188 736
rect 1236 733 1269 736
rect 132 723 157 726
rect 194 723 220 726
rect 250 723 260 726
rect 434 723 444 726
rect 732 723 773 726
rect 812 723 821 726
rect 924 723 941 726
rect 986 723 1028 726
rect 1068 723 1093 726
rect 500 713 541 716
rect 548 713 557 716
rect 1074 713 1100 716
rect 1074 683 1077 713
rect 1106 706 1109 725
rect 1178 716 1181 733
rect 1196 723 1205 726
rect 1212 723 1221 726
rect 1322 723 1325 734
rect 1338 733 1356 736
rect 1388 733 1397 736
rect 1402 733 1412 736
rect 1490 733 1499 736
rect 1514 733 1524 736
rect 1548 733 1581 736
rect 1586 726 1589 734
rect 1746 733 1764 736
rect 1788 733 1820 736
rect 1834 733 1844 736
rect 1954 733 1980 736
rect 2002 733 2028 736
rect 2052 733 2060 736
rect 2098 733 2124 736
rect 2242 733 2284 736
rect 2442 733 2460 736
rect 1338 723 1364 726
rect 1434 723 1460 726
rect 1476 723 1485 726
rect 1516 723 1525 726
rect 1546 723 1589 726
rect 1602 723 1612 726
rect 1658 723 1668 726
rect 1882 723 1900 726
rect 1948 723 1972 726
rect 1996 723 2029 726
rect 2148 723 2165 726
rect 2282 723 2292 726
rect 2298 723 2316 726
rect 2322 723 2348 726
rect 2450 723 2468 726
rect 1124 713 1133 716
rect 1148 713 1157 716
rect 1172 713 1181 716
rect 1324 713 1333 716
rect 1338 706 1341 723
rect 2490 716 2493 734
rect 2514 733 2524 736
rect 2546 733 2564 736
rect 2604 733 2621 736
rect 2650 733 2660 736
rect 2674 733 2684 736
rect 2794 733 2820 736
rect 2954 733 2972 736
rect 2988 733 3005 736
rect 3010 733 3020 736
rect 3162 733 3172 736
rect 3002 726 3005 733
rect 2532 723 2556 726
rect 2612 723 2645 726
rect 2676 723 2685 726
rect 2748 723 2765 726
rect 2772 723 2805 726
rect 2940 723 2964 726
rect 3002 723 3028 726
rect 3082 723 3100 726
rect 3140 723 3173 726
rect 3338 723 3373 726
rect 2236 713 2245 716
rect 2300 713 2309 716
rect 2324 713 2333 716
rect 2402 713 2412 716
rect 2476 713 2493 716
rect 2762 713 2765 723
rect 3108 713 3117 716
rect 3154 713 3157 723
rect 3370 716 3373 723
rect 3188 713 3197 716
rect 3266 713 3276 716
rect 3370 713 3389 716
rect 1082 703 1109 706
rect 1130 703 1164 706
rect 1330 703 1341 706
rect 3370 703 3396 706
rect 3410 703 3428 706
rect 14 667 3506 673
rect 1114 633 1140 636
rect 1594 633 1612 636
rect 2570 633 2588 636
rect 3010 633 3036 636
rect 1562 623 1596 626
rect 1716 623 1725 626
rect 1740 623 1749 626
rect 1970 623 1980 626
rect 2562 623 2572 626
rect 3130 623 3149 626
rect 146 613 156 616
rect 162 613 228 616
rect 340 613 357 616
rect 396 613 421 616
rect 428 613 437 616
rect 692 613 709 616
rect 762 613 772 616
rect 804 613 829 616
rect 868 613 877 616
rect 932 613 957 616
rect 994 613 1020 616
rect 1084 613 1101 616
rect 1180 613 1213 616
rect 1228 613 1237 616
rect 1292 613 1301 616
rect 1330 613 1340 616
rect 1396 613 1405 616
rect 1460 613 1493 616
rect 1556 613 1589 616
rect 1626 613 1636 616
rect 1658 613 1692 616
rect 1756 613 1781 616
rect 1786 613 1812 616
rect 2010 613 2036 616
rect 2050 613 2068 616
rect 2082 613 2125 616
rect 2146 613 2157 616
rect 2164 613 2173 616
rect 2178 613 2196 616
rect 2282 613 2292 616
rect 2354 613 2388 616
rect 2460 613 2469 616
rect 234 603 252 606
rect 418 605 421 613
rect 434 595 437 613
rect 444 603 477 606
rect 714 603 732 606
rect 754 603 780 606
rect 1076 603 1093 606
rect 1220 603 1253 606
rect 1260 603 1269 606
rect 1284 603 1301 606
rect 1322 603 1332 606
rect 1394 603 1420 606
rect 1652 603 1677 606
rect 1858 603 1876 606
rect 1906 603 1940 606
rect 2010 603 2028 606
rect 2082 605 2085 613
rect 2090 603 2124 606
rect 2146 605 2149 613
rect 2236 603 2245 606
rect 2274 603 2284 606
rect 2348 603 2357 606
rect 2370 603 2380 606
rect 2466 605 2469 613
rect 2482 606 2485 616
rect 2506 613 2540 616
rect 2556 613 2565 616
rect 2658 613 2677 616
rect 2684 613 2708 616
rect 2732 613 2757 616
rect 2764 613 2789 616
rect 2836 613 2861 616
rect 2866 613 2909 616
rect 2954 613 2980 616
rect 2498 603 2532 606
rect 2618 603 2636 606
rect 2660 603 2669 606
rect 2674 605 2677 613
rect 2906 606 2909 613
rect 2690 603 2716 606
rect 2778 603 2812 606
rect 2834 603 2868 606
rect 2906 603 2924 606
rect 3074 603 3084 606
rect 1186 593 1212 596
rect 1226 593 1252 596
rect 2354 583 2357 603
rect 3090 596 3093 615
rect 3116 613 3133 616
rect 3146 606 3149 623
rect 3180 613 3189 616
rect 3226 613 3260 616
rect 3314 613 3324 616
rect 3372 613 3389 616
rect 3410 613 3428 616
rect 3108 603 3141 606
rect 3146 603 3172 606
rect 3196 603 3221 606
rect 2426 593 2436 596
rect 3058 593 3076 596
rect 3090 593 3100 596
rect 3122 593 3164 596
rect 3178 593 3188 596
rect 38 567 3482 573
rect 2402 553 2421 556
rect 202 526 205 534
rect 218 526 221 545
rect 1788 543 1797 546
rect 2314 536 2317 546
rect 228 533 261 536
rect 388 533 405 536
rect 1010 533 1028 536
rect 1212 533 1237 536
rect 1244 533 1285 536
rect 1290 533 1300 536
rect 1484 533 1525 536
rect 1586 533 1604 536
rect 1708 533 1716 536
rect 1754 533 1772 536
rect 1836 533 1844 536
rect 1938 533 1948 536
rect 2036 533 2044 536
rect 2164 533 2173 536
rect 2212 533 2220 536
rect 2314 533 2324 536
rect 2362 533 2372 536
rect 180 523 205 526
rect 212 523 221 526
rect 500 523 525 526
rect 578 523 612 526
rect 660 523 677 526
rect 828 523 853 526
rect 940 523 965 526
rect 1002 523 1036 526
rect 1220 523 1229 526
rect 1426 523 1444 526
rect 1506 523 1540 526
rect 1612 523 1621 526
rect 1666 523 1692 526
rect 1738 523 1764 526
rect 1788 523 1813 526
rect 1930 523 1940 526
rect 1978 523 2020 526
rect 2162 523 2196 526
rect 2218 523 2228 526
rect 2298 523 2332 526
rect 2402 516 2405 553
rect 2594 543 2620 546
rect 2682 543 2716 546
rect 2474 533 2492 536
rect 2724 533 2749 536
rect 2794 533 2812 536
rect 2826 533 2852 536
rect 2884 533 2909 536
rect 3018 533 3068 536
rect 3146 533 3156 536
rect 3180 533 3213 536
rect 2410 523 2436 526
rect 2482 523 2500 526
rect 2572 523 2581 526
rect 2588 523 2597 526
rect 2676 523 2717 526
rect 2746 523 2764 526
rect 2802 523 2820 526
rect 3018 523 3076 526
rect 3082 523 3092 526
rect 3140 523 3157 526
rect 3218 523 3228 526
rect 3242 523 3260 526
rect 3274 523 3316 526
rect 3346 523 3364 526
rect 506 513 532 516
rect 1084 513 1093 516
rect 1098 513 1116 516
rect 1154 513 1172 516
rect 1412 513 1421 516
rect 1868 513 1893 516
rect 2108 513 2117 516
rect 2236 513 2253 516
rect 2402 513 2413 516
rect 1090 503 1132 506
rect 2098 503 2124 506
rect 2594 503 2597 523
rect 2746 503 2749 523
rect 3242 515 3245 523
rect 3346 515 3349 523
rect 3372 513 3389 516
rect 14 467 3506 473
rect 530 433 564 436
rect 698 433 748 436
rect 324 423 349 426
rect 364 423 389 426
rect 548 423 557 426
rect 692 423 732 426
rect 794 423 812 426
rect 1130 423 1164 426
rect 1194 425 1197 436
rect 1250 433 1276 436
rect 2034 433 2052 436
rect 2506 433 2524 436
rect 3226 433 3252 436
rect 1234 423 1260 426
rect 2036 423 2045 426
rect 2132 423 2141 426
rect 2276 423 2317 426
rect 346 416 349 423
rect 386 416 389 423
rect 794 416 797 423
rect 188 413 213 416
rect 244 413 285 416
rect 292 413 308 416
rect 346 413 356 416
rect 386 413 404 416
rect 596 413 605 416
rect 666 413 684 416
rect 772 413 797 416
rect 892 413 933 416
rect 972 413 989 416
rect 1034 413 1060 416
rect 1124 413 1172 416
rect 1306 413 1348 416
rect 1404 413 1429 416
rect 1434 413 1452 416
rect 1562 413 1572 416
rect 1612 413 1645 416
rect 1652 413 1669 416
rect 1714 413 1772 416
rect 1794 413 1804 416
rect 1810 413 1820 416
rect 1826 413 1884 416
rect 1908 413 1925 416
rect 2066 413 2124 416
rect 2164 413 2189 416
rect 2194 413 2237 416
rect 2244 413 2261 416
rect 2268 413 2301 416
rect 282 405 285 413
rect 338 403 348 406
rect 410 403 420 406
rect 634 403 644 406
rect 866 403 884 406
rect 1314 403 1332 406
rect 1378 403 1388 406
rect 1578 403 1604 406
rect 1618 403 1644 406
rect 1666 403 1669 413
rect 2314 406 2317 423
rect 1722 403 1764 406
rect 1826 403 1892 406
rect 1962 403 2004 406
rect 2066 403 2116 406
rect 2130 403 2140 406
rect 2170 403 2196 406
rect 2250 403 2260 406
rect 2298 405 2317 406
rect 2330 406 2333 425
rect 2508 423 2517 426
rect 2532 423 2565 426
rect 3218 423 3236 426
rect 2362 413 2388 416
rect 2476 413 2516 416
rect 2538 413 2572 416
rect 2708 413 2733 416
rect 2818 413 2829 416
rect 2866 413 2908 416
rect 3098 413 3140 416
rect 3330 413 3348 416
rect 2298 403 2316 405
rect 2330 403 2348 406
rect 2418 403 2452 406
rect 2826 405 2829 413
rect 2882 403 2900 406
rect 2964 403 2997 406
rect 3170 403 3180 406
rect 436 393 445 396
rect 1370 393 1380 396
rect 38 367 3482 373
rect 330 326 333 345
rect 452 343 469 346
rect 474 343 484 346
rect 474 336 477 343
rect 1314 336 1317 346
rect 1978 336 1981 345
rect 2074 336 2077 345
rect 340 333 349 336
rect 410 333 436 336
rect 450 333 477 336
rect 652 333 669 336
rect 698 333 740 336
rect 756 333 765 336
rect 770 333 788 336
rect 826 333 860 336
rect 890 333 900 336
rect 116 323 141 326
rect 172 323 205 326
rect 244 323 253 326
rect 300 323 333 326
rect 364 323 381 326
rect 418 323 428 326
rect 452 323 461 326
rect 500 323 525 326
rect 666 325 669 333
rect 914 326 917 334
rect 930 333 964 336
rect 1284 333 1317 336
rect 1418 333 1452 336
rect 1514 333 1524 336
rect 1972 333 1981 336
rect 2066 333 2077 336
rect 2084 333 2109 336
rect 2210 333 2220 336
rect 2284 333 2308 336
rect 2362 333 2380 336
rect 2730 333 2756 336
rect 2922 333 2948 336
rect 3138 333 3172 336
rect 1162 326 1180 327
rect 1226 326 1244 327
rect 700 323 725 326
rect 778 323 796 326
rect 858 323 868 326
rect 908 323 917 326
rect 1084 323 1109 326
rect 1140 324 1180 326
rect 1212 324 1244 326
rect 1140 323 1165 324
rect 1212 323 1229 324
rect 1356 323 1381 326
rect 1498 323 1508 326
rect 1604 323 1629 326
rect 1660 323 1677 326
rect 1716 323 1741 326
rect 1828 323 1853 326
rect 2010 323 2044 326
rect 2050 323 2060 326
rect 540 313 549 316
rect 1012 313 1045 316
rect 1146 313 1172 316
rect 1226 313 1236 316
rect 986 303 1004 306
rect 1178 303 1188 306
rect 1218 303 1252 306
rect 1498 303 1501 323
rect 1890 313 1916 316
rect 2066 315 2069 333
rect 2210 326 2213 333
rect 3226 326 3229 345
rect 2148 323 2173 326
rect 2204 323 2213 326
rect 2244 323 2253 326
rect 2332 323 2357 326
rect 2362 323 2388 326
rect 2426 323 2436 326
rect 2668 323 2693 326
rect 2730 323 2764 326
rect 2844 323 2869 326
rect 2906 323 2956 326
rect 3196 323 3229 326
rect 3346 323 3372 326
rect 3386 323 3404 326
rect 3410 323 3420 326
rect 2362 313 2365 323
rect 2780 313 2805 316
rect 3410 313 3413 323
rect 1898 303 1932 306
rect 14 267 3506 273
rect 698 223 708 226
rect 2036 223 2045 226
rect 2106 216 2109 226
rect 2738 216 2741 225
rect 164 213 189 216
rect 284 213 309 216
rect 340 213 349 216
rect 362 213 380 216
rect 820 213 853 216
rect 898 213 908 216
rect 980 213 1005 216
rect 1036 213 1053 216
rect 1084 213 1101 216
rect 1196 213 1237 216
rect 1252 213 1261 216
rect 1268 213 1277 216
rect 1290 213 1300 216
rect 1364 213 1381 216
rect 1386 213 1404 216
rect 1458 213 1509 216
rect 1546 213 1580 216
rect 1636 213 1645 216
rect 1740 213 1749 216
rect 1802 213 1876 216
rect 1938 213 1948 216
rect 1978 213 2044 216
rect 2066 213 2076 216
rect 2106 213 2125 216
rect 362 206 365 213
rect 1050 206 1053 213
rect 346 203 365 206
rect 412 203 453 206
rect 842 203 860 206
rect 890 203 900 206
rect 1050 203 1060 206
rect 1234 195 1237 213
rect 1244 203 1260 206
rect 1282 203 1292 206
rect 1316 203 1341 206
rect 1466 203 1492 206
rect 1506 205 1509 213
rect 1540 203 1557 206
rect 1562 203 1572 206
rect 1602 203 1612 206
rect 1906 203 1940 206
rect 2122 205 2125 213
rect 2146 213 2157 216
rect 2210 213 2228 216
rect 2258 213 2268 216
rect 2410 213 2428 216
rect 2434 213 2444 216
rect 2508 213 2516 216
rect 2540 213 2573 216
rect 2580 213 2596 216
rect 2634 213 2676 216
rect 2690 213 2724 216
rect 2738 213 2805 216
rect 2836 213 2884 216
rect 2970 213 2988 216
rect 3060 213 3069 216
rect 3076 213 3124 216
rect 3220 213 3245 216
rect 3372 213 3445 216
rect 2146 205 2149 213
rect 2252 203 2260 206
rect 2346 203 2356 206
rect 2386 203 2420 206
rect 2500 203 2517 206
rect 2570 205 2573 213
rect 2586 203 2604 206
rect 2634 203 2668 206
rect 2698 203 2716 206
rect 2770 203 2804 206
rect 2858 203 2892 206
rect 2956 203 2973 206
rect 3004 203 3021 206
rect 3098 203 3116 206
rect 3140 203 3189 206
rect 3244 203 3277 206
rect 1562 196 1565 203
rect 1546 193 1565 196
rect 2274 193 2316 196
rect 2922 193 2948 196
rect 38 167 3482 173
rect 434 133 452 136
rect 1050 133 1060 136
rect 1306 133 1332 136
rect 1346 133 1356 136
rect 1412 133 1420 136
rect 1492 133 1500 136
rect 1540 133 1573 136
rect 1674 133 1684 136
rect 1730 133 1756 136
rect 1050 126 1053 133
rect 1786 126 1789 145
rect 1802 143 1812 146
rect 1796 133 1813 136
rect 1820 133 1845 136
rect 1946 133 1956 136
rect 2002 133 2020 136
rect 2194 133 2204 136
rect 2442 133 2460 136
rect 2554 133 2580 136
rect 2650 133 2668 136
rect 2730 133 2740 136
rect 2764 133 2789 136
rect 2866 133 2884 136
rect 2932 133 2948 136
rect 3010 133 3020 136
rect 3042 133 3076 136
rect 3098 133 3108 136
rect 3132 133 3141 136
rect 124 123 149 126
rect 186 123 212 126
rect 218 123 228 126
rect 292 123 317 126
rect 348 123 357 126
rect 548 123 573 126
rect 716 123 725 126
rect 828 123 837 126
rect 988 123 1013 126
rect 1044 123 1053 126
rect 1084 123 1093 126
rect 1188 123 1221 126
rect 1266 123 1276 126
rect 1340 123 1357 126
rect 1364 123 1381 126
rect 1418 123 1428 126
rect 1434 123 1476 126
rect 1490 123 1508 126
rect 1514 123 1524 126
rect 1612 123 1637 126
rect 1732 123 1757 126
rect 1764 123 1773 126
rect 1780 123 1789 126
rect 1882 123 1892 126
rect 1908 124 1924 127
rect 1954 123 1964 126
rect 2050 123 2060 126
rect 2154 123 2164 126
rect 2212 123 2221 126
rect 2546 123 2588 126
rect 2676 123 2685 126
rect 2770 123 2804 126
rect 2908 123 2949 126
rect 2972 123 3012 126
rect 3050 123 3068 126
rect 3100 123 3116 126
rect 3244 123 3253 126
rect 1292 113 1301 116
rect 1852 113 1861 116
rect 1940 113 1949 116
rect 2100 113 2117 116
rect 2500 113 2509 116
rect 2540 113 2589 116
rect 2604 113 2613 116
rect 2644 113 2661 116
rect 2820 113 2829 116
rect 2860 113 2877 116
rect 1834 103 1868 106
rect 1914 103 1932 106
rect 2066 103 2092 106
rect 2106 103 2140 106
rect 14 67 3506 73
rect 38 37 3482 57
rect 14 13 3506 33
<< metal2 >>
rect 14 13 34 3427
rect 38 37 58 3403
rect 266 3363 309 3366
rect 210 3343 237 3346
rect 82 3256 85 3336
rect 130 3323 133 3336
rect 82 3253 93 3256
rect 90 2776 93 3253
rect 178 3193 181 3206
rect 202 3196 205 3336
rect 210 3323 213 3343
rect 218 3333 229 3336
rect 266 3333 269 3363
rect 282 3333 285 3346
rect 226 3226 229 3316
rect 218 3223 229 3226
rect 218 3206 221 3223
rect 194 3193 205 3196
rect 214 3203 221 3206
rect 130 3086 133 3126
rect 122 3083 133 3086
rect 122 3036 125 3083
rect 138 3076 141 3116
rect 170 3113 173 3126
rect 138 3073 149 3076
rect 122 3033 133 3036
rect 130 3013 133 3033
rect 146 3026 149 3073
rect 138 3023 149 3026
rect 138 3003 141 3023
rect 194 2996 197 3193
rect 214 3146 217 3203
rect 214 3143 221 3146
rect 218 3123 221 3143
rect 226 3133 229 3216
rect 258 3156 261 3216
rect 266 3163 269 3326
rect 306 3323 309 3363
rect 682 3363 725 3366
rect 362 3293 365 3326
rect 378 3256 381 3346
rect 426 3323 429 3346
rect 466 3336 469 3346
rect 450 3333 469 3336
rect 474 3333 477 3346
rect 378 3253 389 3256
rect 306 3193 309 3206
rect 354 3193 357 3216
rect 386 3206 389 3253
rect 450 3213 453 3333
rect 466 3313 469 3326
rect 482 3303 485 3326
rect 514 3276 517 3336
rect 562 3323 565 3346
rect 634 3343 661 3346
rect 594 3333 629 3336
rect 514 3273 525 3276
rect 370 3203 389 3206
rect 370 3166 373 3203
rect 234 3153 261 3156
rect 234 3133 237 3153
rect 250 3133 253 3146
rect 258 3143 285 3146
rect 258 3123 261 3143
rect 266 3133 277 3136
rect 258 3096 261 3116
rect 250 3093 261 3096
rect 250 3036 253 3093
rect 274 3036 277 3116
rect 314 3113 317 3166
rect 362 3163 373 3166
rect 378 3163 421 3166
rect 362 3106 365 3163
rect 378 3133 381 3163
rect 362 3103 373 3106
rect 218 3023 221 3036
rect 250 3033 261 3036
rect 202 3013 221 3016
rect 210 3003 221 3006
rect 194 2993 229 2996
rect 130 2923 133 2956
rect 210 2916 213 2936
rect 218 2923 221 2936
rect 202 2913 213 2916
rect 130 2803 133 2816
rect 90 2773 101 2776
rect 98 2756 101 2773
rect 98 2753 117 2756
rect 98 2736 101 2753
rect 82 2733 101 2736
rect 114 2733 117 2753
rect 82 2646 85 2733
rect 154 2716 157 2816
rect 162 2723 165 2746
rect 154 2713 165 2716
rect 162 2676 165 2713
rect 162 2673 181 2676
rect 82 2643 101 2646
rect 98 2566 101 2643
rect 146 2593 149 2616
rect 178 2576 181 2673
rect 202 2636 205 2913
rect 202 2633 213 2636
rect 202 2603 205 2616
rect 90 2563 101 2566
rect 170 2573 181 2576
rect 90 2356 93 2563
rect 138 2513 141 2526
rect 170 2486 173 2573
rect 210 2546 213 2633
rect 218 2603 221 2626
rect 226 2606 229 2993
rect 234 2933 237 2956
rect 242 2933 245 2946
rect 234 2903 237 2916
rect 250 2823 253 2836
rect 234 2796 237 2816
rect 258 2813 261 3033
rect 270 3033 277 3036
rect 270 2966 273 3033
rect 282 3003 285 3026
rect 306 2976 309 3076
rect 370 3073 373 3103
rect 394 3073 397 3136
rect 418 3123 421 3163
rect 442 3143 445 3206
rect 466 3193 469 3206
rect 498 3043 501 3126
rect 506 3116 509 3226
rect 522 3183 525 3273
rect 570 3153 573 3216
rect 530 3133 549 3136
rect 586 3133 589 3236
rect 594 3133 597 3333
rect 634 3323 637 3343
rect 666 3336 669 3346
rect 658 3333 669 3336
rect 682 3333 685 3363
rect 650 3226 653 3316
rect 650 3223 661 3226
rect 602 3193 645 3196
rect 530 3123 541 3126
rect 506 3113 541 3116
rect 330 3013 333 3026
rect 442 3013 445 3026
rect 266 2963 273 2966
rect 290 2973 333 2976
rect 266 2893 269 2963
rect 274 2933 277 2956
rect 290 2933 293 2973
rect 314 2923 317 2956
rect 330 2916 333 2973
rect 378 2923 381 2966
rect 322 2913 333 2916
rect 242 2803 253 2806
rect 234 2793 261 2796
rect 298 2786 301 2816
rect 306 2803 309 2826
rect 298 2783 317 2786
rect 282 2736 285 2746
rect 234 2613 237 2626
rect 226 2603 237 2606
rect 242 2603 253 2606
rect 66 2353 93 2356
rect 162 2483 173 2486
rect 194 2543 213 2546
rect 234 2596 237 2603
rect 266 2596 269 2736
rect 282 2733 293 2736
rect 274 2723 285 2726
rect 298 2723 301 2746
rect 290 2713 301 2716
rect 298 2653 301 2713
rect 314 2676 317 2783
rect 322 2686 325 2913
rect 402 2853 405 2976
rect 410 2933 421 2936
rect 418 2893 421 2926
rect 426 2916 429 2936
rect 434 2923 437 2996
rect 442 2933 445 2946
rect 442 2916 445 2926
rect 426 2913 445 2916
rect 450 2886 453 3016
rect 466 3013 469 3036
rect 458 2983 461 3006
rect 466 2933 469 2956
rect 482 2926 485 3016
rect 490 2986 493 3016
rect 498 2993 501 3006
rect 490 2983 501 2986
rect 418 2883 453 2886
rect 346 2813 349 2826
rect 402 2776 405 2846
rect 402 2773 409 2776
rect 354 2763 397 2766
rect 322 2683 333 2686
rect 306 2656 309 2676
rect 314 2673 325 2676
rect 306 2653 313 2656
rect 298 2623 301 2636
rect 282 2613 301 2616
rect 234 2593 269 2596
rect 298 2593 301 2606
rect 66 2176 69 2353
rect 74 2253 77 2316
rect 90 2176 93 2346
rect 138 2313 141 2326
rect 114 2193 117 2216
rect 66 2173 77 2176
rect 90 2173 101 2176
rect 74 1966 77 2173
rect 98 1966 101 2173
rect 162 2166 165 2483
rect 194 2416 197 2543
rect 234 2536 237 2593
rect 310 2586 313 2653
rect 306 2583 313 2586
rect 210 2523 213 2536
rect 218 2533 237 2536
rect 194 2413 205 2416
rect 186 2393 197 2396
rect 186 2246 189 2366
rect 194 2323 197 2393
rect 186 2243 193 2246
rect 162 2163 169 2166
rect 146 2123 149 2136
rect 166 2086 169 2163
rect 162 2083 169 2086
rect 162 2056 165 2083
rect 162 2053 169 2056
rect 146 1993 149 2016
rect 166 1976 169 2053
rect 66 1963 77 1966
rect 90 1963 101 1966
rect 162 1973 169 1976
rect 66 1896 69 1963
rect 66 1893 77 1896
rect 74 1646 77 1893
rect 90 1756 93 1963
rect 138 1923 141 1936
rect 162 1876 165 1973
rect 178 1886 181 2236
rect 190 2186 193 2243
rect 202 2226 205 2413
rect 218 2306 221 2533
rect 242 2523 245 2536
rect 250 2533 253 2546
rect 242 2503 245 2516
rect 266 2496 269 2576
rect 298 2513 301 2536
rect 242 2493 293 2496
rect 242 2413 245 2493
rect 242 2393 245 2406
rect 258 2353 261 2406
rect 282 2393 285 2416
rect 242 2323 245 2336
rect 266 2333 269 2346
rect 218 2303 229 2306
rect 250 2303 253 2316
rect 226 2256 229 2303
rect 290 2296 293 2493
rect 306 2456 309 2583
rect 322 2573 325 2673
rect 330 2666 333 2683
rect 330 2663 337 2666
rect 334 2586 337 2663
rect 330 2583 337 2586
rect 330 2566 333 2583
rect 218 2253 229 2256
rect 282 2293 293 2296
rect 302 2453 309 2456
rect 322 2563 333 2566
rect 322 2456 325 2563
rect 322 2453 333 2456
rect 218 2233 221 2253
rect 202 2223 229 2226
rect 250 2223 253 2236
rect 218 2203 221 2216
rect 226 2206 229 2223
rect 226 2203 237 2206
rect 190 2183 205 2186
rect 202 1956 205 2183
rect 234 1966 237 2203
rect 250 2193 253 2206
rect 258 2193 261 2206
rect 242 2143 269 2146
rect 242 2123 245 2143
rect 250 2133 261 2136
rect 258 2103 261 2116
rect 258 2023 261 2036
rect 242 2013 261 2016
rect 258 1993 261 2006
rect 274 2003 277 2026
rect 154 1873 165 1876
rect 174 1883 181 1886
rect 194 1953 205 1956
rect 226 1963 237 1966
rect 154 1816 157 1873
rect 154 1813 165 1816
rect 146 1783 149 1796
rect 162 1766 165 1813
rect 174 1786 177 1883
rect 194 1876 197 1953
rect 218 1923 221 1936
rect 226 1906 229 1963
rect 282 1956 285 2293
rect 302 2286 305 2453
rect 330 2386 333 2453
rect 322 2383 333 2386
rect 346 2383 349 2736
rect 354 2733 357 2763
rect 370 2686 373 2746
rect 394 2723 397 2763
rect 406 2716 409 2773
rect 402 2713 409 2716
rect 370 2683 381 2686
rect 362 2593 365 2606
rect 378 2603 381 2683
rect 354 2513 357 2526
rect 402 2516 405 2713
rect 418 2696 421 2883
rect 434 2803 437 2816
rect 442 2786 445 2856
rect 458 2843 461 2926
rect 474 2903 477 2926
rect 482 2923 493 2926
rect 498 2923 501 2983
rect 458 2813 461 2836
rect 414 2693 421 2696
rect 438 2783 445 2786
rect 414 2636 417 2693
rect 438 2686 441 2783
rect 426 2683 441 2686
rect 414 2633 421 2636
rect 410 2593 413 2616
rect 418 2583 421 2633
rect 418 2523 421 2546
rect 394 2513 405 2516
rect 394 2456 397 2513
rect 394 2453 405 2456
rect 386 2413 389 2436
rect 394 2413 397 2426
rect 322 2363 325 2383
rect 394 2363 397 2406
rect 314 2323 317 2346
rect 330 2286 333 2356
rect 298 2283 305 2286
rect 322 2283 333 2286
rect 298 2226 301 2283
rect 290 2223 301 2226
rect 290 2176 293 2223
rect 298 2193 301 2206
rect 322 2176 325 2283
rect 346 2193 349 2216
rect 290 2173 301 2176
rect 322 2173 333 2176
rect 298 1966 301 2173
rect 314 2133 317 2146
rect 330 2056 333 2173
rect 354 2123 357 2146
rect 322 2053 333 2056
rect 322 1966 325 2053
rect 346 2013 349 2026
rect 362 1966 365 2356
rect 386 2323 389 2336
rect 394 2283 397 2336
rect 402 2266 405 2453
rect 410 2413 413 2506
rect 418 2403 421 2496
rect 426 2396 429 2683
rect 434 2506 437 2536
rect 442 2523 445 2636
rect 450 2606 453 2806
rect 458 2613 461 2796
rect 466 2763 469 2806
rect 482 2756 485 2923
rect 506 2863 509 3006
rect 514 2973 517 3106
rect 538 3013 541 3113
rect 546 3103 549 3133
rect 554 3106 557 3126
rect 602 3123 605 3193
rect 618 3133 621 3156
rect 618 3106 621 3126
rect 554 3103 565 3106
rect 562 3036 565 3103
rect 610 3103 621 3106
rect 554 3033 565 3036
rect 546 2946 549 3006
rect 554 3003 557 3033
rect 586 3013 589 3056
rect 562 2946 565 3006
rect 602 2983 605 3006
rect 610 2973 613 3103
rect 626 3036 629 3136
rect 634 3133 653 3136
rect 634 3113 637 3133
rect 650 3116 653 3133
rect 658 3123 661 3223
rect 674 3213 677 3326
rect 682 3176 685 3206
rect 698 3203 701 3356
rect 722 3323 725 3363
rect 722 3176 725 3216
rect 682 3173 725 3176
rect 650 3113 657 3116
rect 634 3086 637 3106
rect 634 3083 645 3086
rect 618 3033 629 3036
rect 522 2923 525 2936
rect 530 2933 533 2946
rect 538 2943 549 2946
rect 554 2943 565 2946
rect 538 2926 541 2943
rect 546 2933 557 2936
rect 562 2933 565 2943
rect 538 2923 565 2926
rect 570 2923 573 2936
rect 586 2933 589 2956
rect 514 2913 557 2916
rect 498 2813 501 2826
rect 514 2813 517 2913
rect 474 2753 485 2756
rect 466 2606 469 2736
rect 474 2703 477 2753
rect 482 2723 485 2746
rect 498 2736 501 2756
rect 522 2746 525 2906
rect 562 2896 565 2923
rect 554 2893 565 2896
rect 570 2913 589 2916
rect 506 2743 525 2746
rect 490 2733 525 2736
rect 506 2713 509 2726
rect 522 2723 525 2733
rect 474 2613 477 2626
rect 450 2603 461 2606
rect 466 2603 477 2606
rect 450 2533 453 2556
rect 434 2503 445 2506
rect 442 2436 445 2503
rect 434 2433 445 2436
rect 434 2403 437 2433
rect 458 2416 461 2576
rect 466 2506 469 2586
rect 474 2526 477 2603
rect 482 2533 485 2616
rect 498 2613 501 2656
rect 490 2586 493 2606
rect 490 2583 497 2586
rect 474 2523 485 2526
rect 466 2503 473 2506
rect 394 2263 405 2266
rect 410 2393 429 2396
rect 394 2176 397 2263
rect 394 2173 401 2176
rect 398 2116 401 2173
rect 398 2113 405 2116
rect 402 2093 405 2113
rect 410 2086 413 2393
rect 418 2333 421 2346
rect 426 2333 429 2346
rect 442 2336 445 2416
rect 434 2333 445 2336
rect 450 2413 461 2416
rect 434 2316 437 2333
rect 418 2263 421 2316
rect 430 2313 437 2316
rect 430 2236 433 2313
rect 442 2273 445 2326
rect 450 2283 453 2413
rect 458 2393 461 2406
rect 470 2366 473 2503
rect 482 2423 485 2523
rect 494 2516 497 2583
rect 506 2533 509 2616
rect 490 2513 497 2516
rect 490 2413 493 2513
rect 514 2496 517 2606
rect 522 2573 525 2706
rect 530 2643 533 2836
rect 554 2826 557 2893
rect 538 2626 541 2826
rect 554 2823 565 2826
rect 546 2733 549 2806
rect 562 2773 565 2823
rect 570 2813 573 2913
rect 586 2813 589 2836
rect 578 2793 581 2806
rect 586 2726 589 2786
rect 594 2736 597 2946
rect 602 2813 605 2826
rect 618 2813 621 3033
rect 642 3026 645 3083
rect 654 3036 657 3113
rect 666 3083 669 3136
rect 654 3033 661 3036
rect 626 2986 629 3026
rect 634 3023 645 3026
rect 634 3006 637 3023
rect 658 3013 661 3033
rect 634 3003 645 3006
rect 626 2983 637 2986
rect 626 2923 629 2976
rect 634 2926 637 2983
rect 642 2933 645 3003
rect 650 2986 653 3006
rect 666 3003 669 3036
rect 674 3003 677 3126
rect 682 3053 685 3136
rect 730 3106 733 3366
rect 722 3103 733 3106
rect 722 3056 725 3103
rect 746 3096 749 3156
rect 762 3146 765 3440
rect 810 3406 813 3440
rect 774 3403 813 3406
rect 774 3346 777 3403
rect 834 3366 837 3440
rect 826 3363 837 3366
rect 850 3363 853 3440
rect 866 3426 869 3440
rect 866 3423 877 3426
rect 770 3343 777 3346
rect 770 3196 773 3343
rect 778 3203 781 3326
rect 770 3193 781 3196
rect 762 3143 773 3146
rect 770 3096 773 3143
rect 742 3093 749 3096
rect 762 3093 773 3096
rect 722 3053 733 3056
rect 650 2983 657 2986
rect 634 2923 645 2926
rect 642 2906 645 2923
rect 634 2903 645 2906
rect 634 2846 637 2903
rect 654 2876 657 2983
rect 666 2913 669 2926
rect 674 2923 677 2996
rect 682 2993 685 3016
rect 690 2936 693 3006
rect 698 2973 701 3016
rect 706 3013 709 3026
rect 722 3016 725 3036
rect 718 3013 725 3016
rect 682 2933 693 2936
rect 674 2896 677 2906
rect 682 2903 685 2933
rect 698 2923 701 2966
rect 690 2903 693 2916
rect 674 2893 693 2896
rect 650 2873 657 2876
rect 650 2853 653 2873
rect 634 2843 645 2846
rect 642 2813 645 2843
rect 658 2813 661 2836
rect 666 2813 669 2826
rect 634 2783 637 2806
rect 658 2786 661 2806
rect 682 2803 685 2826
rect 690 2813 693 2893
rect 706 2843 709 3006
rect 718 2956 721 3013
rect 730 2993 733 3053
rect 742 3016 745 3093
rect 742 3013 749 3016
rect 746 2993 749 3013
rect 714 2953 721 2956
rect 714 2916 717 2953
rect 746 2946 749 2956
rect 722 2943 749 2946
rect 722 2923 725 2943
rect 730 2923 733 2936
rect 738 2923 741 2936
rect 746 2933 749 2943
rect 714 2913 725 2916
rect 706 2813 709 2836
rect 722 2823 725 2913
rect 658 2783 665 2786
rect 618 2743 637 2746
rect 634 2736 637 2743
rect 594 2733 621 2736
rect 634 2733 645 2736
rect 546 2713 549 2726
rect 554 2723 597 2726
rect 610 2723 637 2726
rect 530 2623 541 2626
rect 530 2593 533 2623
rect 554 2616 557 2723
rect 610 2716 613 2723
rect 570 2713 613 2716
rect 538 2613 557 2616
rect 562 2613 565 2636
rect 538 2526 541 2613
rect 570 2606 573 2713
rect 642 2706 645 2733
rect 634 2703 645 2706
rect 610 2646 613 2666
rect 546 2603 573 2606
rect 554 2593 565 2596
rect 554 2533 557 2566
rect 578 2536 581 2606
rect 586 2586 589 2636
rect 594 2593 597 2646
rect 606 2643 613 2646
rect 586 2583 597 2586
rect 570 2533 581 2536
rect 570 2526 573 2533
rect 530 2523 541 2526
rect 498 2493 517 2496
rect 498 2403 501 2493
rect 506 2413 509 2426
rect 522 2413 525 2446
rect 546 2436 549 2526
rect 554 2523 573 2526
rect 554 2506 557 2523
rect 578 2513 581 2526
rect 554 2503 581 2506
rect 586 2453 589 2526
rect 530 2433 549 2436
rect 466 2363 473 2366
rect 458 2333 461 2346
rect 466 2266 469 2363
rect 514 2356 517 2406
rect 530 2393 533 2433
rect 538 2386 541 2426
rect 578 2413 581 2446
rect 594 2423 597 2583
rect 606 2536 609 2643
rect 618 2553 621 2646
rect 634 2626 637 2703
rect 626 2623 637 2626
rect 606 2533 613 2536
rect 610 2516 613 2533
rect 626 2523 629 2623
rect 602 2446 605 2516
rect 610 2513 629 2516
rect 602 2443 621 2446
rect 530 2383 541 2386
rect 546 2386 549 2406
rect 546 2383 553 2386
rect 506 2353 517 2356
rect 482 2313 485 2336
rect 386 2083 413 2086
rect 426 2233 433 2236
rect 442 2263 469 2266
rect 386 2056 389 2083
rect 386 2053 397 2056
rect 394 1976 397 2053
rect 274 1953 285 1956
rect 290 1963 301 1966
rect 314 1963 325 1966
rect 354 1963 365 1966
rect 386 1973 397 1976
rect 250 1933 253 1946
rect 258 1933 261 1946
rect 250 1913 253 1926
rect 226 1903 245 1906
rect 186 1873 197 1876
rect 174 1783 181 1786
rect 162 1763 169 1766
rect 90 1753 101 1756
rect 98 1656 101 1753
rect 146 1723 149 1746
rect 166 1686 169 1763
rect 66 1643 77 1646
rect 90 1653 101 1656
rect 162 1683 169 1686
rect 66 1576 69 1643
rect 66 1573 77 1576
rect 74 1446 77 1573
rect 66 1443 77 1446
rect 66 1296 69 1443
rect 66 1293 77 1296
rect 74 1136 77 1293
rect 90 1286 93 1653
rect 114 1533 117 1616
rect 162 1613 165 1683
rect 122 1533 125 1606
rect 170 1603 173 1616
rect 178 1576 181 1783
rect 186 1776 189 1873
rect 202 1813 205 1856
rect 194 1793 197 1806
rect 218 1803 221 1816
rect 186 1773 197 1776
rect 194 1666 197 1773
rect 218 1723 221 1786
rect 242 1776 245 1903
rect 274 1853 277 1953
rect 282 1933 285 1946
rect 290 1866 293 1963
rect 286 1863 293 1866
rect 258 1793 261 1816
rect 226 1773 245 1776
rect 186 1663 197 1666
rect 186 1586 189 1663
rect 202 1593 205 1606
rect 186 1583 197 1586
rect 178 1573 189 1576
rect 154 1543 181 1546
rect 146 1453 149 1536
rect 154 1523 157 1543
rect 162 1533 173 1536
rect 178 1493 181 1516
rect 186 1476 189 1573
rect 194 1556 197 1583
rect 226 1576 229 1773
rect 286 1766 289 1863
rect 286 1763 293 1766
rect 250 1733 253 1746
rect 282 1726 285 1746
rect 274 1723 285 1726
rect 250 1693 253 1716
rect 274 1666 277 1723
rect 274 1663 285 1666
rect 282 1623 285 1663
rect 218 1573 229 1576
rect 194 1553 205 1556
rect 202 1496 205 1553
rect 170 1473 189 1476
rect 194 1493 205 1496
rect 114 1393 117 1416
rect 114 1323 117 1346
rect 90 1283 101 1286
rect 98 1173 101 1283
rect 122 1246 125 1376
rect 170 1266 173 1473
rect 170 1263 181 1266
rect 122 1243 133 1246
rect 130 1196 133 1243
rect 122 1193 133 1196
rect 146 1193 149 1216
rect 122 1146 125 1193
rect 178 1186 181 1263
rect 194 1193 197 1493
rect 218 1476 221 1573
rect 210 1473 221 1476
rect 242 1476 245 1616
rect 250 1593 253 1616
rect 250 1503 253 1536
rect 242 1473 253 1476
rect 210 1296 213 1473
rect 234 1423 237 1436
rect 218 1413 237 1416
rect 234 1393 237 1406
rect 250 1356 253 1473
rect 266 1366 269 1536
rect 290 1533 293 1763
rect 290 1503 293 1526
rect 298 1496 301 1856
rect 314 1746 317 1963
rect 338 1923 341 1946
rect 338 1836 341 1916
rect 354 1886 357 1963
rect 354 1883 365 1886
rect 306 1743 317 1746
rect 330 1833 341 1836
rect 306 1706 309 1743
rect 314 1723 317 1736
rect 322 1713 325 1726
rect 306 1703 313 1706
rect 290 1493 301 1496
rect 274 1373 277 1416
rect 290 1413 293 1493
rect 310 1486 313 1703
rect 322 1613 325 1626
rect 330 1616 333 1833
rect 346 1803 349 1816
rect 338 1733 341 1746
rect 354 1733 357 1816
rect 362 1776 365 1883
rect 370 1793 373 1806
rect 362 1773 369 1776
rect 366 1726 369 1773
rect 378 1733 381 1906
rect 386 1813 389 1973
rect 402 1923 405 1956
rect 410 1906 413 1936
rect 418 1913 421 2006
rect 426 1943 429 2233
rect 434 2213 437 2226
rect 442 2193 445 2263
rect 458 2213 461 2236
rect 450 2183 453 2206
rect 466 2203 469 2256
rect 474 2213 477 2286
rect 482 2213 485 2246
rect 498 2213 501 2266
rect 450 2143 461 2146
rect 450 2133 453 2143
rect 434 2113 437 2126
rect 434 2003 437 2016
rect 442 2013 445 2126
rect 458 2103 461 2126
rect 458 2013 461 2036
rect 450 1993 453 2006
rect 466 2003 469 2156
rect 474 2133 477 2206
rect 474 2016 477 2126
rect 482 2106 485 2196
rect 490 2133 493 2206
rect 506 2203 509 2326
rect 514 2323 517 2346
rect 482 2103 489 2106
rect 486 2026 489 2103
rect 498 2093 501 2136
rect 486 2023 493 2026
rect 474 2013 485 2016
rect 426 1923 437 1926
rect 442 1923 445 1986
rect 450 1906 453 1966
rect 458 1933 461 1946
rect 466 1926 469 1976
rect 410 1903 437 1906
rect 394 1853 421 1856
rect 394 1823 397 1853
rect 402 1816 405 1846
rect 394 1813 405 1816
rect 418 1813 421 1853
rect 394 1796 397 1813
rect 390 1793 397 1796
rect 390 1736 393 1793
rect 410 1783 413 1806
rect 426 1803 429 1896
rect 434 1813 437 1903
rect 446 1903 453 1906
rect 458 1923 469 1926
rect 446 1836 449 1903
rect 446 1833 453 1836
rect 390 1733 397 1736
rect 346 1693 349 1726
rect 362 1723 369 1726
rect 362 1636 365 1723
rect 354 1633 365 1636
rect 354 1616 357 1633
rect 362 1623 389 1626
rect 330 1613 349 1616
rect 354 1613 365 1616
rect 322 1603 333 1606
rect 346 1586 349 1613
rect 354 1593 357 1606
rect 346 1583 357 1586
rect 354 1533 357 1583
rect 362 1503 365 1613
rect 370 1543 373 1616
rect 386 1613 389 1623
rect 378 1593 381 1606
rect 394 1603 397 1733
rect 402 1566 405 1776
rect 410 1603 413 1736
rect 418 1723 421 1796
rect 402 1563 413 1566
rect 394 1533 397 1546
rect 410 1526 413 1563
rect 418 1533 421 1636
rect 426 1613 429 1786
rect 450 1773 453 1833
rect 458 1793 461 1923
rect 474 1886 477 2006
rect 482 1963 485 2013
rect 466 1883 477 1886
rect 466 1726 469 1883
rect 482 1876 485 1946
rect 474 1873 485 1876
rect 474 1743 477 1873
rect 490 1853 493 2023
rect 498 1903 501 2026
rect 506 2003 509 2126
rect 514 2103 517 2236
rect 522 2203 525 2356
rect 530 2276 533 2383
rect 538 2373 541 2383
rect 550 2286 553 2383
rect 602 2336 605 2426
rect 618 2403 621 2443
rect 626 2343 629 2513
rect 634 2443 637 2606
rect 642 2593 645 2616
rect 650 2613 653 2766
rect 662 2666 665 2783
rect 674 2723 677 2776
rect 690 2723 693 2796
rect 658 2663 665 2666
rect 698 2663 701 2806
rect 722 2766 725 2786
rect 714 2763 725 2766
rect 658 2643 661 2663
rect 706 2653 709 2726
rect 714 2723 717 2763
rect 738 2746 741 2826
rect 746 2773 749 2876
rect 754 2783 757 3086
rect 762 2996 765 3093
rect 778 3083 781 3193
rect 770 3013 773 3056
rect 762 2993 769 2996
rect 766 2896 769 2993
rect 778 2923 781 3006
rect 786 2903 789 3286
rect 794 3153 797 3346
rect 826 3316 829 3363
rect 874 3356 877 3423
rect 842 3323 845 3356
rect 866 3353 877 3356
rect 866 3336 869 3353
rect 862 3333 869 3336
rect 882 3333 901 3336
rect 906 3333 909 3356
rect 922 3333 925 3346
rect 826 3313 837 3316
rect 802 3183 805 3216
rect 810 3213 813 3296
rect 834 3283 837 3313
rect 862 3256 865 3333
rect 862 3253 869 3256
rect 826 3213 845 3216
rect 850 3213 853 3226
rect 858 3213 861 3236
rect 794 3123 797 3146
rect 810 3066 813 3206
rect 834 3136 837 3206
rect 842 3186 845 3213
rect 866 3206 869 3253
rect 874 3223 877 3326
rect 882 3213 885 3316
rect 890 3213 893 3326
rect 858 3203 869 3206
rect 842 3183 849 3186
rect 794 3063 813 3066
rect 818 3133 837 3136
rect 794 3003 797 3063
rect 802 3013 805 3056
rect 810 3013 813 3046
rect 818 3026 821 3133
rect 826 3053 829 3126
rect 834 3063 837 3126
rect 818 3023 837 3026
rect 818 3013 829 3016
rect 762 2893 769 2896
rect 762 2873 765 2893
rect 802 2846 805 2996
rect 794 2843 805 2846
rect 762 2833 773 2836
rect 770 2753 773 2826
rect 786 2813 789 2826
rect 778 2763 781 2806
rect 738 2743 745 2746
rect 682 2643 717 2646
rect 682 2636 685 2643
rect 666 2633 685 2636
rect 658 2583 661 2616
rect 666 2613 669 2633
rect 674 2593 677 2606
rect 682 2556 685 2616
rect 690 2583 693 2636
rect 714 2623 717 2643
rect 642 2553 685 2556
rect 642 2496 645 2553
rect 698 2546 701 2616
rect 706 2603 717 2606
rect 722 2593 725 2736
rect 730 2603 733 2736
rect 742 2656 745 2743
rect 754 2703 757 2726
rect 762 2723 765 2736
rect 770 2706 773 2726
rect 766 2703 773 2706
rect 738 2653 745 2656
rect 738 2613 741 2653
rect 766 2636 769 2703
rect 746 2633 769 2636
rect 778 2633 781 2736
rect 794 2673 797 2843
rect 802 2813 805 2836
rect 810 2736 813 2806
rect 802 2733 813 2736
rect 810 2693 813 2726
rect 706 2553 717 2556
rect 650 2543 693 2546
rect 698 2543 733 2546
rect 650 2533 653 2543
rect 650 2513 669 2516
rect 642 2493 653 2496
rect 562 2323 565 2336
rect 546 2283 553 2286
rect 530 2273 537 2276
rect 534 2216 537 2273
rect 530 2213 537 2216
rect 530 2196 533 2213
rect 522 2193 533 2196
rect 522 2106 525 2193
rect 546 2123 549 2283
rect 570 2243 573 2326
rect 586 2266 589 2336
rect 602 2333 613 2336
rect 594 2303 597 2326
rect 586 2263 597 2266
rect 562 2223 589 2226
rect 562 2123 565 2223
rect 578 2186 581 2216
rect 586 2213 589 2223
rect 594 2216 597 2263
rect 602 2223 605 2246
rect 594 2213 605 2216
rect 610 2213 613 2333
rect 618 2233 621 2326
rect 626 2213 629 2246
rect 634 2213 637 2416
rect 642 2373 645 2416
rect 650 2353 653 2493
rect 674 2456 677 2536
rect 690 2513 693 2536
rect 714 2533 733 2536
rect 714 2503 717 2533
rect 738 2513 741 2566
rect 746 2456 749 2633
rect 754 2623 805 2626
rect 754 2613 757 2623
rect 674 2453 685 2456
rect 674 2423 677 2446
rect 682 2416 685 2453
rect 730 2453 749 2456
rect 674 2413 685 2416
rect 650 2326 653 2346
rect 658 2333 661 2366
rect 642 2233 645 2326
rect 650 2323 661 2326
rect 658 2303 661 2316
rect 650 2233 653 2256
rect 658 2216 661 2236
rect 602 2203 605 2213
rect 578 2183 585 2186
rect 570 2123 573 2176
rect 582 2126 585 2183
rect 594 2173 605 2176
rect 594 2133 597 2146
rect 602 2133 605 2173
rect 582 2123 605 2126
rect 610 2123 613 2206
rect 626 2203 637 2206
rect 626 2133 629 2203
rect 642 2146 645 2216
rect 650 2203 653 2216
rect 658 2213 665 2216
rect 662 2156 665 2213
rect 674 2173 677 2413
rect 682 2303 685 2326
rect 690 2286 693 2406
rect 698 2333 701 2406
rect 722 2376 725 2416
rect 730 2396 733 2453
rect 738 2423 741 2446
rect 738 2403 741 2416
rect 754 2413 757 2606
rect 762 2593 765 2606
rect 770 2583 773 2606
rect 778 2573 781 2616
rect 786 2606 789 2616
rect 810 2613 813 2626
rect 786 2603 813 2606
rect 818 2603 821 2856
rect 834 2826 837 3023
rect 846 2996 849 3183
rect 858 3116 861 3203
rect 898 3196 901 3333
rect 906 3313 909 3326
rect 954 3306 957 3326
rect 950 3303 957 3306
rect 950 3236 953 3303
rect 950 3233 957 3236
rect 962 3233 965 3440
rect 1018 3333 1021 3346
rect 1002 3276 1005 3326
rect 1066 3323 1069 3336
rect 1082 3333 1109 3336
rect 1138 3333 1149 3336
rect 994 3273 1005 3276
rect 866 3193 901 3196
rect 906 3223 941 3226
rect 866 3133 869 3193
rect 890 3133 893 3146
rect 858 3113 869 3116
rect 890 3113 893 3126
rect 898 3123 901 3186
rect 866 3056 869 3113
rect 858 3053 869 3056
rect 858 3033 861 3053
rect 906 3046 909 3223
rect 922 3176 925 3216
rect 930 3183 933 3206
rect 938 3203 941 3223
rect 954 3213 957 3233
rect 994 3226 997 3273
rect 962 3223 997 3226
rect 962 3213 965 3223
rect 970 3203 973 3216
rect 986 3213 1005 3216
rect 1018 3213 1021 3296
rect 922 3173 941 3176
rect 914 3103 917 3126
rect 922 3056 925 3156
rect 930 3123 933 3146
rect 938 3133 941 3173
rect 994 3153 997 3206
rect 1002 3183 1005 3213
rect 1026 3176 1029 3196
rect 1034 3186 1037 3216
rect 1042 3193 1045 3206
rect 1034 3183 1045 3186
rect 1022 3173 1029 3176
rect 978 3096 981 3126
rect 970 3093 981 3096
rect 922 3053 929 3056
rect 906 3043 917 3046
rect 874 3013 877 3026
rect 842 2993 849 2996
rect 890 2993 893 3006
rect 842 2973 845 2993
rect 914 2956 917 3043
rect 850 2923 853 2946
rect 882 2923 885 2936
rect 890 2906 893 2936
rect 898 2923 901 2956
rect 906 2953 917 2956
rect 906 2916 909 2953
rect 926 2946 929 3053
rect 970 3046 973 3093
rect 970 3043 981 3046
rect 938 2993 941 3016
rect 970 3013 973 3026
rect 978 2996 981 3043
rect 974 2993 981 2996
rect 914 2933 917 2946
rect 922 2943 929 2946
rect 922 2926 925 2943
rect 882 2903 893 2906
rect 898 2913 909 2916
rect 914 2923 925 2926
rect 826 2823 837 2826
rect 826 2773 829 2823
rect 786 2566 789 2603
rect 778 2563 789 2566
rect 762 2453 765 2546
rect 770 2446 773 2556
rect 778 2523 781 2563
rect 786 2523 789 2546
rect 762 2443 773 2446
rect 730 2393 741 2396
rect 714 2356 717 2376
rect 722 2373 729 2376
rect 710 2353 717 2356
rect 686 2283 693 2286
rect 686 2226 689 2283
rect 682 2223 689 2226
rect 682 2203 685 2223
rect 662 2153 669 2156
rect 642 2143 653 2146
rect 578 2113 597 2116
rect 522 2103 533 2106
rect 530 2046 533 2103
rect 514 2043 533 2046
rect 514 1996 517 2043
rect 506 1993 517 1996
rect 482 1833 501 1836
rect 482 1803 485 1833
rect 490 1813 493 1826
rect 498 1783 501 1826
rect 506 1813 509 1993
rect 522 1973 525 2026
rect 530 2003 533 2026
rect 538 1996 541 2016
rect 570 2013 573 2026
rect 538 1993 549 1996
rect 546 1946 549 1993
rect 538 1943 549 1946
rect 522 1933 533 1936
rect 522 1913 525 1933
rect 538 1906 541 1943
rect 530 1903 541 1906
rect 514 1736 517 1856
rect 530 1846 533 1903
rect 526 1843 533 1846
rect 526 1766 529 1843
rect 522 1763 529 1766
rect 522 1743 525 1763
rect 538 1736 541 1826
rect 546 1746 549 1826
rect 554 1803 557 1926
rect 562 1896 565 1926
rect 570 1913 573 1946
rect 578 1923 581 2113
rect 602 2033 605 2123
rect 618 2026 621 2116
rect 594 2023 621 2026
rect 562 1893 573 1896
rect 570 1806 573 1893
rect 562 1803 573 1806
rect 562 1786 565 1803
rect 586 1793 589 2006
rect 594 2003 597 2023
rect 626 2016 629 2036
rect 634 2023 637 2126
rect 602 1983 605 2016
rect 618 2013 629 2016
rect 594 1813 597 1836
rect 562 1783 581 1786
rect 546 1743 565 1746
rect 434 1706 437 1726
rect 450 1723 469 1726
rect 434 1703 445 1706
rect 450 1703 453 1716
rect 458 1666 461 1723
rect 474 1706 477 1736
rect 506 1716 509 1736
rect 514 1733 525 1736
rect 450 1663 461 1666
rect 470 1703 477 1706
rect 450 1613 453 1663
rect 470 1646 473 1703
rect 470 1643 477 1646
rect 466 1616 469 1626
rect 458 1613 469 1616
rect 306 1483 313 1486
rect 282 1366 285 1396
rect 290 1376 293 1406
rect 306 1393 309 1483
rect 378 1443 381 1526
rect 386 1486 389 1526
rect 394 1523 405 1526
rect 410 1523 421 1526
rect 394 1493 397 1523
rect 402 1496 405 1516
rect 402 1493 409 1496
rect 386 1483 397 1486
rect 394 1426 397 1483
rect 386 1423 397 1426
rect 330 1376 333 1416
rect 386 1406 389 1423
rect 290 1373 333 1376
rect 378 1403 389 1406
rect 266 1363 293 1366
rect 250 1353 261 1356
rect 234 1333 237 1346
rect 218 1323 237 1326
rect 226 1313 237 1316
rect 258 1296 261 1353
rect 274 1333 277 1346
rect 210 1293 221 1296
rect 258 1293 277 1296
rect 218 1226 221 1293
rect 210 1223 221 1226
rect 258 1223 261 1256
rect 274 1236 277 1293
rect 290 1236 293 1363
rect 378 1356 381 1403
rect 394 1363 397 1416
rect 406 1366 409 1493
rect 418 1433 421 1523
rect 426 1496 429 1586
rect 434 1533 437 1566
rect 442 1513 445 1526
rect 458 1523 461 1613
rect 466 1516 469 1606
rect 474 1593 477 1643
rect 482 1606 485 1716
rect 498 1713 509 1716
rect 498 1666 501 1713
rect 498 1663 509 1666
rect 490 1613 493 1626
rect 498 1623 501 1646
rect 506 1633 509 1663
rect 482 1603 501 1606
rect 506 1603 509 1626
rect 450 1513 469 1516
rect 426 1493 437 1496
rect 426 1413 429 1426
rect 418 1373 421 1406
rect 434 1403 437 1493
rect 406 1363 429 1366
rect 378 1353 389 1356
rect 322 1323 325 1346
rect 378 1316 381 1336
rect 386 1323 389 1353
rect 410 1333 413 1346
rect 426 1333 429 1363
rect 442 1333 445 1436
rect 450 1403 453 1513
rect 458 1413 461 1506
rect 474 1416 477 1426
rect 466 1413 477 1416
rect 482 1413 485 1536
rect 490 1523 493 1576
rect 370 1313 381 1316
rect 274 1233 285 1236
rect 290 1233 333 1236
rect 210 1206 213 1223
rect 242 1213 269 1216
rect 210 1203 237 1206
rect 178 1183 189 1186
rect 66 1133 77 1136
rect 98 1133 101 1146
rect 122 1143 133 1146
rect 66 693 69 1133
rect 74 1096 77 1116
rect 130 1096 133 1143
rect 178 1126 181 1146
rect 74 1093 85 1096
rect 82 966 85 1093
rect 122 1093 133 1096
rect 122 1016 125 1093
rect 146 1076 149 1126
rect 170 1123 181 1126
rect 146 1073 157 1076
rect 122 1013 133 1016
rect 98 993 101 1006
rect 114 993 117 1006
rect 74 963 85 966
rect 74 896 77 963
rect 74 893 81 896
rect 78 756 81 893
rect 90 836 93 946
rect 90 833 109 836
rect 74 753 81 756
rect 74 696 77 753
rect 82 723 85 736
rect 90 713 93 796
rect 74 693 85 696
rect 82 636 85 693
rect 74 633 85 636
rect 74 496 77 633
rect 106 616 109 833
rect 122 813 125 1013
rect 138 1003 141 1066
rect 146 1003 149 1016
rect 154 996 157 1073
rect 170 1046 173 1123
rect 170 1043 181 1046
rect 162 1013 165 1026
rect 130 993 157 996
rect 162 966 165 1006
rect 138 963 165 966
rect 138 923 141 963
rect 170 923 173 996
rect 178 916 181 1043
rect 170 913 181 916
rect 154 776 157 806
rect 170 803 173 913
rect 186 883 189 1183
rect 210 1133 213 1146
rect 194 1093 197 1126
rect 234 1063 237 1203
rect 258 1183 261 1206
rect 266 1193 269 1213
rect 282 1186 285 1233
rect 306 1203 309 1226
rect 330 1203 333 1233
rect 354 1213 357 1226
rect 282 1183 293 1186
rect 242 1056 245 1126
rect 290 1086 293 1183
rect 370 1176 373 1313
rect 394 1283 397 1326
rect 418 1313 421 1326
rect 434 1323 445 1326
rect 314 1123 317 1136
rect 338 1133 341 1176
rect 370 1173 381 1176
rect 378 1136 381 1173
rect 282 1083 293 1086
rect 194 1036 197 1056
rect 234 1053 245 1056
rect 194 1033 201 1036
rect 198 966 201 1033
rect 210 993 213 1006
rect 226 993 229 1006
rect 234 1003 237 1053
rect 242 1013 245 1026
rect 250 986 253 1066
rect 258 1003 261 1016
rect 194 963 201 966
rect 242 983 253 986
rect 194 876 197 963
rect 210 933 213 946
rect 242 916 245 983
rect 274 976 277 1006
rect 258 973 277 976
rect 258 923 261 973
rect 242 913 253 916
rect 194 873 205 876
rect 194 776 197 816
rect 202 806 205 873
rect 202 803 213 806
rect 154 773 197 776
rect 210 756 213 803
rect 202 753 213 756
rect 154 723 157 736
rect 178 723 189 726
rect 194 713 197 726
rect 202 616 205 753
rect 210 713 213 736
rect 218 733 229 736
rect 234 723 237 896
rect 234 616 237 626
rect 90 613 109 616
rect 90 566 93 613
rect 106 583 109 606
rect 90 563 101 566
rect 98 523 101 563
rect 114 553 117 616
rect 122 613 133 616
rect 138 613 149 616
rect 154 613 165 616
rect 202 613 237 616
rect 122 523 125 606
rect 138 603 141 613
rect 154 606 157 613
rect 146 603 157 606
rect 146 583 149 603
rect 210 596 213 613
rect 218 603 237 606
rect 202 593 213 596
rect 202 536 205 593
rect 218 543 221 556
rect 202 533 213 536
rect 74 493 85 496
rect 82 436 85 493
rect 74 433 85 436
rect 74 413 77 433
rect 90 413 101 416
rect 90 403 93 413
rect 114 376 117 406
rect 162 403 165 526
rect 210 433 213 533
rect 234 523 237 596
rect 242 443 245 886
rect 250 876 253 913
rect 250 873 261 876
rect 258 806 261 873
rect 282 826 285 1083
rect 322 1046 325 1126
rect 346 1053 349 1136
rect 354 1133 381 1136
rect 354 1123 357 1133
rect 378 1083 381 1126
rect 386 1116 389 1126
rect 394 1123 405 1126
rect 386 1113 401 1116
rect 298 1023 309 1026
rect 290 923 293 996
rect 298 953 301 1006
rect 306 943 309 1016
rect 314 923 317 1046
rect 322 1043 349 1046
rect 322 1013 333 1016
rect 338 1013 341 1036
rect 322 1003 333 1006
rect 330 933 333 1003
rect 338 993 341 1006
rect 346 913 349 1043
rect 362 1013 365 1026
rect 386 1023 389 1106
rect 398 1036 401 1113
rect 398 1033 405 1036
rect 370 1013 397 1016
rect 370 1006 373 1013
rect 354 953 357 1006
rect 362 1003 373 1006
rect 378 993 381 1006
rect 386 986 389 1006
rect 362 983 389 986
rect 354 933 357 946
rect 362 943 365 983
rect 394 946 397 1013
rect 402 963 405 1033
rect 370 933 373 946
rect 394 943 405 946
rect 394 933 397 943
rect 274 823 285 826
rect 274 806 277 823
rect 298 816 301 826
rect 250 803 261 806
rect 270 803 277 806
rect 250 783 253 803
rect 270 746 273 803
rect 282 773 285 816
rect 298 813 309 816
rect 290 793 293 806
rect 298 756 301 813
rect 306 793 309 806
rect 314 803 317 846
rect 322 803 325 816
rect 354 813 357 826
rect 330 783 333 806
rect 338 803 349 806
rect 294 753 301 756
rect 270 743 277 746
rect 250 733 261 736
rect 250 713 253 726
rect 258 696 261 733
rect 274 726 277 743
rect 274 723 285 726
rect 254 693 261 696
rect 254 626 257 693
rect 250 623 257 626
rect 250 603 253 623
rect 266 616 269 716
rect 282 616 285 723
rect 294 706 297 753
rect 294 703 301 706
rect 258 613 269 616
rect 274 613 285 616
rect 258 576 261 613
rect 274 593 277 613
rect 298 586 301 703
rect 298 583 309 586
rect 250 573 261 576
rect 250 496 253 573
rect 258 563 301 566
rect 258 533 261 563
rect 274 533 277 546
rect 298 523 301 563
rect 306 533 309 583
rect 250 493 261 496
rect 258 436 261 493
rect 250 433 261 436
rect 210 393 213 416
rect 250 403 253 433
rect 298 403 301 416
rect 306 413 309 426
rect 314 383 317 766
rect 338 723 341 803
rect 354 686 357 706
rect 346 683 357 686
rect 346 636 349 683
rect 346 633 357 636
rect 354 613 357 633
rect 362 613 365 926
rect 370 816 373 916
rect 378 823 381 926
rect 410 913 413 1266
rect 426 1203 429 1246
rect 434 1183 437 1323
rect 450 1303 453 1336
rect 450 1246 453 1276
rect 458 1253 461 1326
rect 442 1243 461 1246
rect 442 1206 445 1243
rect 450 1213 453 1226
rect 458 1213 461 1243
rect 466 1213 469 1413
rect 474 1333 477 1406
rect 482 1263 485 1406
rect 490 1323 493 1386
rect 498 1306 501 1603
rect 506 1533 509 1566
rect 514 1513 517 1726
rect 522 1686 525 1733
rect 530 1696 533 1736
rect 538 1733 557 1736
rect 530 1693 541 1696
rect 522 1683 533 1686
rect 522 1613 525 1666
rect 506 1466 509 1486
rect 506 1463 513 1466
rect 510 1376 513 1463
rect 506 1373 513 1376
rect 506 1333 509 1373
rect 494 1303 501 1306
rect 482 1223 485 1246
rect 494 1226 497 1303
rect 494 1223 501 1226
rect 474 1213 485 1216
rect 474 1206 477 1213
rect 498 1206 501 1223
rect 442 1203 453 1206
rect 418 1083 421 1126
rect 418 923 421 1076
rect 426 973 429 1136
rect 434 1073 437 1126
rect 442 1043 445 1136
rect 442 1016 445 1026
rect 434 1013 445 1016
rect 434 953 437 1013
rect 442 936 445 1006
rect 450 993 453 1203
rect 450 943 453 956
rect 442 933 453 936
rect 458 933 461 1206
rect 466 1203 477 1206
rect 490 1203 501 1206
rect 466 1023 469 1186
rect 474 1113 477 1203
rect 506 1196 509 1326
rect 514 1313 517 1356
rect 522 1333 525 1606
rect 530 1423 533 1683
rect 538 1643 541 1693
rect 538 1506 541 1626
rect 546 1573 549 1726
rect 554 1563 557 1733
rect 562 1523 565 1743
rect 538 1503 549 1506
rect 570 1503 573 1776
rect 578 1663 581 1783
rect 594 1746 597 1806
rect 586 1743 597 1746
rect 586 1666 589 1743
rect 602 1713 605 1806
rect 610 1753 613 1946
rect 618 1893 621 2013
rect 634 1943 637 2006
rect 642 1933 645 2136
rect 650 2126 653 2143
rect 650 2123 657 2126
rect 654 2066 657 2123
rect 650 2063 657 2066
rect 650 2033 653 2063
rect 666 2046 669 2153
rect 690 2123 693 2216
rect 698 2126 701 2326
rect 710 2306 713 2353
rect 710 2303 717 2306
rect 706 2206 709 2236
rect 714 2223 717 2303
rect 726 2236 729 2373
rect 738 2253 741 2393
rect 746 2343 749 2406
rect 746 2246 749 2326
rect 754 2296 757 2356
rect 762 2323 765 2443
rect 778 2426 781 2446
rect 794 2443 797 2576
rect 802 2506 805 2566
rect 810 2523 813 2603
rect 818 2533 821 2596
rect 802 2503 809 2506
rect 770 2423 781 2426
rect 770 2413 773 2423
rect 778 2413 789 2416
rect 794 2413 797 2436
rect 806 2426 809 2503
rect 802 2423 809 2426
rect 770 2333 773 2406
rect 778 2353 781 2413
rect 786 2376 789 2406
rect 802 2403 805 2423
rect 786 2373 797 2376
rect 778 2323 781 2346
rect 794 2333 797 2373
rect 762 2303 765 2316
rect 786 2303 789 2326
rect 754 2293 773 2296
rect 746 2243 757 2246
rect 726 2233 733 2236
rect 730 2213 733 2233
rect 706 2203 725 2206
rect 714 2193 725 2196
rect 706 2133 717 2136
rect 722 2133 725 2146
rect 698 2123 717 2126
rect 658 2043 669 2046
rect 650 2006 653 2016
rect 658 2013 661 2043
rect 666 2023 693 2026
rect 650 2003 661 2006
rect 650 1933 653 1946
rect 610 1723 613 1736
rect 618 1733 621 1816
rect 626 1793 629 1916
rect 586 1663 593 1666
rect 578 1603 581 1616
rect 590 1596 593 1663
rect 626 1656 629 1726
rect 634 1696 637 1896
rect 642 1833 645 1926
rect 650 1773 653 1926
rect 658 1886 661 2003
rect 666 1923 669 2023
rect 698 1993 701 2006
rect 706 2003 709 2036
rect 714 2016 717 2123
rect 722 2093 725 2126
rect 730 2123 733 2166
rect 738 2143 741 2236
rect 746 2213 749 2226
rect 746 2133 749 2186
rect 754 2163 757 2243
rect 730 2113 749 2116
rect 754 2113 757 2126
rect 714 2013 725 2016
rect 674 1933 677 1966
rect 682 1933 685 1946
rect 714 1936 717 2013
rect 658 1883 669 1886
rect 666 1836 669 1883
rect 662 1833 669 1836
rect 662 1756 665 1833
rect 674 1783 677 1816
rect 642 1733 645 1746
rect 650 1733 653 1756
rect 658 1753 665 1756
rect 658 1726 661 1753
rect 666 1733 677 1736
rect 650 1723 661 1726
rect 666 1723 677 1726
rect 642 1703 645 1716
rect 674 1703 677 1723
rect 682 1696 685 1926
rect 690 1823 693 1836
rect 690 1803 693 1816
rect 698 1813 701 1936
rect 706 1933 717 1936
rect 706 1923 709 1933
rect 714 1906 717 1926
rect 730 1923 733 2113
rect 754 2076 757 2096
rect 746 2073 757 2076
rect 746 2006 749 2073
rect 762 2016 765 2286
rect 770 2186 773 2293
rect 802 2283 805 2326
rect 810 2323 813 2336
rect 818 2323 821 2446
rect 778 2203 781 2246
rect 770 2183 777 2186
rect 774 2046 777 2183
rect 786 2163 789 2216
rect 810 2213 813 2236
rect 818 2213 821 2256
rect 794 2173 797 2206
rect 810 2196 813 2206
rect 770 2043 777 2046
rect 770 2026 773 2043
rect 786 2033 789 2146
rect 770 2023 781 2026
rect 762 2013 773 2016
rect 746 2003 765 2006
rect 738 1933 741 1966
rect 762 1946 765 2003
rect 778 1976 781 2023
rect 786 1983 789 2026
rect 794 1993 797 2136
rect 802 2103 805 2196
rect 810 2193 821 2196
rect 810 2133 813 2176
rect 818 2163 821 2193
rect 818 2133 821 2146
rect 810 2016 813 2036
rect 818 2023 821 2126
rect 826 2026 829 2756
rect 834 2753 837 2816
rect 842 2746 845 2816
rect 858 2803 861 2866
rect 882 2836 885 2903
rect 882 2833 893 2836
rect 866 2793 869 2826
rect 882 2763 885 2816
rect 890 2753 893 2833
rect 898 2786 901 2913
rect 914 2833 917 2923
rect 922 2826 925 2916
rect 930 2873 933 2916
rect 946 2866 949 2966
rect 974 2916 977 2993
rect 974 2913 981 2916
rect 978 2893 981 2913
rect 986 2876 989 3006
rect 994 2963 997 3136
rect 1022 3036 1025 3173
rect 1034 3123 1037 3156
rect 1042 3116 1045 3183
rect 1050 3173 1053 3216
rect 1082 3206 1085 3333
rect 1098 3293 1101 3326
rect 1114 3256 1117 3326
rect 1138 3313 1149 3316
rect 1154 3296 1157 3326
rect 1106 3253 1117 3256
rect 1146 3293 1157 3296
rect 1074 3203 1085 3206
rect 1074 3123 1077 3146
rect 1082 3133 1085 3203
rect 1090 3166 1093 3236
rect 1098 3203 1101 3216
rect 1106 3183 1109 3253
rect 1114 3166 1117 3226
rect 1090 3163 1101 3166
rect 1034 3113 1045 3116
rect 1022 3033 1029 3036
rect 1026 3016 1029 3033
rect 1034 3023 1037 3113
rect 1042 3023 1053 3026
rect 1018 2953 1021 3016
rect 1026 3013 1037 3016
rect 1026 2996 1029 3013
rect 1042 3006 1045 3016
rect 1034 3003 1045 3006
rect 1026 2993 1037 2996
rect 994 2923 997 2946
rect 1034 2936 1037 2993
rect 1050 2983 1053 3023
rect 1066 2993 1069 3006
rect 1074 2966 1077 3116
rect 1082 3103 1085 3126
rect 1098 3096 1101 3163
rect 1090 3093 1101 3096
rect 1110 3163 1117 3166
rect 1110 3096 1113 3163
rect 1122 3133 1125 3156
rect 1110 3093 1117 3096
rect 1018 2933 1037 2936
rect 1018 2876 1021 2933
rect 986 2873 997 2876
rect 946 2863 965 2866
rect 906 2823 941 2826
rect 906 2803 909 2823
rect 922 2803 925 2816
rect 938 2813 941 2823
rect 930 2786 933 2806
rect 898 2783 933 2786
rect 922 2766 925 2783
rect 914 2763 925 2766
rect 834 2723 837 2746
rect 842 2743 885 2746
rect 834 2703 837 2716
rect 850 2706 853 2736
rect 866 2723 869 2743
rect 882 2736 885 2743
rect 850 2703 861 2706
rect 834 2563 837 2636
rect 842 2626 845 2696
rect 858 2656 861 2703
rect 874 2666 877 2736
rect 882 2733 893 2736
rect 890 2703 893 2726
rect 874 2663 893 2666
rect 850 2653 861 2656
rect 850 2633 853 2653
rect 842 2623 869 2626
rect 842 2613 845 2623
rect 834 2533 837 2546
rect 850 2536 853 2606
rect 858 2603 861 2616
rect 866 2593 869 2623
rect 874 2553 877 2616
rect 882 2536 885 2656
rect 890 2583 893 2663
rect 898 2613 901 2726
rect 914 2676 917 2763
rect 914 2673 925 2676
rect 922 2653 925 2673
rect 930 2646 933 2776
rect 946 2756 949 2836
rect 962 2776 965 2863
rect 938 2753 949 2756
rect 954 2773 965 2776
rect 938 2723 941 2753
rect 914 2576 917 2646
rect 930 2643 941 2646
rect 850 2533 861 2536
rect 834 2513 837 2526
rect 842 2493 845 2526
rect 858 2456 861 2533
rect 834 2333 837 2406
rect 842 2393 845 2456
rect 850 2453 861 2456
rect 874 2533 885 2536
rect 898 2573 925 2576
rect 898 2533 901 2573
rect 922 2556 925 2573
rect 922 2553 929 2556
rect 874 2456 877 2533
rect 890 2486 893 2506
rect 926 2496 929 2553
rect 938 2503 941 2643
rect 946 2626 949 2656
rect 954 2643 957 2773
rect 946 2623 953 2626
rect 950 2566 953 2623
rect 962 2613 965 2626
rect 950 2563 965 2566
rect 946 2523 949 2546
rect 922 2493 929 2496
rect 890 2483 897 2486
rect 874 2453 885 2456
rect 850 2333 853 2453
rect 866 2413 869 2436
rect 874 2413 877 2426
rect 882 2406 885 2453
rect 858 2393 861 2406
rect 874 2403 885 2406
rect 858 2326 861 2336
rect 834 2093 837 2326
rect 842 2323 861 2326
rect 842 2213 845 2323
rect 866 2313 869 2326
rect 874 2303 877 2403
rect 894 2396 897 2483
rect 890 2393 897 2396
rect 850 2126 853 2246
rect 866 2203 869 2296
rect 882 2243 885 2346
rect 890 2176 893 2393
rect 850 2123 857 2126
rect 826 2023 837 2026
rect 802 2003 805 2016
rect 810 2013 821 2016
rect 834 2013 837 2023
rect 842 2013 845 2116
rect 818 1976 821 2006
rect 826 1983 829 2006
rect 778 1973 789 1976
rect 818 1973 829 1976
rect 746 1933 749 1946
rect 762 1943 773 1946
rect 714 1903 725 1906
rect 746 1903 749 1926
rect 706 1816 709 1836
rect 706 1813 717 1816
rect 634 1693 645 1696
rect 626 1653 637 1656
rect 602 1643 629 1646
rect 602 1623 605 1643
rect 602 1603 605 1616
rect 610 1613 613 1636
rect 626 1613 629 1643
rect 590 1593 597 1596
rect 546 1436 549 1503
rect 578 1496 581 1536
rect 586 1523 589 1576
rect 594 1513 597 1593
rect 618 1573 621 1606
rect 602 1533 629 1536
rect 578 1493 589 1496
rect 538 1433 549 1436
rect 586 1436 589 1493
rect 586 1433 597 1436
rect 538 1393 541 1433
rect 530 1326 533 1336
rect 522 1323 533 1326
rect 522 1296 525 1323
rect 498 1193 509 1196
rect 518 1293 525 1296
rect 482 1113 485 1146
rect 490 1103 493 1126
rect 474 1023 493 1026
rect 466 1003 469 1016
rect 474 1013 477 1023
rect 482 1003 485 1016
rect 466 986 469 996
rect 490 993 493 1023
rect 498 986 501 1193
rect 466 983 501 986
rect 442 893 445 926
rect 450 896 453 933
rect 450 893 461 896
rect 458 866 461 893
rect 450 863 461 866
rect 466 863 469 983
rect 506 963 509 1186
rect 518 1166 521 1293
rect 530 1273 533 1316
rect 538 1226 541 1336
rect 546 1323 549 1416
rect 554 1356 557 1416
rect 562 1403 565 1416
rect 570 1393 573 1416
rect 586 1383 589 1406
rect 554 1353 589 1356
rect 554 1333 557 1353
rect 530 1223 541 1226
rect 518 1163 525 1166
rect 522 1143 525 1163
rect 530 1136 533 1223
rect 546 1216 549 1256
rect 514 1133 533 1136
rect 538 1213 549 1216
rect 554 1213 557 1276
rect 562 1263 565 1326
rect 570 1303 573 1336
rect 578 1333 581 1346
rect 586 1333 589 1353
rect 594 1316 597 1433
rect 538 1133 541 1213
rect 514 1003 517 1133
rect 522 1073 525 1116
rect 530 1056 533 1126
rect 546 1123 549 1186
rect 522 1053 533 1056
rect 514 956 517 996
rect 522 973 525 1053
rect 554 1026 557 1176
rect 570 1136 573 1206
rect 578 1183 581 1316
rect 590 1313 597 1316
rect 590 1216 593 1313
rect 602 1253 605 1533
rect 610 1266 613 1526
rect 618 1523 629 1526
rect 618 1353 621 1523
rect 626 1503 629 1516
rect 626 1343 629 1406
rect 618 1333 629 1336
rect 634 1333 637 1653
rect 642 1633 645 1693
rect 666 1693 685 1696
rect 642 1523 645 1606
rect 650 1536 653 1666
rect 666 1613 669 1693
rect 690 1686 693 1796
rect 674 1683 693 1686
rect 674 1596 677 1683
rect 698 1676 701 1806
rect 682 1673 701 1676
rect 682 1606 685 1673
rect 690 1613 701 1616
rect 682 1603 693 1606
rect 698 1596 701 1606
rect 674 1593 701 1596
rect 650 1533 661 1536
rect 650 1513 653 1526
rect 658 1506 661 1533
rect 666 1513 669 1556
rect 650 1503 661 1506
rect 650 1413 653 1503
rect 658 1413 661 1426
rect 650 1356 653 1406
rect 642 1353 653 1356
rect 642 1333 645 1353
rect 626 1326 629 1333
rect 618 1293 621 1326
rect 626 1323 637 1326
rect 650 1323 653 1346
rect 626 1313 637 1316
rect 626 1273 629 1313
rect 650 1296 653 1306
rect 642 1293 653 1296
rect 610 1263 629 1266
rect 590 1213 597 1216
rect 602 1213 605 1236
rect 610 1223 621 1226
rect 626 1223 629 1263
rect 642 1236 645 1293
rect 634 1233 645 1236
rect 594 1196 597 1213
rect 610 1203 613 1216
rect 586 1193 613 1196
rect 570 1133 577 1136
rect 586 1133 589 1193
rect 594 1133 597 1146
rect 562 1083 565 1126
rect 574 1056 577 1133
rect 570 1053 577 1056
rect 570 1033 573 1053
rect 546 1023 565 1026
rect 506 953 517 956
rect 490 933 493 946
rect 506 926 509 953
rect 474 923 493 926
rect 506 923 517 926
rect 474 913 477 923
rect 490 896 493 923
rect 482 893 493 896
rect 370 813 381 816
rect 378 736 381 813
rect 386 743 389 806
rect 378 733 389 736
rect 338 536 341 556
rect 338 533 345 536
rect 342 486 345 533
rect 354 523 357 586
rect 378 526 381 546
rect 370 523 381 526
rect 338 483 345 486
rect 322 393 325 406
rect 338 403 341 483
rect 370 446 373 523
rect 370 443 381 446
rect 370 413 373 426
rect 378 423 381 443
rect 90 373 117 376
rect 90 333 93 373
rect 218 333 221 376
rect 258 356 261 376
rect 258 353 265 356
rect 138 256 141 326
rect 202 313 205 326
rect 138 253 181 256
rect 178 226 181 253
rect 170 223 181 226
rect 138 176 141 206
rect 98 173 141 176
rect 170 176 173 223
rect 186 176 189 216
rect 218 213 221 306
rect 250 303 253 326
rect 262 296 265 353
rect 346 333 349 346
rect 346 313 349 326
rect 258 293 265 296
rect 258 203 261 293
rect 354 256 357 336
rect 378 313 381 326
rect 346 253 357 256
rect 306 213 309 226
rect 346 213 349 253
rect 170 173 181 176
rect 186 173 213 176
rect 98 133 101 173
rect 146 86 149 126
rect 178 123 181 173
rect 186 86 189 126
rect 202 113 205 136
rect 210 126 213 173
rect 218 133 221 146
rect 266 133 269 176
rect 346 166 349 206
rect 314 163 349 166
rect 210 123 221 126
rect 314 123 317 163
rect 354 123 357 226
rect 370 203 373 236
rect 386 226 389 733
rect 394 723 397 846
rect 402 733 405 786
rect 410 586 413 856
rect 434 793 437 816
rect 450 756 453 863
rect 482 796 485 893
rect 498 803 501 916
rect 514 866 517 923
rect 530 916 533 926
rect 538 923 541 1016
rect 546 1013 549 1023
rect 546 963 549 1006
rect 554 933 557 956
rect 546 923 557 926
rect 570 923 573 1016
rect 578 993 581 1016
rect 586 956 589 1126
rect 602 1123 605 1186
rect 610 1123 613 1193
rect 618 1156 621 1223
rect 634 1163 637 1233
rect 642 1203 645 1216
rect 618 1153 637 1156
rect 650 1153 653 1216
rect 658 1173 661 1386
rect 618 1133 621 1146
rect 594 993 597 1006
rect 586 953 597 956
rect 586 933 589 946
rect 594 923 597 953
rect 546 916 549 923
rect 530 913 549 916
rect 554 913 589 916
rect 506 863 517 866
rect 482 793 493 796
rect 450 753 461 756
rect 434 613 437 726
rect 450 703 453 736
rect 458 723 461 753
rect 466 733 469 746
rect 482 723 485 736
rect 490 723 493 793
rect 506 743 509 863
rect 514 726 517 826
rect 522 813 525 846
rect 506 723 517 726
rect 450 593 453 616
rect 474 593 477 606
rect 394 583 413 586
rect 394 543 397 583
rect 402 563 445 566
rect 394 523 397 536
rect 402 533 405 563
rect 418 533 421 546
rect 442 523 445 563
rect 490 503 493 696
rect 506 666 509 723
rect 506 663 517 666
rect 514 613 517 663
rect 522 596 525 806
rect 530 753 533 866
rect 554 846 557 913
rect 546 843 557 846
rect 538 803 541 816
rect 546 736 549 843
rect 562 816 565 826
rect 554 813 565 816
rect 570 813 573 826
rect 578 813 581 836
rect 586 826 589 913
rect 586 823 597 826
rect 554 796 557 813
rect 570 803 581 806
rect 554 793 569 796
rect 506 593 525 596
rect 506 486 509 593
rect 522 523 525 576
rect 530 553 533 736
rect 538 733 549 736
rect 566 736 569 793
rect 578 743 581 803
rect 566 733 573 736
rect 538 713 541 733
rect 546 723 557 726
rect 546 656 549 723
rect 538 653 549 656
rect 538 576 541 653
rect 554 616 557 716
rect 570 713 573 733
rect 578 723 581 736
rect 586 723 589 823
rect 602 813 605 1016
rect 610 1003 613 1076
rect 618 1033 621 1126
rect 618 966 621 1016
rect 626 983 629 1126
rect 634 1086 637 1153
rect 642 1123 645 1146
rect 666 1136 669 1456
rect 674 1403 677 1546
rect 706 1536 709 1776
rect 722 1756 725 1903
rect 730 1793 733 1806
rect 714 1753 725 1756
rect 714 1696 717 1753
rect 730 1733 733 1766
rect 754 1736 757 1926
rect 770 1923 773 1943
rect 778 1933 781 1966
rect 786 1923 789 1973
rect 770 1836 773 1896
rect 766 1833 773 1836
rect 766 1756 769 1833
rect 786 1766 789 1806
rect 810 1803 813 1816
rect 810 1766 813 1786
rect 778 1763 789 1766
rect 802 1763 813 1766
rect 766 1753 773 1756
rect 754 1733 765 1736
rect 754 1713 757 1726
rect 762 1696 765 1733
rect 714 1693 725 1696
rect 722 1636 725 1693
rect 758 1693 765 1696
rect 758 1636 761 1693
rect 722 1633 749 1636
rect 758 1633 765 1636
rect 690 1533 709 1536
rect 690 1483 693 1533
rect 698 1516 701 1526
rect 706 1516 709 1526
rect 698 1513 709 1516
rect 674 1333 677 1376
rect 674 1183 677 1316
rect 682 1143 685 1426
rect 690 1353 693 1396
rect 690 1333 693 1346
rect 650 1123 653 1136
rect 666 1133 681 1136
rect 658 1103 661 1126
rect 666 1113 669 1126
rect 634 1083 645 1086
rect 634 1013 637 1056
rect 642 1043 645 1083
rect 678 1076 681 1133
rect 690 1083 693 1326
rect 698 1313 701 1513
rect 706 1403 709 1506
rect 714 1503 717 1606
rect 722 1603 725 1616
rect 738 1613 741 1626
rect 746 1616 749 1633
rect 746 1613 753 1616
rect 738 1593 741 1606
rect 722 1513 725 1566
rect 722 1413 725 1486
rect 730 1423 733 1536
rect 738 1523 741 1556
rect 750 1546 753 1613
rect 762 1553 765 1633
rect 746 1543 753 1546
rect 746 1523 749 1543
rect 738 1413 741 1446
rect 706 1263 709 1346
rect 714 1226 717 1326
rect 722 1243 725 1406
rect 730 1333 733 1406
rect 754 1386 757 1526
rect 770 1443 773 1753
rect 778 1686 781 1763
rect 802 1706 805 1763
rect 818 1733 821 1926
rect 826 1916 829 1973
rect 834 1933 837 2006
rect 842 1923 845 1956
rect 854 1936 857 2123
rect 850 1933 857 1936
rect 866 1933 869 2176
rect 874 2173 893 2176
rect 898 2173 901 2356
rect 906 2283 909 2446
rect 922 2386 925 2493
rect 962 2443 965 2563
rect 978 2536 981 2846
rect 994 2776 997 2873
rect 1010 2873 1021 2876
rect 1010 2796 1013 2873
rect 1026 2813 1029 2926
rect 1042 2913 1045 2926
rect 1050 2823 1053 2966
rect 1058 2963 1077 2966
rect 1058 2926 1061 2963
rect 1082 2956 1085 3016
rect 1090 2973 1093 3093
rect 1114 3073 1117 3093
rect 1122 3083 1125 3116
rect 1130 3103 1133 3136
rect 1074 2953 1085 2956
rect 1066 2933 1069 2946
rect 1058 2923 1069 2926
rect 1066 2913 1069 2923
rect 1074 2896 1077 2953
rect 1106 2933 1109 3026
rect 1138 3023 1141 3126
rect 1146 3013 1149 3293
rect 1162 3236 1165 3336
rect 1242 3333 1245 3356
rect 1186 3303 1189 3316
rect 1242 3313 1245 3326
rect 1162 3233 1181 3236
rect 1066 2893 1077 2896
rect 1034 2813 1053 2816
rect 1066 2813 1069 2893
rect 1082 2836 1085 2926
rect 1098 2893 1101 2916
rect 1106 2886 1109 2926
rect 1098 2883 1109 2886
rect 1082 2833 1089 2836
rect 1026 2803 1061 2806
rect 1010 2793 1021 2796
rect 990 2773 997 2776
rect 990 2706 993 2773
rect 1002 2723 1005 2746
rect 1018 2736 1021 2793
rect 1018 2733 1029 2736
rect 1042 2733 1045 2756
rect 990 2703 997 2706
rect 994 2636 997 2703
rect 1026 2686 1029 2733
rect 1042 2693 1045 2726
rect 1050 2723 1053 2736
rect 1058 2696 1061 2803
rect 1066 2783 1069 2806
rect 1066 2716 1069 2756
rect 1074 2726 1077 2816
rect 1086 2776 1089 2833
rect 1082 2773 1089 2776
rect 1082 2753 1085 2773
rect 1090 2733 1093 2746
rect 1074 2723 1093 2726
rect 1066 2713 1085 2716
rect 1058 2693 1069 2696
rect 986 2633 997 2636
rect 1018 2683 1029 2686
rect 986 2586 989 2633
rect 994 2603 997 2616
rect 1002 2593 1005 2616
rect 986 2583 997 2586
rect 970 2533 981 2536
rect 970 2496 973 2533
rect 978 2513 981 2526
rect 986 2523 989 2576
rect 994 2566 997 2583
rect 994 2563 1001 2566
rect 998 2516 1001 2563
rect 1018 2516 1021 2683
rect 1034 2556 1037 2646
rect 1050 2623 1053 2676
rect 1066 2636 1069 2693
rect 1082 2646 1085 2713
rect 1090 2703 1093 2716
rect 1058 2633 1069 2636
rect 1078 2643 1085 2646
rect 1050 2603 1053 2616
rect 994 2513 1001 2516
rect 1010 2513 1021 2516
rect 1030 2553 1037 2556
rect 970 2493 977 2496
rect 946 2386 949 2406
rect 922 2383 949 2386
rect 922 2256 925 2383
rect 974 2376 977 2493
rect 994 2436 997 2513
rect 970 2373 977 2376
rect 986 2433 997 2436
rect 970 2356 973 2373
rect 962 2353 973 2356
rect 930 2266 933 2286
rect 930 2263 937 2266
rect 906 2253 925 2256
rect 874 2106 877 2173
rect 906 2166 909 2253
rect 914 2193 917 2216
rect 934 2176 937 2263
rect 946 2213 949 2236
rect 962 2226 965 2353
rect 970 2323 973 2346
rect 986 2276 989 2433
rect 994 2413 997 2426
rect 978 2273 989 2276
rect 962 2223 969 2226
rect 890 2163 909 2166
rect 930 2173 937 2176
rect 874 2103 881 2106
rect 878 2036 881 2103
rect 890 2036 893 2163
rect 930 2066 933 2173
rect 954 2163 957 2216
rect 966 2156 969 2223
rect 962 2153 969 2156
rect 938 2123 941 2146
rect 962 2136 965 2153
rect 958 2133 965 2136
rect 958 2086 961 2133
rect 970 2113 973 2126
rect 946 2083 961 2086
rect 930 2063 937 2066
rect 878 2033 885 2036
rect 890 2033 909 2036
rect 826 1913 833 1916
rect 830 1746 833 1913
rect 850 1856 853 1933
rect 858 1923 869 1926
rect 874 1906 877 1936
rect 870 1903 877 1906
rect 870 1856 873 1903
rect 882 1866 885 2033
rect 906 1976 909 2033
rect 906 1973 917 1976
rect 890 1876 893 1936
rect 898 1913 901 1926
rect 914 1883 917 1973
rect 934 1956 937 2063
rect 946 1966 949 2083
rect 978 2036 981 2273
rect 986 2173 989 2206
rect 994 2156 997 2356
rect 1002 2313 1005 2326
rect 1010 2296 1013 2513
rect 1030 2506 1033 2553
rect 1042 2533 1045 2546
rect 1050 2533 1053 2586
rect 1042 2513 1045 2526
rect 1030 2503 1037 2506
rect 1018 2306 1021 2446
rect 1026 2413 1029 2436
rect 1034 2353 1037 2503
rect 1050 2443 1053 2526
rect 1042 2333 1045 2406
rect 1050 2373 1053 2416
rect 1026 2313 1029 2326
rect 1018 2303 1029 2306
rect 1006 2293 1013 2296
rect 1006 2236 1009 2293
rect 1002 2233 1009 2236
rect 1002 2173 1005 2233
rect 1010 2213 1013 2226
rect 1010 2193 1013 2206
rect 1018 2203 1021 2296
rect 1026 2216 1029 2303
rect 1042 2223 1045 2256
rect 1026 2213 1045 2216
rect 1050 2183 1053 2326
rect 990 2153 997 2156
rect 990 2046 993 2153
rect 1002 2116 1005 2136
rect 1026 2133 1029 2146
rect 1050 2133 1053 2176
rect 1010 2123 1021 2126
rect 1002 2113 1013 2116
rect 990 2043 997 2046
rect 974 2033 981 2036
rect 954 2003 957 2016
rect 974 1976 977 2033
rect 986 2013 989 2026
rect 974 1973 981 1976
rect 946 1963 953 1966
rect 934 1953 941 1956
rect 938 1896 941 1953
rect 950 1916 953 1963
rect 962 1923 965 1946
rect 930 1893 941 1896
rect 946 1913 953 1916
rect 946 1893 949 1913
rect 890 1873 917 1876
rect 882 1863 893 1866
rect 850 1853 861 1856
rect 870 1853 877 1856
rect 858 1776 861 1853
rect 850 1773 861 1776
rect 850 1756 853 1773
rect 874 1756 877 1853
rect 890 1816 893 1863
rect 826 1743 833 1746
rect 846 1753 853 1756
rect 858 1753 877 1756
rect 886 1813 893 1816
rect 886 1756 889 1813
rect 886 1753 893 1756
rect 818 1713 821 1726
rect 802 1703 813 1706
rect 778 1683 789 1686
rect 786 1603 789 1683
rect 810 1636 813 1703
rect 810 1633 821 1636
rect 810 1613 813 1626
rect 778 1413 781 1426
rect 770 1393 773 1406
rect 754 1383 781 1386
rect 738 1323 741 1366
rect 746 1246 749 1336
rect 754 1323 757 1356
rect 762 1256 765 1336
rect 770 1303 773 1326
rect 778 1313 781 1383
rect 786 1256 789 1546
rect 794 1413 797 1426
rect 802 1403 805 1566
rect 810 1523 813 1586
rect 810 1336 813 1446
rect 794 1323 797 1336
rect 802 1333 813 1336
rect 802 1306 805 1333
rect 762 1253 789 1256
rect 798 1303 805 1306
rect 746 1243 765 1246
rect 698 1223 717 1226
rect 698 1123 701 1223
rect 706 1213 733 1216
rect 706 1176 709 1213
rect 722 1193 725 1206
rect 746 1203 749 1236
rect 754 1213 757 1226
rect 762 1203 765 1243
rect 706 1173 717 1176
rect 714 1126 717 1173
rect 746 1146 749 1166
rect 770 1146 773 1246
rect 778 1203 781 1253
rect 786 1196 789 1246
rect 798 1236 801 1303
rect 794 1233 801 1236
rect 794 1206 797 1233
rect 802 1213 805 1226
rect 794 1203 805 1206
rect 730 1143 749 1146
rect 714 1123 725 1126
rect 730 1106 733 1143
rect 722 1103 733 1106
rect 678 1073 685 1076
rect 650 1003 653 1066
rect 682 1056 685 1073
rect 682 1053 693 1056
rect 610 913 613 966
rect 618 963 625 966
rect 622 906 625 963
rect 634 923 645 926
rect 658 913 661 1006
rect 674 993 677 1006
rect 674 946 677 956
rect 666 943 677 946
rect 666 906 669 936
rect 618 903 625 906
rect 650 903 669 906
rect 610 803 613 826
rect 594 743 605 746
rect 594 706 597 736
rect 562 703 597 706
rect 602 636 605 743
rect 610 723 613 756
rect 618 713 621 903
rect 674 886 677 943
rect 682 933 685 1046
rect 690 956 693 1053
rect 722 1036 725 1103
rect 722 1033 733 1036
rect 698 963 701 1016
rect 706 983 709 1016
rect 690 953 701 956
rect 670 883 677 886
rect 670 826 673 883
rect 658 813 661 826
rect 670 823 677 826
rect 634 763 637 806
rect 666 733 669 806
rect 674 733 677 823
rect 642 723 677 726
rect 586 633 605 636
rect 554 613 573 616
rect 538 573 549 576
rect 466 483 509 486
rect 394 423 437 426
rect 394 403 397 423
rect 402 413 421 416
rect 434 413 437 423
rect 402 403 413 406
rect 402 243 405 386
rect 410 363 413 403
rect 418 353 421 413
rect 442 393 445 446
rect 410 313 413 336
rect 418 323 421 346
rect 434 326 437 346
rect 434 323 441 326
rect 378 223 389 226
rect 146 83 189 86
rect 378 23 381 223
rect 386 213 397 216
rect 402 213 405 236
rect 418 213 421 226
rect 394 196 397 206
rect 394 193 413 196
rect 394 133 397 176
rect 402 123 405 136
rect 410 133 413 193
rect 418 123 421 146
rect 426 133 429 306
rect 438 206 441 323
rect 434 203 441 206
rect 434 133 437 203
rect 450 136 453 336
rect 458 323 461 426
rect 466 406 469 483
rect 474 413 525 416
rect 466 403 493 406
rect 498 393 501 406
rect 506 346 509 406
rect 530 403 533 436
rect 538 416 541 526
rect 546 446 549 573
rect 554 523 557 613
rect 562 516 565 536
rect 570 523 573 536
rect 578 533 581 606
rect 586 576 589 633
rect 586 573 597 576
rect 578 516 581 526
rect 554 453 557 516
rect 562 513 581 516
rect 594 506 597 573
rect 586 503 597 506
rect 546 443 573 446
rect 554 423 565 426
rect 570 423 573 443
rect 562 416 565 423
rect 538 413 557 416
rect 562 413 581 416
rect 466 333 469 346
rect 482 343 509 346
rect 538 343 541 413
rect 466 143 469 246
rect 490 213 493 336
rect 522 273 525 326
rect 546 323 557 326
rect 546 296 549 316
rect 554 313 557 323
rect 562 313 565 406
rect 578 396 581 413
rect 586 403 589 503
rect 578 393 597 396
rect 602 393 605 416
rect 554 303 565 306
rect 570 296 573 326
rect 578 313 581 326
rect 586 303 589 336
rect 594 313 597 393
rect 610 296 613 606
rect 634 593 637 616
rect 642 546 645 723
rect 682 636 685 926
rect 690 903 693 936
rect 698 783 701 953
rect 714 926 717 996
rect 722 943 725 1006
rect 690 723 693 736
rect 698 723 701 776
rect 706 763 709 926
rect 714 923 721 926
rect 718 836 721 923
rect 714 833 721 836
rect 714 796 717 833
rect 722 803 725 816
rect 714 793 725 796
rect 706 656 709 756
rect 722 733 725 793
rect 730 726 733 1033
rect 738 853 741 1136
rect 746 1133 749 1143
rect 754 1143 773 1146
rect 778 1193 789 1196
rect 746 1073 749 1126
rect 754 1106 757 1143
rect 762 1123 765 1136
rect 754 1103 765 1106
rect 746 993 749 1056
rect 754 1013 757 1096
rect 762 1063 765 1103
rect 770 1096 773 1136
rect 778 1113 781 1193
rect 794 1136 797 1196
rect 802 1173 805 1203
rect 786 1133 797 1136
rect 802 1133 805 1166
rect 770 1093 781 1096
rect 746 933 749 956
rect 754 923 757 976
rect 762 873 765 1026
rect 770 1016 773 1086
rect 778 1023 781 1093
rect 786 1053 789 1133
rect 794 1043 797 1126
rect 802 1103 805 1126
rect 770 1013 789 1016
rect 794 1013 797 1026
rect 802 1013 805 1036
rect 770 933 773 1006
rect 778 946 781 1006
rect 786 1003 789 1013
rect 810 996 813 1326
rect 818 1243 821 1633
rect 826 1583 829 1743
rect 834 1593 837 1726
rect 846 1666 849 1753
rect 846 1663 853 1666
rect 826 1533 845 1536
rect 826 1496 829 1526
rect 834 1513 837 1526
rect 826 1493 833 1496
rect 830 1426 833 1493
rect 826 1423 833 1426
rect 826 1366 829 1423
rect 834 1383 837 1406
rect 842 1403 845 1533
rect 826 1363 833 1366
rect 830 1276 833 1363
rect 842 1333 845 1396
rect 850 1343 853 1663
rect 858 1573 861 1753
rect 874 1733 877 1746
rect 866 1713 869 1726
rect 866 1613 869 1646
rect 866 1536 869 1596
rect 858 1533 869 1536
rect 858 1513 861 1533
rect 874 1453 877 1726
rect 882 1693 885 1726
rect 890 1626 893 1753
rect 898 1736 901 1806
rect 906 1793 909 1816
rect 914 1746 917 1873
rect 930 1806 933 1893
rect 938 1813 941 1826
rect 930 1803 941 1806
rect 914 1743 925 1746
rect 898 1733 933 1736
rect 906 1713 909 1726
rect 890 1623 909 1626
rect 882 1603 893 1606
rect 890 1586 893 1603
rect 886 1583 893 1586
rect 886 1506 889 1583
rect 898 1563 901 1616
rect 906 1543 909 1623
rect 914 1566 917 1726
rect 922 1613 925 1646
rect 922 1586 925 1606
rect 930 1603 933 1733
rect 938 1723 941 1803
rect 954 1616 957 1886
rect 978 1696 981 1973
rect 970 1693 981 1696
rect 938 1596 941 1616
rect 946 1603 949 1616
rect 954 1613 965 1616
rect 954 1596 957 1606
rect 938 1593 957 1596
rect 962 1586 965 1613
rect 922 1583 965 1586
rect 970 1583 973 1693
rect 986 1663 989 1996
rect 978 1596 981 1616
rect 986 1613 989 1636
rect 994 1623 997 2043
rect 1002 1983 1005 2106
rect 1010 1953 1013 2113
rect 1026 2103 1029 2116
rect 1018 1993 1021 2036
rect 1002 1913 1005 1926
rect 1018 1923 1021 1976
rect 1026 1916 1029 2026
rect 1018 1913 1029 1916
rect 1018 1856 1021 1913
rect 1018 1853 1025 1856
rect 1002 1803 1005 1816
rect 1022 1796 1025 1853
rect 1018 1793 1025 1796
rect 1002 1703 1005 1726
rect 1002 1613 1005 1696
rect 1010 1606 1013 1686
rect 986 1603 997 1606
rect 978 1593 989 1596
rect 914 1563 933 1566
rect 886 1503 893 1506
rect 890 1446 893 1503
rect 890 1443 897 1446
rect 866 1383 869 1406
rect 882 1346 885 1396
rect 894 1366 897 1443
rect 906 1383 909 1536
rect 914 1393 917 1416
rect 930 1376 933 1563
rect 874 1343 885 1346
rect 890 1363 897 1366
rect 906 1373 933 1376
rect 842 1323 853 1326
rect 842 1283 845 1323
rect 830 1273 853 1276
rect 826 1193 829 1206
rect 806 993 813 996
rect 778 943 797 946
rect 794 933 797 943
rect 770 843 773 926
rect 786 903 789 926
rect 746 793 749 806
rect 778 753 781 876
rect 806 866 809 993
rect 806 863 813 866
rect 714 723 733 726
rect 706 653 717 656
rect 682 633 693 636
rect 706 613 709 626
rect 650 566 653 606
rect 714 603 717 653
rect 722 583 725 616
rect 730 596 733 606
rect 738 603 741 616
rect 746 603 749 736
rect 786 733 789 856
rect 794 813 797 826
rect 770 713 773 726
rect 754 613 757 646
rect 810 636 813 863
rect 818 746 821 1186
rect 850 1176 853 1273
rect 858 1246 861 1336
rect 866 1263 869 1326
rect 858 1243 865 1246
rect 874 1243 877 1343
rect 882 1283 885 1336
rect 826 1173 853 1176
rect 826 976 829 1173
rect 862 1166 865 1243
rect 874 1173 877 1216
rect 862 1163 877 1166
rect 834 986 837 1146
rect 850 1133 853 1146
rect 850 986 853 1006
rect 874 1003 877 1163
rect 882 996 885 1166
rect 890 1106 893 1363
rect 898 1163 901 1346
rect 906 1333 909 1373
rect 938 1353 941 1566
rect 946 1516 949 1576
rect 954 1523 957 1546
rect 986 1523 989 1593
rect 994 1523 997 1603
rect 1002 1603 1013 1606
rect 946 1513 957 1516
rect 946 1413 949 1426
rect 922 1333 925 1346
rect 906 1233 909 1326
rect 906 1213 909 1226
rect 898 1123 901 1146
rect 890 1103 897 1106
rect 894 1036 897 1103
rect 834 983 853 986
rect 866 993 885 996
rect 890 1033 897 1036
rect 890 993 893 1033
rect 898 1003 901 1016
rect 826 973 837 976
rect 826 813 829 926
rect 834 923 837 973
rect 834 813 837 906
rect 842 793 845 983
rect 866 933 869 993
rect 914 976 917 1286
rect 890 973 917 976
rect 890 933 893 973
rect 914 943 917 966
rect 898 933 917 936
rect 850 906 853 926
rect 858 923 869 926
rect 874 923 885 926
rect 850 903 857 906
rect 854 826 857 903
rect 850 823 857 826
rect 850 803 853 823
rect 866 806 869 923
rect 882 833 885 923
rect 898 853 901 926
rect 914 916 917 933
rect 910 913 917 916
rect 910 856 913 913
rect 922 873 925 1276
rect 930 1136 933 1246
rect 946 1193 949 1386
rect 954 1323 957 1513
rect 1002 1506 1005 1603
rect 1018 1596 1021 1793
rect 1026 1603 1029 1706
rect 1018 1593 1029 1596
rect 1018 1566 1021 1586
rect 994 1503 1005 1506
rect 1014 1563 1021 1566
rect 1014 1506 1017 1563
rect 1026 1513 1029 1593
rect 1014 1503 1021 1506
rect 962 1383 965 1436
rect 994 1426 997 1503
rect 994 1423 1005 1426
rect 1010 1423 1013 1456
rect 1002 1406 1005 1423
rect 962 1323 965 1346
rect 970 1196 973 1406
rect 986 1403 1005 1406
rect 1010 1393 1013 1406
rect 1018 1366 1021 1503
rect 986 1363 1021 1366
rect 986 1236 989 1363
rect 994 1273 997 1356
rect 1002 1303 1005 1326
rect 962 1193 973 1196
rect 978 1233 989 1236
rect 930 1133 941 1136
rect 930 1043 933 1126
rect 938 1093 941 1133
rect 930 1013 933 1026
rect 938 1013 941 1086
rect 946 1063 949 1186
rect 954 1046 957 1166
rect 962 1106 965 1193
rect 962 1103 969 1106
rect 950 1043 957 1046
rect 930 886 933 996
rect 950 956 953 1043
rect 966 1016 969 1103
rect 978 1016 981 1233
rect 986 1193 989 1216
rect 986 1133 989 1176
rect 1002 1136 1005 1176
rect 994 1133 1005 1136
rect 1010 1156 1013 1356
rect 1018 1163 1021 1336
rect 1026 1323 1029 1446
rect 1034 1396 1037 2126
rect 1042 2003 1053 2006
rect 1058 1966 1061 2633
rect 1066 2563 1069 2616
rect 1078 2576 1081 2643
rect 1090 2623 1093 2636
rect 1078 2573 1085 2576
rect 1066 2553 1077 2556
rect 1066 2496 1069 2546
rect 1074 2513 1077 2553
rect 1066 2493 1073 2496
rect 1070 2416 1073 2493
rect 1066 2413 1073 2416
rect 1066 2393 1069 2413
rect 1066 2333 1069 2346
rect 1074 2333 1077 2356
rect 1066 2313 1069 2326
rect 1074 2236 1077 2326
rect 1066 2233 1077 2236
rect 1066 2123 1069 2233
rect 1074 2203 1077 2226
rect 1074 2033 1077 2196
rect 1082 2176 1085 2573
rect 1090 2543 1093 2576
rect 1098 2526 1101 2883
rect 1106 2793 1109 2806
rect 1114 2726 1117 3006
rect 1138 2993 1141 3006
rect 1146 2956 1149 3006
rect 1138 2953 1149 2956
rect 1138 2936 1141 2953
rect 1130 2933 1141 2936
rect 1138 2906 1141 2926
rect 1146 2923 1149 2946
rect 1154 2916 1157 3166
rect 1162 3116 1165 3216
rect 1178 3213 1181 3233
rect 1194 3203 1197 3216
rect 1202 3193 1205 3206
rect 1218 3203 1221 3236
rect 1258 3226 1261 3316
rect 1274 3236 1277 3326
rect 1298 3313 1301 3416
rect 1306 3323 1309 3336
rect 1314 3333 1365 3336
rect 1370 3333 1373 3366
rect 1274 3233 1281 3236
rect 1170 3133 1173 3166
rect 1202 3123 1205 3156
rect 1162 3113 1173 3116
rect 1170 3056 1173 3113
rect 1166 3053 1173 3056
rect 1166 2956 1169 3053
rect 1202 3036 1205 3116
rect 1210 3103 1213 3146
rect 1226 3133 1229 3176
rect 1226 3106 1229 3126
rect 1222 3103 1229 3106
rect 1222 3036 1225 3103
rect 1186 3033 1205 3036
rect 1210 3033 1225 3036
rect 1178 2963 1181 3006
rect 1162 2953 1169 2956
rect 1186 2956 1189 3033
rect 1194 3003 1197 3016
rect 1186 2953 1197 2956
rect 1162 2923 1165 2953
rect 1170 2916 1173 2936
rect 1178 2923 1181 2936
rect 1186 2923 1189 2946
rect 1194 2916 1197 2953
rect 1154 2913 1165 2916
rect 1170 2913 1181 2916
rect 1130 2903 1141 2906
rect 1130 2846 1133 2903
rect 1146 2876 1149 2896
rect 1162 2893 1173 2896
rect 1146 2873 1153 2876
rect 1130 2843 1141 2846
rect 1122 2813 1125 2826
rect 1138 2796 1141 2843
rect 1106 2723 1117 2726
rect 1130 2793 1141 2796
rect 1106 2553 1109 2723
rect 1130 2716 1133 2793
rect 1150 2786 1153 2873
rect 1146 2783 1153 2786
rect 1146 2723 1149 2783
rect 1162 2746 1165 2893
rect 1178 2883 1181 2913
rect 1186 2913 1197 2916
rect 1202 2913 1205 2976
rect 1170 2813 1173 2876
rect 1186 2826 1189 2913
rect 1210 2833 1213 3033
rect 1218 2873 1221 3026
rect 1226 2856 1229 3016
rect 1234 2993 1237 3166
rect 1242 3033 1245 3226
rect 1258 3223 1269 3226
rect 1266 3186 1269 3206
rect 1262 3183 1269 3186
rect 1250 3013 1253 3136
rect 1262 3036 1265 3183
rect 1278 3176 1281 3233
rect 1274 3173 1281 3176
rect 1262 3033 1269 3036
rect 1266 3013 1269 3033
rect 1222 2853 1229 2856
rect 1234 2853 1237 2946
rect 1258 2943 1261 3006
rect 1182 2823 1189 2826
rect 1202 2823 1213 2826
rect 1182 2756 1185 2823
rect 1182 2753 1189 2756
rect 1162 2743 1169 2746
rect 1114 2546 1117 2716
rect 1130 2713 1141 2716
rect 1122 2603 1125 2616
rect 1130 2603 1133 2636
rect 1122 2593 1133 2596
rect 1138 2586 1141 2713
rect 1154 2706 1157 2736
rect 1150 2703 1157 2706
rect 1150 2606 1153 2703
rect 1166 2696 1169 2743
rect 1162 2693 1169 2696
rect 1150 2603 1157 2606
rect 1130 2583 1141 2586
rect 1154 2586 1157 2603
rect 1162 2596 1165 2693
rect 1170 2613 1173 2626
rect 1162 2593 1173 2596
rect 1154 2583 1165 2586
rect 1094 2523 1101 2526
rect 1106 2543 1117 2546
rect 1094 2456 1097 2523
rect 1094 2453 1101 2456
rect 1106 2453 1109 2543
rect 1114 2523 1117 2536
rect 1122 2516 1125 2566
rect 1114 2513 1125 2516
rect 1090 2423 1093 2436
rect 1090 2403 1093 2416
rect 1090 2193 1093 2396
rect 1098 2296 1101 2453
rect 1114 2446 1117 2513
rect 1106 2443 1117 2446
rect 1106 2413 1109 2443
rect 1106 2313 1109 2406
rect 1114 2393 1117 2436
rect 1122 2423 1125 2496
rect 1098 2293 1105 2296
rect 1102 2186 1105 2293
rect 1114 2223 1117 2306
rect 1122 2276 1125 2416
rect 1130 2286 1133 2583
rect 1138 2413 1141 2546
rect 1146 2463 1149 2536
rect 1154 2513 1157 2526
rect 1138 2333 1141 2346
rect 1146 2303 1149 2456
rect 1154 2403 1157 2426
rect 1162 2323 1165 2583
rect 1170 2573 1173 2593
rect 1178 2566 1181 2736
rect 1186 2723 1189 2753
rect 1194 2733 1197 2816
rect 1202 2796 1205 2823
rect 1202 2793 1213 2796
rect 1210 2736 1213 2793
rect 1222 2756 1225 2853
rect 1242 2843 1245 2936
rect 1250 2916 1253 2936
rect 1266 2926 1269 3006
rect 1274 2993 1277 3173
rect 1290 3156 1293 3226
rect 1306 3183 1309 3216
rect 1314 3203 1317 3333
rect 1362 3326 1365 3333
rect 1338 3236 1341 3256
rect 1334 3233 1341 3236
rect 1286 3153 1293 3156
rect 1286 3086 1289 3153
rect 1298 3133 1301 3146
rect 1322 3126 1325 3216
rect 1334 3156 1337 3233
rect 1334 3153 1341 3156
rect 1298 3093 1301 3126
rect 1306 3123 1325 3126
rect 1286 3083 1293 3086
rect 1290 3026 1293 3083
rect 1290 3023 1301 3026
rect 1274 2933 1277 2956
rect 1290 2936 1293 3016
rect 1298 2976 1301 3023
rect 1306 3013 1309 3123
rect 1322 3093 1325 3116
rect 1330 3076 1333 3136
rect 1322 3073 1333 3076
rect 1322 3006 1325 3073
rect 1322 3003 1333 3006
rect 1330 2983 1333 3003
rect 1298 2973 1317 2976
rect 1266 2923 1277 2926
rect 1250 2913 1257 2916
rect 1254 2846 1257 2913
rect 1274 2876 1277 2923
rect 1266 2873 1277 2876
rect 1282 2873 1285 2936
rect 1290 2933 1301 2936
rect 1250 2843 1257 2846
rect 1222 2753 1229 2756
rect 1202 2733 1213 2736
rect 1226 2733 1229 2753
rect 1202 2653 1205 2733
rect 1234 2666 1237 2806
rect 1226 2663 1237 2666
rect 1226 2646 1229 2663
rect 1222 2643 1229 2646
rect 1186 2603 1189 2616
rect 1170 2563 1181 2566
rect 1194 2596 1197 2616
rect 1202 2603 1205 2626
rect 1210 2596 1213 2616
rect 1194 2593 1213 2596
rect 1170 2413 1173 2563
rect 1178 2533 1189 2536
rect 1194 2526 1197 2593
rect 1222 2556 1225 2643
rect 1222 2553 1229 2556
rect 1186 2523 1197 2526
rect 1186 2413 1189 2516
rect 1194 2453 1197 2523
rect 1210 2513 1213 2536
rect 1218 2456 1221 2536
rect 1214 2453 1221 2456
rect 1226 2456 1229 2553
rect 1234 2503 1237 2656
rect 1242 2636 1245 2836
rect 1250 2643 1253 2843
rect 1258 2823 1277 2826
rect 1282 2823 1285 2836
rect 1258 2813 1261 2823
rect 1274 2816 1277 2823
rect 1258 2793 1261 2806
rect 1266 2803 1269 2816
rect 1274 2813 1285 2816
rect 1290 2803 1293 2926
rect 1298 2896 1301 2933
rect 1306 2913 1309 2946
rect 1298 2893 1305 2896
rect 1314 2893 1317 2973
rect 1322 2943 1325 2976
rect 1302 2816 1305 2893
rect 1314 2826 1317 2876
rect 1314 2823 1325 2826
rect 1302 2813 1309 2816
rect 1258 2743 1269 2746
rect 1290 2733 1293 2766
rect 1298 2726 1301 2806
rect 1242 2633 1253 2636
rect 1242 2593 1245 2606
rect 1242 2486 1245 2566
rect 1250 2543 1253 2633
rect 1242 2483 1253 2486
rect 1226 2453 1245 2456
rect 1202 2406 1205 2426
rect 1170 2403 1181 2406
rect 1186 2403 1205 2406
rect 1130 2283 1157 2286
rect 1122 2273 1141 2276
rect 1114 2203 1117 2216
rect 1098 2183 1105 2186
rect 1082 2173 1089 2176
rect 1086 2046 1089 2173
rect 1082 2043 1089 2046
rect 1066 1993 1069 2026
rect 1082 2023 1085 2043
rect 1074 1993 1077 2006
rect 1050 1963 1069 1966
rect 1082 1963 1085 2006
rect 1098 2003 1101 2183
rect 1122 2146 1125 2236
rect 1130 2213 1133 2246
rect 1138 2213 1141 2273
rect 1122 2143 1141 2146
rect 1106 2096 1109 2116
rect 1122 2113 1125 2136
rect 1106 2093 1125 2096
rect 1106 1996 1109 2086
rect 1122 2076 1125 2093
rect 1098 1993 1109 1996
rect 1118 2073 1125 2076
rect 1118 1996 1121 2073
rect 1118 1993 1125 1996
rect 1042 1923 1045 1936
rect 1050 1893 1053 1963
rect 1066 1956 1069 1963
rect 1042 1813 1045 1826
rect 1050 1793 1053 1816
rect 1042 1713 1045 1726
rect 1050 1693 1053 1736
rect 1058 1683 1061 1956
rect 1066 1953 1093 1956
rect 1082 1933 1085 1946
rect 1090 1933 1093 1953
rect 1098 1943 1101 1993
rect 1066 1923 1077 1926
rect 1082 1913 1093 1916
rect 1098 1906 1101 1926
rect 1114 1913 1117 1976
rect 1122 1923 1125 1993
rect 1130 1906 1133 2136
rect 1090 1903 1101 1906
rect 1090 1853 1093 1903
rect 1066 1796 1069 1826
rect 1090 1823 1093 1836
rect 1074 1813 1093 1816
rect 1082 1803 1093 1806
rect 1066 1793 1085 1796
rect 1082 1736 1085 1793
rect 1082 1733 1093 1736
rect 1066 1653 1069 1726
rect 1082 1706 1085 1726
rect 1074 1703 1085 1706
rect 1090 1703 1093 1733
rect 1074 1646 1077 1703
rect 1098 1696 1101 1896
rect 1106 1886 1109 1906
rect 1126 1903 1133 1906
rect 1106 1883 1117 1886
rect 1114 1836 1117 1883
rect 1106 1833 1117 1836
rect 1126 1836 1129 1903
rect 1126 1833 1133 1836
rect 1106 1813 1109 1833
rect 1130 1813 1133 1833
rect 1114 1793 1117 1806
rect 1122 1773 1125 1806
rect 1106 1723 1109 1766
rect 1066 1643 1077 1646
rect 1082 1693 1101 1696
rect 1042 1563 1045 1626
rect 1058 1583 1061 1626
rect 1042 1516 1045 1546
rect 1050 1523 1053 1536
rect 1042 1513 1053 1516
rect 1042 1413 1045 1426
rect 1034 1393 1041 1396
rect 1038 1316 1041 1393
rect 1034 1313 1041 1316
rect 1050 1316 1053 1486
rect 1058 1323 1061 1536
rect 1066 1443 1069 1643
rect 1082 1586 1085 1693
rect 1106 1653 1109 1716
rect 1090 1623 1093 1636
rect 1098 1603 1101 1616
rect 1106 1596 1109 1606
rect 1098 1593 1109 1596
rect 1074 1576 1077 1586
rect 1082 1583 1101 1586
rect 1074 1573 1093 1576
rect 1074 1533 1085 1536
rect 1090 1513 1093 1573
rect 1074 1373 1077 1436
rect 1082 1403 1085 1426
rect 1090 1393 1093 1416
rect 1066 1333 1069 1366
rect 1098 1353 1101 1583
rect 1106 1513 1109 1556
rect 1114 1433 1117 1756
rect 1130 1753 1133 1806
rect 1138 1746 1141 2143
rect 1146 2123 1149 2276
rect 1154 2106 1157 2283
rect 1162 2216 1165 2306
rect 1170 2233 1173 2336
rect 1186 2326 1189 2403
rect 1214 2346 1217 2453
rect 1202 2326 1205 2346
rect 1214 2343 1221 2346
rect 1186 2323 1197 2326
rect 1202 2323 1209 2326
rect 1186 2303 1189 2316
rect 1194 2313 1197 2323
rect 1162 2213 1169 2216
rect 1166 2146 1169 2213
rect 1178 2203 1181 2246
rect 1150 2103 1157 2106
rect 1162 2143 1169 2146
rect 1150 2016 1153 2103
rect 1150 2013 1157 2016
rect 1146 1823 1149 1996
rect 1146 1756 1149 1816
rect 1154 1803 1157 2013
rect 1162 1966 1165 2143
rect 1170 2013 1173 2126
rect 1178 2113 1181 2126
rect 1178 2003 1181 2026
rect 1186 2016 1189 2236
rect 1194 2116 1197 2286
rect 1206 2246 1209 2323
rect 1218 2273 1221 2343
rect 1202 2243 1209 2246
rect 1202 2173 1205 2243
rect 1226 2226 1229 2416
rect 1234 2303 1237 2446
rect 1242 2283 1245 2453
rect 1210 2126 1213 2226
rect 1222 2223 1229 2226
rect 1222 2156 1225 2223
rect 1250 2216 1253 2483
rect 1258 2286 1261 2726
rect 1274 2713 1277 2726
rect 1282 2723 1301 2726
rect 1306 2723 1309 2813
rect 1322 2746 1325 2823
rect 1338 2803 1341 3153
rect 1346 3113 1349 3226
rect 1354 3123 1357 3326
rect 1362 3323 1373 3326
rect 1370 3283 1373 3316
rect 1386 3306 1389 3356
rect 1442 3333 1445 3386
rect 1450 3333 1453 3356
rect 1474 3333 1477 3346
rect 1546 3343 1557 3346
rect 1382 3303 1389 3306
rect 1362 3203 1365 3236
rect 1382 3216 1385 3303
rect 1402 3296 1405 3316
rect 1402 3293 1413 3296
rect 1370 3213 1385 3216
rect 1362 3096 1365 3146
rect 1354 3093 1365 3096
rect 1346 2933 1349 2996
rect 1354 2973 1357 3093
rect 1362 3003 1365 3016
rect 1370 2996 1373 3213
rect 1378 3166 1381 3206
rect 1378 3163 1385 3166
rect 1382 3096 1385 3163
rect 1394 3113 1397 3286
rect 1410 3236 1413 3293
rect 1402 3233 1413 3236
rect 1402 3213 1405 3233
rect 1458 3226 1461 3326
rect 1474 3293 1477 3316
rect 1482 3283 1485 3336
rect 1506 3326 1509 3336
rect 1490 3266 1493 3326
rect 1486 3263 1493 3266
rect 1498 3323 1509 3326
rect 1458 3223 1477 3226
rect 1426 3183 1429 3216
rect 1402 3133 1405 3166
rect 1426 3136 1429 3156
rect 1442 3153 1445 3216
rect 1450 3193 1453 3206
rect 1410 3133 1429 3136
rect 1458 3136 1461 3216
rect 1458 3133 1465 3136
rect 1382 3093 1389 3096
rect 1386 3026 1389 3093
rect 1378 3023 1389 3026
rect 1378 3006 1381 3023
rect 1434 3013 1437 3036
rect 1442 3013 1445 3126
rect 1450 3083 1453 3126
rect 1462 3076 1465 3133
rect 1458 3073 1465 3076
rect 1378 3003 1389 3006
rect 1362 2993 1373 2996
rect 1386 2996 1389 3003
rect 1458 2996 1461 3073
rect 1474 3026 1477 3223
rect 1486 3156 1489 3263
rect 1486 3153 1493 3156
rect 1490 3133 1493 3153
rect 1498 3143 1501 3323
rect 1506 3256 1509 3316
rect 1554 3293 1557 3336
rect 1610 3333 1613 3396
rect 1570 3283 1573 3326
rect 1506 3253 1525 3256
rect 1506 3213 1509 3226
rect 1506 3193 1509 3206
rect 1514 3193 1517 3246
rect 1522 3186 1525 3253
rect 1602 3246 1605 3266
rect 1594 3243 1605 3246
rect 1514 3183 1525 3186
rect 1466 3023 1477 3026
rect 1466 3003 1469 3023
rect 1386 2993 1397 2996
rect 1426 2993 1461 2996
rect 1354 2823 1357 2936
rect 1362 2816 1365 2993
rect 1318 2743 1325 2746
rect 1266 2333 1269 2626
rect 1274 2563 1277 2616
rect 1282 2603 1285 2723
rect 1298 2606 1301 2696
rect 1290 2603 1301 2606
rect 1274 2533 1277 2546
rect 1282 2533 1285 2576
rect 1290 2516 1293 2603
rect 1306 2596 1309 2716
rect 1318 2636 1321 2743
rect 1338 2726 1341 2796
rect 1346 2733 1349 2816
rect 1354 2813 1365 2816
rect 1370 2813 1373 2926
rect 1378 2813 1381 2936
rect 1386 2906 1389 2976
rect 1394 2943 1397 2993
rect 1394 2916 1397 2926
rect 1402 2923 1405 2956
rect 1410 2933 1413 2966
rect 1410 2916 1413 2926
rect 1394 2913 1413 2916
rect 1466 2913 1469 2956
rect 1386 2903 1397 2906
rect 1394 2886 1397 2903
rect 1474 2896 1477 2916
rect 1482 2903 1485 2936
rect 1490 2916 1493 3116
rect 1498 3103 1501 3136
rect 1498 3013 1501 3026
rect 1506 3003 1509 3046
rect 1514 3036 1517 3183
rect 1538 3146 1541 3216
rect 1594 3176 1597 3243
rect 1618 3213 1621 3376
rect 1634 3346 1637 3366
rect 1634 3343 1653 3346
rect 1722 3343 1725 3366
rect 1626 3293 1629 3336
rect 1634 3323 1637 3343
rect 1634 3216 1637 3236
rect 1642 3226 1645 3336
rect 1650 3333 1653 3343
rect 1722 3293 1725 3326
rect 1642 3223 1661 3226
rect 1634 3213 1653 3216
rect 1610 3186 1613 3206
rect 1626 3193 1629 3206
rect 1658 3203 1661 3223
rect 1610 3183 1653 3186
rect 1594 3173 1605 3176
rect 1530 3143 1541 3146
rect 1522 3053 1525 3126
rect 1530 3043 1533 3143
rect 1546 3113 1549 3156
rect 1554 3103 1557 3136
rect 1514 3033 1533 3036
rect 1530 3023 1533 3033
rect 1514 3003 1517 3016
rect 1506 2923 1509 2976
rect 1514 2933 1517 2966
rect 1514 2923 1525 2926
rect 1514 2916 1517 2923
rect 1490 2913 1517 2916
rect 1474 2893 1485 2896
rect 1394 2883 1405 2886
rect 1402 2836 1405 2883
rect 1482 2836 1485 2893
rect 1394 2833 1405 2836
rect 1474 2833 1485 2836
rect 1302 2593 1309 2596
rect 1314 2633 1321 2636
rect 1302 2536 1305 2593
rect 1286 2513 1293 2516
rect 1298 2533 1305 2536
rect 1266 2303 1269 2326
rect 1258 2283 1265 2286
rect 1234 2213 1253 2216
rect 1262 2216 1265 2283
rect 1274 2266 1277 2506
rect 1286 2436 1289 2513
rect 1298 2473 1301 2533
rect 1314 2526 1317 2633
rect 1322 2593 1325 2616
rect 1330 2593 1333 2726
rect 1338 2723 1349 2726
rect 1338 2666 1341 2716
rect 1346 2686 1349 2723
rect 1354 2693 1357 2813
rect 1394 2806 1397 2833
rect 1402 2813 1445 2816
rect 1370 2803 1397 2806
rect 1362 2733 1365 2746
rect 1370 2723 1373 2803
rect 1378 2706 1381 2736
rect 1386 2713 1389 2796
rect 1394 2723 1397 2803
rect 1374 2703 1381 2706
rect 1346 2683 1357 2686
rect 1338 2663 1345 2666
rect 1342 2606 1345 2663
rect 1338 2603 1345 2606
rect 1338 2586 1341 2603
rect 1330 2583 1341 2586
rect 1314 2523 1321 2526
rect 1282 2433 1289 2436
rect 1282 2396 1285 2433
rect 1306 2426 1309 2516
rect 1318 2436 1321 2523
rect 1290 2423 1309 2426
rect 1314 2433 1321 2436
rect 1314 2413 1317 2433
rect 1306 2403 1317 2406
rect 1282 2393 1301 2396
rect 1282 2273 1285 2336
rect 1290 2323 1293 2346
rect 1274 2263 1285 2266
rect 1282 2246 1285 2263
rect 1282 2243 1289 2246
rect 1262 2213 1277 2216
rect 1222 2153 1229 2156
rect 1202 2123 1213 2126
rect 1194 2113 1205 2116
rect 1194 2016 1197 2026
rect 1186 2013 1197 2016
rect 1162 1963 1173 1966
rect 1162 1933 1165 1956
rect 1146 1753 1157 1756
rect 1122 1733 1125 1746
rect 1130 1733 1133 1746
rect 1138 1743 1149 1746
rect 1122 1613 1125 1676
rect 1130 1656 1133 1726
rect 1138 1663 1141 1736
rect 1146 1733 1149 1743
rect 1130 1653 1141 1656
rect 1122 1593 1125 1606
rect 1138 1583 1141 1653
rect 1146 1603 1149 1726
rect 1154 1703 1157 1753
rect 1162 1713 1165 1856
rect 1170 1843 1173 1963
rect 1178 1836 1181 1946
rect 1186 1933 1189 2006
rect 1194 1936 1197 2013
rect 1202 1973 1205 2113
rect 1210 2003 1213 2036
rect 1194 1933 1205 1936
rect 1174 1833 1181 1836
rect 1174 1756 1177 1833
rect 1170 1753 1177 1756
rect 1170 1646 1173 1753
rect 1162 1643 1173 1646
rect 1122 1416 1125 1536
rect 1130 1506 1133 1526
rect 1130 1503 1137 1506
rect 1134 1426 1137 1503
rect 1146 1436 1149 1566
rect 1154 1483 1157 1606
rect 1146 1433 1157 1436
rect 1162 1433 1165 1643
rect 1170 1613 1173 1636
rect 1134 1423 1149 1426
rect 1106 1406 1109 1416
rect 1122 1413 1141 1416
rect 1106 1403 1117 1406
rect 1122 1386 1125 1396
rect 1130 1393 1133 1406
rect 1138 1403 1141 1413
rect 1146 1386 1149 1423
rect 1154 1416 1157 1433
rect 1154 1413 1165 1416
rect 1122 1383 1149 1386
rect 1050 1313 1061 1316
rect 1026 1213 1029 1236
rect 1010 1153 1029 1156
rect 986 1113 989 1126
rect 994 1113 997 1126
rect 994 1076 997 1096
rect 994 1073 1001 1076
rect 986 1023 989 1066
rect 966 1013 973 1016
rect 978 1013 989 1016
rect 950 953 957 956
rect 938 903 941 926
rect 946 923 949 936
rect 954 933 957 953
rect 962 923 965 1006
rect 930 883 937 886
rect 906 853 913 856
rect 906 833 909 853
rect 862 803 869 806
rect 818 743 829 746
rect 818 723 821 736
rect 762 613 765 626
rect 786 613 789 636
rect 806 633 813 636
rect 754 596 757 606
rect 794 603 797 616
rect 730 593 757 596
rect 806 586 809 633
rect 826 626 829 743
rect 834 686 837 786
rect 862 746 865 803
rect 862 743 869 746
rect 850 706 853 726
rect 866 723 869 743
rect 874 723 877 826
rect 882 803 885 826
rect 906 766 909 806
rect 934 796 937 883
rect 930 793 937 796
rect 930 766 933 793
rect 898 763 909 766
rect 926 763 933 766
rect 850 703 861 706
rect 834 683 845 686
rect 818 623 829 626
rect 806 583 813 586
rect 650 563 661 566
rect 626 543 645 546
rect 626 533 629 543
rect 634 523 637 536
rect 642 523 645 543
rect 658 516 661 563
rect 690 533 693 546
rect 642 513 661 516
rect 642 406 645 513
rect 674 486 677 526
rect 714 486 717 526
rect 674 483 717 486
rect 666 423 669 436
rect 650 413 669 416
rect 634 313 637 406
rect 642 403 669 406
rect 642 343 669 346
rect 674 343 677 406
rect 658 303 661 326
rect 546 293 573 296
rect 586 293 613 296
rect 538 213 549 216
rect 570 196 573 226
rect 562 193 573 196
rect 450 133 469 136
rect 434 86 437 126
rect 442 93 445 126
rect 450 86 453 133
rect 458 113 461 126
rect 474 123 477 156
rect 562 146 565 193
rect 586 153 589 293
rect 610 166 613 216
rect 658 196 661 216
rect 666 213 669 343
rect 674 333 685 336
rect 682 273 685 326
rect 690 293 693 426
rect 698 423 701 436
rect 714 356 717 436
rect 754 423 757 566
rect 810 563 813 583
rect 802 533 805 546
rect 818 543 821 623
rect 826 583 829 616
rect 834 573 837 616
rect 842 603 845 683
rect 858 646 861 703
rect 898 666 901 763
rect 926 716 929 763
rect 938 723 941 756
rect 926 713 933 716
rect 898 663 909 666
rect 850 643 861 646
rect 850 613 853 643
rect 858 603 861 616
rect 770 426 773 526
rect 850 523 853 566
rect 874 536 877 616
rect 906 576 909 663
rect 930 603 933 713
rect 906 573 917 576
rect 946 573 949 876
rect 954 803 957 816
rect 970 793 973 1013
rect 978 1003 989 1006
rect 998 996 1001 1073
rect 1010 1053 1013 1153
rect 1018 1133 1021 1146
rect 1026 1133 1029 1153
rect 1018 1023 1021 1116
rect 1026 1016 1029 1126
rect 994 993 1001 996
rect 1010 1013 1029 1016
rect 994 936 997 993
rect 982 933 997 936
rect 982 876 985 933
rect 1010 926 1013 1013
rect 1018 933 1021 946
rect 1026 933 1029 956
rect 1034 926 1037 1313
rect 1042 1213 1045 1256
rect 1042 1173 1045 1206
rect 1042 1113 1045 1166
rect 1050 1093 1053 1156
rect 1042 973 1045 1026
rect 1050 963 1053 1006
rect 1058 1003 1061 1306
rect 1066 1293 1069 1326
rect 1074 1323 1077 1336
rect 1090 1333 1093 1346
rect 1098 1316 1101 1336
rect 1090 1313 1101 1316
rect 1082 1213 1085 1226
rect 1082 1193 1085 1206
rect 1090 1153 1093 1313
rect 1106 1296 1109 1376
rect 1154 1366 1157 1406
rect 1102 1293 1109 1296
rect 1102 1156 1105 1293
rect 1102 1153 1109 1156
rect 1082 1133 1085 1146
rect 1106 1136 1109 1153
rect 1090 1133 1109 1136
rect 1066 1123 1085 1126
rect 1114 1123 1117 1366
rect 1122 1363 1157 1366
rect 1082 1103 1085 1116
rect 1066 1033 1085 1036
rect 1066 983 1069 1033
rect 1074 1016 1077 1026
rect 1082 1023 1085 1033
rect 1074 1013 1085 1016
rect 1082 1003 1085 1013
rect 1042 933 1053 936
rect 978 873 985 876
rect 978 786 981 873
rect 986 813 989 856
rect 970 783 981 786
rect 970 706 973 783
rect 978 713 981 726
rect 986 723 989 746
rect 994 726 997 926
rect 1002 923 1021 926
rect 1034 923 1045 926
rect 1010 893 1013 923
rect 1018 903 1021 916
rect 1002 813 1005 836
rect 1034 813 1037 826
rect 1010 733 1013 806
rect 1026 803 1037 806
rect 1042 766 1045 923
rect 1050 913 1053 933
rect 1066 883 1069 936
rect 1082 933 1085 946
rect 1090 936 1093 1096
rect 1114 1073 1117 1116
rect 1098 946 1101 1016
rect 1106 1013 1109 1056
rect 1122 993 1125 1363
rect 1130 1303 1133 1316
rect 1130 1096 1133 1276
rect 1138 1113 1141 1286
rect 1146 1213 1149 1356
rect 1154 1203 1157 1346
rect 1162 1276 1165 1413
rect 1170 1353 1173 1606
rect 1178 1553 1181 1736
rect 1186 1716 1189 1916
rect 1194 1883 1197 1926
rect 1202 1916 1205 1933
rect 1210 1923 1213 1946
rect 1202 1913 1213 1916
rect 1194 1803 1197 1826
rect 1202 1823 1205 1906
rect 1202 1736 1205 1806
rect 1210 1763 1213 1913
rect 1194 1733 1213 1736
rect 1194 1723 1197 1733
rect 1202 1716 1205 1726
rect 1186 1713 1205 1716
rect 1210 1713 1213 1733
rect 1186 1613 1189 1646
rect 1178 1533 1181 1546
rect 1186 1523 1189 1596
rect 1178 1413 1181 1486
rect 1170 1313 1173 1336
rect 1178 1323 1181 1346
rect 1186 1323 1189 1466
rect 1194 1306 1197 1706
rect 1202 1603 1205 1713
rect 1210 1603 1213 1626
rect 1202 1363 1205 1586
rect 1210 1346 1213 1546
rect 1218 1493 1221 2126
rect 1226 1813 1229 2153
rect 1234 2033 1237 2213
rect 1242 2176 1245 2206
rect 1242 2173 1249 2176
rect 1246 2046 1249 2173
rect 1242 2043 1249 2046
rect 1242 2026 1245 2043
rect 1258 2026 1261 2196
rect 1266 2036 1269 2206
rect 1274 2053 1277 2213
rect 1286 2146 1289 2243
rect 1282 2143 1289 2146
rect 1298 2146 1301 2393
rect 1322 2343 1325 2416
rect 1306 2306 1309 2326
rect 1306 2303 1317 2306
rect 1314 2256 1317 2303
rect 1306 2253 1317 2256
rect 1306 2233 1309 2253
rect 1330 2243 1333 2583
rect 1338 2533 1341 2566
rect 1338 2433 1341 2446
rect 1306 2223 1333 2226
rect 1306 2213 1309 2223
rect 1298 2143 1309 2146
rect 1282 2123 1285 2143
rect 1282 2083 1285 2116
rect 1282 2036 1285 2046
rect 1266 2033 1285 2036
rect 1234 2023 1245 2026
rect 1250 2023 1261 2026
rect 1234 1813 1237 2023
rect 1242 2003 1245 2016
rect 1242 1853 1245 1926
rect 1250 1916 1253 2023
rect 1258 2013 1269 2016
rect 1274 2013 1277 2026
rect 1282 2013 1285 2033
rect 1258 1933 1261 1946
rect 1250 1913 1257 1916
rect 1254 1836 1257 1913
rect 1250 1833 1257 1836
rect 1250 1816 1253 1833
rect 1242 1813 1253 1816
rect 1242 1806 1245 1813
rect 1234 1803 1245 1806
rect 1226 1713 1229 1736
rect 1226 1463 1229 1666
rect 1234 1543 1237 1803
rect 1242 1706 1245 1726
rect 1250 1713 1253 1806
rect 1266 1776 1269 1936
rect 1258 1773 1269 1776
rect 1274 1916 1277 1926
rect 1282 1923 1285 2006
rect 1290 2003 1293 2126
rect 1306 2123 1309 2143
rect 1314 2136 1317 2216
rect 1338 2203 1341 2386
rect 1346 2243 1349 2536
rect 1354 2506 1357 2683
rect 1374 2646 1377 2703
rect 1374 2643 1381 2646
rect 1378 2626 1381 2643
rect 1362 2623 1381 2626
rect 1362 2523 1365 2623
rect 1386 2603 1389 2686
rect 1426 2636 1429 2726
rect 1434 2723 1437 2736
rect 1442 2723 1445 2813
rect 1450 2746 1453 2826
rect 1458 2813 1461 2826
rect 1474 2766 1477 2833
rect 1474 2763 1485 2766
rect 1450 2743 1461 2746
rect 1482 2743 1485 2763
rect 1490 2746 1493 2826
rect 1506 2823 1517 2826
rect 1522 2816 1525 2896
rect 1530 2863 1533 3006
rect 1538 3003 1541 3086
rect 1562 3063 1565 3166
rect 1546 2986 1549 3026
rect 1546 2983 1557 2986
rect 1538 2913 1541 2926
rect 1546 2923 1549 2976
rect 1554 2906 1557 2983
rect 1570 2963 1573 3126
rect 1602 3123 1605 3173
rect 1626 3086 1629 3126
rect 1610 3083 1629 3086
rect 1578 2946 1581 3046
rect 1610 3026 1613 3083
rect 1610 3023 1621 3026
rect 1618 3006 1621 3023
rect 1586 3003 1597 3006
rect 1610 3003 1621 3006
rect 1586 2956 1589 2976
rect 1610 2956 1613 3003
rect 1586 2953 1597 2956
rect 1610 2953 1621 2956
rect 1574 2943 1581 2946
rect 1550 2903 1557 2906
rect 1538 2823 1541 2876
rect 1514 2813 1525 2816
rect 1498 2793 1501 2806
rect 1490 2743 1505 2746
rect 1354 2503 1361 2506
rect 1358 2386 1361 2503
rect 1354 2383 1361 2386
rect 1354 2363 1357 2383
rect 1354 2333 1357 2346
rect 1362 2316 1365 2356
rect 1370 2326 1373 2556
rect 1378 2523 1381 2576
rect 1394 2546 1397 2626
rect 1402 2603 1405 2636
rect 1426 2633 1437 2636
rect 1390 2543 1397 2546
rect 1390 2456 1393 2543
rect 1390 2453 1397 2456
rect 1386 2416 1389 2436
rect 1394 2423 1397 2453
rect 1402 2433 1405 2536
rect 1418 2533 1421 2576
rect 1426 2563 1429 2626
rect 1434 2556 1437 2633
rect 1426 2553 1437 2556
rect 1386 2413 1397 2416
rect 1394 2363 1405 2366
rect 1378 2336 1381 2346
rect 1378 2333 1389 2336
rect 1370 2323 1381 2326
rect 1354 2313 1373 2316
rect 1346 2193 1349 2226
rect 1314 2133 1325 2136
rect 1314 2113 1317 2126
rect 1322 2106 1325 2133
rect 1306 2103 1325 2106
rect 1306 2086 1309 2103
rect 1302 2083 1309 2086
rect 1302 2026 1305 2083
rect 1302 2023 1309 2026
rect 1290 1943 1293 1986
rect 1298 1916 1301 2006
rect 1274 1913 1301 1916
rect 1242 1703 1253 1706
rect 1242 1623 1245 1636
rect 1242 1593 1245 1606
rect 1250 1543 1253 1703
rect 1258 1606 1261 1773
rect 1266 1663 1269 1766
rect 1266 1633 1269 1646
rect 1274 1623 1277 1913
rect 1282 1813 1285 1826
rect 1290 1816 1293 1846
rect 1298 1823 1301 1856
rect 1306 1833 1309 2023
rect 1314 2013 1317 2056
rect 1346 2053 1349 2136
rect 1322 2013 1333 2016
rect 1322 1996 1325 2006
rect 1330 2003 1341 2006
rect 1346 1996 1349 2006
rect 1322 1993 1349 1996
rect 1314 1966 1317 1986
rect 1314 1963 1325 1966
rect 1322 1856 1325 1963
rect 1338 1933 1341 1946
rect 1314 1853 1325 1856
rect 1290 1813 1301 1816
rect 1282 1606 1285 1716
rect 1290 1633 1293 1796
rect 1298 1683 1301 1813
rect 1314 1763 1317 1853
rect 1338 1836 1341 1896
rect 1346 1853 1349 1926
rect 1330 1833 1341 1836
rect 1330 1756 1333 1833
rect 1330 1753 1341 1756
rect 1306 1673 1309 1736
rect 1314 1733 1325 1736
rect 1314 1713 1317 1726
rect 1330 1693 1333 1736
rect 1258 1603 1269 1606
rect 1266 1546 1269 1603
rect 1258 1543 1269 1546
rect 1278 1603 1285 1606
rect 1234 1456 1237 1536
rect 1250 1503 1253 1526
rect 1226 1453 1237 1456
rect 1226 1426 1229 1453
rect 1218 1423 1229 1426
rect 1218 1413 1221 1423
rect 1258 1416 1261 1543
rect 1278 1536 1281 1603
rect 1290 1586 1293 1616
rect 1306 1593 1309 1626
rect 1322 1613 1325 1626
rect 1338 1613 1341 1753
rect 1314 1586 1317 1606
rect 1290 1583 1317 1586
rect 1278 1533 1285 1536
rect 1274 1503 1277 1516
rect 1226 1413 1237 1416
rect 1218 1403 1229 1406
rect 1162 1273 1173 1276
rect 1162 1226 1165 1266
rect 1170 1233 1173 1273
rect 1178 1243 1181 1306
rect 1186 1303 1197 1306
rect 1202 1343 1213 1346
rect 1226 1343 1229 1403
rect 1234 1356 1237 1413
rect 1242 1393 1245 1416
rect 1250 1413 1261 1416
rect 1234 1353 1245 1356
rect 1162 1223 1173 1226
rect 1170 1213 1173 1223
rect 1146 1193 1157 1196
rect 1130 1093 1137 1096
rect 1134 1016 1137 1093
rect 1130 1013 1137 1016
rect 1098 943 1109 946
rect 1090 933 1101 936
rect 1026 763 1045 766
rect 994 723 1005 726
rect 970 703 981 706
rect 978 656 981 703
rect 974 653 981 656
rect 1002 656 1005 723
rect 1026 716 1029 763
rect 1042 733 1045 756
rect 1050 743 1053 836
rect 1058 793 1061 806
rect 1018 713 1029 716
rect 1042 713 1053 716
rect 1002 653 1013 656
rect 954 593 957 616
rect 974 606 977 653
rect 986 613 989 646
rect 994 633 1005 636
rect 974 603 981 606
rect 994 603 997 616
rect 870 533 877 536
rect 870 476 873 533
rect 882 506 885 526
rect 882 503 893 506
rect 870 473 877 476
rect 874 453 877 473
rect 890 456 893 503
rect 914 466 917 573
rect 962 523 965 536
rect 978 476 981 603
rect 974 473 981 476
rect 914 463 949 466
rect 882 453 893 456
rect 882 436 885 453
rect 826 433 885 436
rect 762 423 773 426
rect 710 353 717 356
rect 698 313 701 336
rect 710 266 713 353
rect 722 323 725 346
rect 730 323 733 396
rect 738 333 741 416
rect 762 393 765 423
rect 818 403 821 416
rect 834 406 837 426
rect 834 403 845 406
rect 762 343 781 346
rect 762 333 765 343
rect 746 306 749 326
rect 762 316 765 326
rect 722 303 749 306
rect 754 313 765 316
rect 710 263 717 266
rect 698 213 701 226
rect 714 213 717 263
rect 722 233 725 303
rect 722 223 733 226
rect 738 206 741 286
rect 754 226 757 313
rect 770 306 773 336
rect 746 223 757 226
rect 762 303 773 306
rect 762 223 765 303
rect 778 283 781 343
rect 802 333 805 346
rect 810 323 813 376
rect 850 366 853 416
rect 818 363 853 366
rect 818 276 821 363
rect 810 273 821 276
rect 746 213 749 223
rect 722 203 741 206
rect 762 203 765 216
rect 810 203 813 273
rect 826 223 829 336
rect 858 323 861 376
rect 866 333 869 406
rect 874 343 893 346
rect 874 303 877 343
rect 882 333 893 336
rect 882 313 885 326
rect 658 193 669 196
rect 602 163 613 166
rect 522 133 525 146
rect 562 143 573 146
rect 570 123 573 143
rect 602 123 605 163
rect 634 133 637 156
rect 666 146 669 193
rect 658 143 669 146
rect 658 123 661 143
rect 722 123 725 203
rect 746 133 749 156
rect 770 93 773 126
rect 834 123 837 276
rect 850 213 869 216
rect 842 166 845 206
rect 874 203 877 246
rect 890 223 893 296
rect 898 283 901 426
rect 930 393 933 416
rect 946 403 949 463
rect 974 396 977 473
rect 986 413 989 526
rect 994 523 997 586
rect 1002 523 1005 633
rect 1010 533 1013 653
rect 1018 483 1021 713
rect 1034 616 1037 626
rect 1026 613 1037 616
rect 1026 576 1029 613
rect 1034 593 1037 606
rect 1042 603 1045 706
rect 1058 673 1061 736
rect 1066 703 1069 846
rect 1074 696 1077 896
rect 1082 703 1085 806
rect 1090 753 1093 866
rect 1090 706 1093 726
rect 1098 713 1101 933
rect 1106 923 1109 943
rect 1106 896 1109 916
rect 1114 903 1117 916
rect 1106 893 1117 896
rect 1106 813 1109 856
rect 1114 813 1117 893
rect 1114 773 1117 806
rect 1090 703 1101 706
rect 1074 693 1085 696
rect 1066 683 1077 686
rect 1026 573 1033 576
rect 1030 496 1033 573
rect 1050 563 1053 616
rect 1058 566 1061 626
rect 1066 583 1069 683
rect 1082 613 1085 693
rect 1090 603 1093 703
rect 1098 593 1101 616
rect 1058 563 1069 566
rect 1066 556 1069 563
rect 1042 533 1053 536
rect 1026 493 1033 496
rect 1050 493 1053 516
rect 1026 473 1029 493
rect 1026 413 1029 456
rect 1058 416 1061 556
rect 1066 553 1085 556
rect 1066 523 1069 553
rect 1082 523 1085 536
rect 1090 513 1093 536
rect 974 393 981 396
rect 978 376 981 393
rect 930 333 933 376
rect 978 373 1013 376
rect 962 333 989 336
rect 906 273 909 326
rect 922 293 925 326
rect 970 253 973 326
rect 978 293 981 316
rect 986 313 989 333
rect 994 313 997 326
rect 986 273 989 306
rect 1010 296 1013 373
rect 1002 293 1013 296
rect 1002 273 1005 293
rect 882 196 885 216
rect 898 213 901 226
rect 1002 213 1005 226
rect 850 193 885 196
rect 842 163 877 166
rect 850 133 853 146
rect 874 123 877 163
rect 434 83 453 86
rect 890 73 893 206
rect 954 176 957 206
rect 954 173 965 176
rect 962 133 965 173
rect 1034 166 1037 416
rect 1050 413 1061 416
rect 1050 383 1053 413
rect 1074 406 1077 506
rect 1082 503 1093 506
rect 1082 423 1085 503
rect 1098 496 1101 516
rect 1090 493 1101 496
rect 1090 413 1093 493
rect 1058 403 1077 406
rect 1098 406 1101 436
rect 1106 423 1109 706
rect 1114 686 1117 756
rect 1122 693 1125 986
rect 1130 923 1133 1013
rect 1130 833 1133 906
rect 1138 826 1141 946
rect 1146 923 1149 1193
rect 1162 1156 1165 1206
rect 1178 1193 1181 1206
rect 1154 1133 1157 1156
rect 1162 1153 1181 1156
rect 1178 1143 1181 1153
rect 1162 1133 1181 1136
rect 1154 1116 1157 1126
rect 1154 1113 1173 1116
rect 1154 983 1157 1086
rect 1146 833 1149 866
rect 1130 773 1133 826
rect 1138 823 1149 826
rect 1154 823 1157 936
rect 1130 713 1133 756
rect 1130 686 1133 706
rect 1114 683 1133 686
rect 1114 623 1117 683
rect 1122 613 1125 626
rect 1122 506 1125 526
rect 1130 513 1133 666
rect 1138 596 1141 816
rect 1146 663 1149 823
rect 1154 723 1157 736
rect 1162 716 1165 1106
rect 1170 983 1173 1113
rect 1178 1103 1181 1133
rect 1170 863 1173 926
rect 1178 846 1181 1096
rect 1186 913 1189 1303
rect 1194 1193 1197 1236
rect 1194 1103 1197 1126
rect 1194 1013 1197 1036
rect 1194 933 1197 946
rect 1202 926 1205 1343
rect 1210 1323 1213 1336
rect 1218 1266 1221 1326
rect 1226 1273 1229 1336
rect 1234 1333 1237 1353
rect 1210 1263 1221 1266
rect 1210 1213 1213 1246
rect 1210 1123 1213 1146
rect 1218 1103 1221 1126
rect 1226 1096 1229 1206
rect 1234 1133 1237 1326
rect 1210 1093 1229 1096
rect 1210 1003 1213 1093
rect 1234 1086 1237 1106
rect 1218 1083 1237 1086
rect 1218 1006 1221 1083
rect 1226 1013 1237 1016
rect 1218 1003 1229 1006
rect 1210 936 1213 996
rect 1218 946 1221 996
rect 1226 953 1229 1003
rect 1218 943 1229 946
rect 1210 933 1221 936
rect 1194 893 1197 926
rect 1202 923 1213 926
rect 1202 876 1205 916
rect 1186 853 1189 876
rect 1198 873 1205 876
rect 1178 843 1189 846
rect 1178 813 1181 836
rect 1186 813 1189 843
rect 1170 726 1173 806
rect 1198 796 1201 873
rect 1210 863 1213 923
rect 1218 836 1221 933
rect 1210 833 1221 836
rect 1186 733 1189 796
rect 1198 793 1205 796
rect 1170 723 1177 726
rect 1154 713 1165 716
rect 1154 683 1157 713
rect 1146 623 1149 636
rect 1138 593 1149 596
rect 1138 513 1141 586
rect 1118 503 1125 506
rect 1118 436 1121 503
rect 1118 433 1125 436
rect 1122 413 1125 433
rect 1098 403 1117 406
rect 1058 333 1061 403
rect 1114 366 1117 403
rect 1114 363 1125 366
rect 1042 263 1045 316
rect 1106 313 1109 326
rect 1122 316 1125 363
rect 1130 336 1133 506
rect 1146 403 1149 593
rect 1154 563 1157 616
rect 1162 613 1165 696
rect 1174 656 1177 723
rect 1174 653 1181 656
rect 1170 603 1173 636
rect 1178 536 1181 653
rect 1186 576 1189 686
rect 1194 676 1197 776
rect 1202 733 1205 793
rect 1202 693 1205 726
rect 1194 673 1201 676
rect 1198 586 1201 673
rect 1210 616 1213 833
rect 1218 813 1221 826
rect 1226 766 1229 943
rect 1234 816 1237 946
rect 1242 903 1245 1346
rect 1250 1046 1253 1413
rect 1258 1323 1261 1406
rect 1266 1403 1269 1416
rect 1274 1413 1277 1496
rect 1282 1396 1285 1533
rect 1290 1503 1293 1536
rect 1298 1523 1301 1583
rect 1314 1563 1317 1583
rect 1330 1543 1333 1606
rect 1306 1533 1325 1536
rect 1322 1526 1325 1533
rect 1322 1523 1333 1526
rect 1346 1523 1349 1846
rect 1354 1723 1357 2313
rect 1362 2196 1365 2276
rect 1370 2213 1373 2286
rect 1378 2256 1381 2323
rect 1386 2266 1389 2333
rect 1394 2283 1397 2326
rect 1402 2273 1405 2363
rect 1386 2263 1405 2266
rect 1378 2253 1389 2256
rect 1362 2193 1369 2196
rect 1366 2106 1369 2193
rect 1378 2143 1381 2236
rect 1378 2113 1381 2126
rect 1386 2123 1389 2253
rect 1394 2123 1397 2226
rect 1366 2103 1381 2106
rect 1322 1496 1325 1516
rect 1290 1493 1325 1496
rect 1290 1476 1293 1493
rect 1290 1473 1297 1476
rect 1270 1393 1285 1396
rect 1270 1316 1273 1393
rect 1282 1323 1285 1366
rect 1294 1346 1297 1473
rect 1290 1343 1297 1346
rect 1306 1426 1309 1436
rect 1306 1423 1325 1426
rect 1266 1313 1273 1316
rect 1258 1133 1261 1266
rect 1266 1133 1269 1313
rect 1290 1273 1293 1343
rect 1298 1313 1301 1326
rect 1306 1283 1309 1423
rect 1330 1416 1333 1523
rect 1354 1516 1357 1656
rect 1350 1513 1357 1516
rect 1314 1333 1317 1416
rect 1322 1413 1333 1416
rect 1338 1413 1341 1486
rect 1350 1426 1353 1513
rect 1346 1423 1353 1426
rect 1322 1333 1325 1413
rect 1330 1323 1333 1376
rect 1338 1316 1341 1396
rect 1330 1313 1341 1316
rect 1330 1276 1333 1313
rect 1346 1296 1349 1423
rect 1354 1306 1357 1406
rect 1362 1323 1365 2026
rect 1370 1933 1373 2076
rect 1370 1893 1373 1926
rect 1370 1793 1373 1876
rect 1370 1733 1373 1766
rect 1378 1733 1381 2103
rect 1394 2066 1397 2116
rect 1402 2073 1405 2263
rect 1394 2063 1405 2066
rect 1386 1826 1389 2056
rect 1394 1863 1397 2056
rect 1402 1986 1405 2063
rect 1410 2053 1413 2496
rect 1426 2483 1429 2553
rect 1434 2513 1437 2536
rect 1442 2533 1445 2556
rect 1450 2466 1453 2736
rect 1458 2733 1461 2743
rect 1490 2716 1493 2736
rect 1482 2713 1493 2716
rect 1482 2646 1485 2713
rect 1482 2643 1493 2646
rect 1466 2613 1469 2626
rect 1490 2623 1493 2643
rect 1458 2586 1461 2606
rect 1458 2583 1465 2586
rect 1462 2516 1465 2583
rect 1458 2513 1465 2516
rect 1458 2493 1461 2513
rect 1450 2463 1469 2466
rect 1418 2056 1421 2416
rect 1426 2226 1429 2456
rect 1434 2343 1437 2406
rect 1434 2253 1437 2326
rect 1426 2223 1437 2226
rect 1426 2133 1429 2216
rect 1434 2173 1437 2223
rect 1442 2156 1445 2416
rect 1458 2413 1461 2456
rect 1450 2403 1461 2406
rect 1450 2323 1453 2346
rect 1466 2246 1469 2463
rect 1474 2413 1477 2616
rect 1502 2606 1505 2743
rect 1498 2603 1505 2606
rect 1514 2603 1517 2813
rect 1550 2796 1553 2903
rect 1562 2813 1565 2936
rect 1574 2836 1577 2943
rect 1594 2906 1597 2953
rect 1618 2933 1621 2953
rect 1586 2903 1597 2906
rect 1610 2906 1613 2926
rect 1626 2923 1629 3006
rect 1634 2983 1637 3136
rect 1650 3083 1653 3183
rect 1682 3143 1685 3156
rect 1682 3123 1701 3126
rect 1642 3003 1645 3056
rect 1690 3013 1693 3066
rect 1666 2966 1669 3006
rect 1682 3003 1693 3006
rect 1666 2963 1677 2966
rect 1642 2913 1645 2926
rect 1650 2906 1653 2926
rect 1610 2903 1653 2906
rect 1586 2853 1589 2903
rect 1574 2833 1581 2836
rect 1570 2803 1573 2816
rect 1578 2803 1581 2833
rect 1594 2823 1597 2886
rect 1626 2816 1629 2836
rect 1618 2813 1629 2816
rect 1530 2733 1533 2796
rect 1550 2793 1557 2796
rect 1546 2733 1549 2766
rect 1522 2603 1525 2636
rect 1490 2523 1493 2596
rect 1498 2473 1501 2603
rect 1530 2556 1533 2726
rect 1546 2713 1549 2726
rect 1554 2713 1557 2793
rect 1578 2723 1581 2776
rect 1618 2756 1621 2813
rect 1618 2753 1629 2756
rect 1586 2733 1605 2736
rect 1626 2723 1629 2753
rect 1602 2683 1605 2716
rect 1634 2666 1637 2903
rect 1642 2713 1645 2746
rect 1650 2723 1653 2816
rect 1658 2803 1661 2896
rect 1666 2803 1669 2936
rect 1674 2803 1677 2963
rect 1682 2923 1685 2936
rect 1706 2893 1709 3276
rect 1730 3166 1733 3396
rect 1738 3263 1741 3326
rect 1730 3163 1741 3166
rect 1738 3123 1741 3163
rect 1714 3033 1717 3046
rect 1722 2933 1725 3066
rect 1730 2923 1733 3016
rect 1746 2956 1749 3406
rect 1850 3346 1853 3366
rect 1802 3343 1837 3346
rect 1802 3333 1805 3343
rect 1834 3333 1837 3343
rect 1754 3116 1757 3306
rect 1762 3203 1765 3216
rect 1770 3213 1773 3326
rect 1842 3323 1845 3346
rect 1850 3343 1861 3346
rect 1826 3273 1829 3316
rect 1874 3296 1877 3416
rect 1930 3343 1933 3366
rect 1938 3333 1941 3396
rect 1866 3293 1877 3296
rect 1898 3293 1901 3326
rect 1786 3216 1789 3246
rect 1786 3213 1797 3216
rect 1770 3193 1773 3206
rect 1794 3203 1797 3213
rect 1802 3193 1805 3206
rect 1810 3193 1821 3196
rect 1762 3133 1765 3166
rect 1810 3153 1813 3193
rect 1786 3143 1813 3146
rect 1786 3136 1789 3143
rect 1778 3133 1789 3136
rect 1754 3113 1765 3116
rect 1742 2953 1749 2956
rect 1742 2906 1745 2953
rect 1762 2946 1765 3113
rect 1786 3083 1789 3126
rect 1802 3116 1805 3136
rect 1798 3113 1805 3116
rect 1786 3013 1789 3026
rect 1798 2956 1801 3113
rect 1810 3003 1813 3143
rect 1818 2996 1821 3146
rect 1826 3023 1829 3236
rect 1866 3216 1869 3293
rect 1858 3213 1869 3216
rect 1810 2993 1821 2996
rect 1798 2953 1805 2956
rect 1738 2903 1745 2906
rect 1754 2943 1765 2946
rect 1690 2836 1693 2856
rect 1738 2846 1741 2903
rect 1754 2856 1757 2943
rect 1762 2896 1765 2926
rect 1762 2893 1773 2896
rect 1754 2853 1761 2856
rect 1738 2843 1749 2846
rect 1690 2833 1697 2836
rect 1682 2783 1685 2826
rect 1694 2756 1697 2833
rect 1746 2826 1749 2843
rect 1626 2663 1637 2666
rect 1538 2613 1541 2646
rect 1538 2593 1541 2606
rect 1546 2573 1549 2626
rect 1626 2616 1629 2663
rect 1650 2623 1653 2656
rect 1554 2603 1557 2616
rect 1626 2613 1637 2616
rect 1634 2573 1637 2613
rect 1658 2593 1661 2666
rect 1490 2403 1493 2446
rect 1506 2426 1509 2536
rect 1514 2526 1517 2556
rect 1530 2553 1541 2556
rect 1522 2533 1525 2546
rect 1514 2523 1525 2526
rect 1514 2496 1517 2523
rect 1522 2513 1525 2523
rect 1514 2493 1525 2496
rect 1522 2436 1525 2493
rect 1498 2423 1509 2426
rect 1514 2433 1525 2436
rect 1490 2336 1493 2346
rect 1474 2333 1493 2336
rect 1438 2153 1445 2156
rect 1450 2243 1469 2246
rect 1426 2113 1429 2126
rect 1438 2076 1441 2153
rect 1438 2073 1445 2076
rect 1418 2053 1437 2056
rect 1410 2003 1421 2006
rect 1402 1983 1409 1986
rect 1406 1866 1409 1983
rect 1402 1863 1409 1866
rect 1402 1843 1405 1863
rect 1418 1853 1421 1966
rect 1426 1943 1429 2046
rect 1386 1823 1421 1826
rect 1386 1803 1389 1823
rect 1402 1803 1405 1816
rect 1410 1793 1413 1816
rect 1386 1733 1397 1736
rect 1402 1733 1405 1756
rect 1370 1393 1373 1706
rect 1378 1463 1381 1726
rect 1394 1723 1405 1726
rect 1410 1723 1413 1746
rect 1386 1363 1389 1686
rect 1394 1493 1397 1696
rect 1402 1683 1405 1723
rect 1410 1613 1413 1666
rect 1418 1653 1421 1823
rect 1426 1643 1429 1756
rect 1426 1613 1429 1626
rect 1402 1603 1413 1606
rect 1402 1523 1405 1536
rect 1410 1513 1413 1596
rect 1418 1583 1421 1606
rect 1434 1596 1437 2053
rect 1442 1983 1445 2073
rect 1450 1963 1453 2243
rect 1458 2223 1461 2236
rect 1474 2216 1477 2276
rect 1458 2213 1477 2216
rect 1458 2203 1461 2213
rect 1482 2203 1485 2316
rect 1490 2276 1493 2333
rect 1498 2326 1501 2423
rect 1506 2386 1509 2416
rect 1514 2403 1517 2433
rect 1538 2416 1541 2553
rect 1562 2543 1581 2546
rect 1538 2413 1549 2416
rect 1562 2413 1565 2543
rect 1570 2516 1573 2526
rect 1578 2523 1581 2543
rect 1586 2523 1597 2526
rect 1586 2516 1589 2523
rect 1570 2513 1589 2516
rect 1522 2403 1533 2406
rect 1530 2393 1533 2403
rect 1506 2383 1517 2386
rect 1506 2333 1509 2346
rect 1498 2323 1509 2326
rect 1506 2293 1509 2323
rect 1514 2276 1517 2383
rect 1538 2373 1541 2396
rect 1546 2353 1549 2413
rect 1546 2323 1549 2346
rect 1570 2326 1573 2436
rect 1578 2413 1581 2446
rect 1554 2323 1573 2326
rect 1522 2286 1525 2306
rect 1522 2283 1533 2286
rect 1490 2273 1501 2276
rect 1498 2216 1501 2273
rect 1490 2213 1501 2216
rect 1510 2273 1517 2276
rect 1458 2193 1469 2196
rect 1458 2183 1461 2193
rect 1482 2156 1485 2176
rect 1474 2153 1485 2156
rect 1458 2103 1461 2136
rect 1474 2036 1477 2153
rect 1490 2146 1493 2213
rect 1510 2166 1513 2273
rect 1530 2236 1533 2283
rect 1522 2233 1533 2236
rect 1510 2163 1517 2166
rect 1490 2143 1509 2146
rect 1498 2123 1501 2136
rect 1490 2046 1493 2116
rect 1506 2103 1509 2143
rect 1490 2043 1501 2046
rect 1474 2033 1485 2036
rect 1458 1943 1461 2006
rect 1474 1983 1477 2006
rect 1442 1933 1461 1936
rect 1442 1903 1445 1926
rect 1450 1893 1453 1926
rect 1442 1783 1445 1796
rect 1450 1776 1453 1796
rect 1442 1773 1453 1776
rect 1442 1693 1445 1773
rect 1450 1703 1453 1736
rect 1430 1593 1437 1596
rect 1442 1593 1445 1656
rect 1394 1406 1397 1466
rect 1410 1413 1413 1436
rect 1418 1413 1421 1526
rect 1430 1496 1433 1593
rect 1442 1543 1445 1576
rect 1450 1556 1453 1686
rect 1458 1653 1461 1933
rect 1466 1903 1469 1926
rect 1474 1903 1477 1976
rect 1482 1923 1485 2033
rect 1490 1943 1493 2006
rect 1498 2003 1501 2043
rect 1514 2016 1517 2163
rect 1506 2013 1517 2016
rect 1506 1976 1509 2013
rect 1502 1973 1509 1976
rect 1522 1973 1525 2233
rect 1530 2036 1533 2216
rect 1538 2103 1541 2136
rect 1546 2123 1549 2206
rect 1554 2176 1557 2323
rect 1562 2223 1565 2246
rect 1570 2226 1573 2316
rect 1570 2223 1589 2226
rect 1594 2216 1597 2516
rect 1610 2403 1613 2416
rect 1618 2413 1621 2546
rect 1626 2503 1629 2536
rect 1634 2523 1645 2526
rect 1618 2366 1621 2406
rect 1634 2403 1637 2456
rect 1642 2376 1645 2486
rect 1658 2463 1661 2526
rect 1650 2403 1653 2446
rect 1642 2373 1653 2376
rect 1658 2373 1661 2416
rect 1618 2363 1645 2366
rect 1602 2313 1605 2326
rect 1610 2323 1613 2356
rect 1626 2336 1629 2356
rect 1642 2346 1645 2363
rect 1650 2356 1653 2373
rect 1674 2366 1677 2756
rect 1690 2753 1697 2756
rect 1706 2823 1749 2826
rect 1690 2733 1693 2753
rect 1706 2736 1709 2823
rect 1702 2733 1709 2736
rect 1690 2513 1693 2696
rect 1702 2626 1705 2733
rect 1702 2623 1709 2626
rect 1706 2603 1709 2623
rect 1714 2613 1717 2726
rect 1722 2613 1725 2736
rect 1730 2733 1733 2806
rect 1730 2556 1733 2726
rect 1738 2663 1741 2816
rect 1746 2723 1749 2806
rect 1758 2756 1761 2853
rect 1754 2753 1761 2756
rect 1754 2623 1757 2753
rect 1770 2736 1773 2893
rect 1794 2846 1797 2936
rect 1786 2843 1797 2846
rect 1786 2796 1789 2843
rect 1802 2803 1805 2953
rect 1810 2803 1813 2993
rect 1818 2913 1821 2936
rect 1826 2883 1829 2926
rect 1834 2876 1837 3166
rect 1858 3116 1861 3213
rect 1882 3123 1885 3206
rect 1890 3193 1893 3286
rect 1922 3226 1925 3326
rect 1954 3323 1957 3356
rect 1922 3223 1933 3226
rect 1906 3203 1909 3216
rect 1914 3143 1917 3166
rect 1890 3133 1917 3136
rect 1898 3123 1909 3126
rect 1858 3113 1877 3116
rect 1842 2913 1845 3096
rect 1874 3026 1877 3113
rect 1906 3076 1909 3123
rect 1914 3083 1917 3133
rect 1930 3076 1933 3223
rect 1970 3213 1973 3326
rect 1986 3286 1989 3336
rect 2002 3326 2005 3376
rect 2010 3333 2013 3366
rect 2002 3323 2013 3326
rect 2026 3296 2029 3376
rect 2090 3336 2093 3396
rect 2106 3346 2109 3386
rect 2138 3356 2141 3416
rect 2354 3393 2365 3396
rect 2138 3353 2149 3356
rect 2106 3343 2125 3346
rect 1986 3283 1997 3286
rect 1978 3213 1981 3226
rect 1994 3206 1997 3283
rect 1954 3133 1957 3206
rect 1986 3203 1997 3206
rect 2018 3203 2021 3296
rect 2026 3293 2037 3296
rect 2034 3226 2037 3293
rect 2082 3263 2085 3336
rect 2090 3333 2101 3336
rect 2090 3266 2093 3326
rect 2106 3323 2109 3343
rect 2114 3276 2117 3336
rect 2122 3333 2125 3343
rect 2114 3273 2125 3276
rect 2090 3263 2117 3266
rect 2098 3236 2101 3256
rect 2098 3233 2105 3236
rect 2026 3223 2037 3226
rect 1978 3116 1981 3136
rect 1986 3123 1989 3203
rect 1994 3133 2005 3136
rect 1906 3073 1933 3076
rect 1970 3113 1981 3116
rect 1850 3013 1853 3026
rect 1874 3023 1885 3026
rect 1850 2903 1853 2936
rect 1858 2923 1861 2936
rect 1866 2896 1869 3016
rect 1882 2936 1885 3023
rect 1882 2933 1901 2936
rect 1890 2896 1893 2916
rect 1830 2873 1837 2876
rect 1842 2893 1869 2896
rect 1882 2893 1893 2896
rect 1818 2813 1821 2866
rect 1830 2806 1833 2873
rect 1826 2803 1833 2806
rect 1786 2793 1797 2796
rect 1766 2733 1773 2736
rect 1730 2553 1737 2556
rect 1698 2543 1725 2546
rect 1698 2533 1701 2543
rect 1722 2533 1725 2543
rect 1722 2503 1725 2516
rect 1734 2496 1737 2553
rect 1754 2543 1757 2606
rect 1766 2536 1769 2733
rect 1762 2533 1769 2536
rect 1746 2513 1749 2526
rect 1730 2493 1737 2496
rect 1698 2396 1701 2416
rect 1694 2393 1701 2396
rect 1674 2363 1685 2366
rect 1650 2353 1669 2356
rect 1642 2343 1661 2346
rect 1618 2333 1629 2336
rect 1626 2286 1629 2326
rect 1562 2193 1565 2216
rect 1578 2213 1597 2216
rect 1618 2283 1629 2286
rect 1554 2173 1561 2176
rect 1558 2106 1561 2173
rect 1578 2156 1581 2213
rect 1570 2153 1581 2156
rect 1570 2113 1573 2153
rect 1586 2113 1589 2126
rect 1558 2103 1573 2106
rect 1530 2033 1565 2036
rect 1458 1613 1461 1646
rect 1458 1573 1461 1606
rect 1450 1553 1457 1556
rect 1430 1493 1437 1496
rect 1394 1403 1405 1406
rect 1370 1333 1389 1336
rect 1386 1326 1389 1333
rect 1378 1313 1381 1326
rect 1386 1323 1397 1326
rect 1402 1306 1405 1403
rect 1354 1303 1365 1306
rect 1298 1273 1333 1276
rect 1342 1293 1349 1296
rect 1274 1203 1277 1216
rect 1282 1196 1285 1226
rect 1290 1213 1293 1246
rect 1298 1203 1301 1273
rect 1314 1223 1333 1226
rect 1314 1216 1317 1223
rect 1306 1213 1317 1216
rect 1258 1093 1261 1116
rect 1274 1103 1277 1196
rect 1282 1193 1289 1196
rect 1266 1093 1277 1096
rect 1250 1043 1261 1046
rect 1250 1023 1253 1036
rect 1258 946 1261 1043
rect 1266 1013 1269 1093
rect 1286 1086 1289 1193
rect 1314 1146 1317 1206
rect 1322 1196 1325 1216
rect 1330 1213 1333 1223
rect 1322 1193 1329 1196
rect 1282 1083 1289 1086
rect 1298 1143 1317 1146
rect 1266 993 1269 1006
rect 1250 826 1253 946
rect 1258 943 1269 946
rect 1258 863 1261 936
rect 1250 823 1261 826
rect 1234 813 1253 816
rect 1258 806 1261 823
rect 1234 793 1237 806
rect 1242 803 1261 806
rect 1266 803 1269 943
rect 1274 893 1277 1016
rect 1282 913 1285 1083
rect 1290 933 1293 1056
rect 1298 993 1301 1143
rect 1298 913 1301 926
rect 1306 906 1309 1116
rect 1314 1083 1317 1136
rect 1326 1076 1329 1193
rect 1342 1156 1345 1293
rect 1362 1256 1365 1303
rect 1398 1303 1405 1306
rect 1354 1253 1365 1256
rect 1342 1153 1349 1156
rect 1346 1133 1349 1153
rect 1338 1083 1341 1126
rect 1354 1116 1357 1253
rect 1378 1203 1381 1226
rect 1386 1213 1389 1286
rect 1398 1246 1401 1303
rect 1394 1243 1401 1246
rect 1394 1206 1397 1243
rect 1402 1223 1405 1236
rect 1386 1203 1397 1206
rect 1370 1143 1373 1166
rect 1370 1123 1381 1126
rect 1346 1113 1365 1116
rect 1322 1073 1329 1076
rect 1314 1003 1317 1016
rect 1314 933 1317 996
rect 1322 926 1325 1073
rect 1378 1053 1381 1106
rect 1330 993 1333 1046
rect 1362 1043 1381 1046
rect 1354 1013 1357 1036
rect 1362 1023 1365 1043
rect 1338 1003 1365 1006
rect 1338 966 1341 1003
rect 1330 963 1341 966
rect 1330 933 1333 963
rect 1322 923 1333 926
rect 1338 923 1341 956
rect 1354 923 1357 996
rect 1290 903 1309 906
rect 1290 823 1293 903
rect 1322 896 1325 916
rect 1318 893 1325 896
rect 1318 836 1321 893
rect 1314 833 1321 836
rect 1314 823 1317 833
rect 1330 826 1333 923
rect 1322 823 1333 826
rect 1226 763 1233 766
rect 1218 743 1221 756
rect 1218 683 1221 726
rect 1230 686 1233 763
rect 1242 743 1245 803
rect 1242 693 1245 726
rect 1226 683 1233 686
rect 1226 663 1229 683
rect 1250 633 1253 776
rect 1258 716 1261 803
rect 1266 733 1269 756
rect 1258 713 1269 716
rect 1210 613 1229 616
rect 1226 593 1229 613
rect 1234 586 1237 616
rect 1198 583 1213 586
rect 1186 573 1197 576
rect 1170 533 1181 536
rect 1154 503 1157 516
rect 1170 453 1173 533
rect 1178 446 1181 526
rect 1194 513 1197 573
rect 1170 443 1181 446
rect 1170 413 1173 443
rect 1186 436 1189 506
rect 1202 496 1205 566
rect 1210 516 1213 583
rect 1226 583 1237 586
rect 1226 523 1229 583
rect 1250 563 1253 606
rect 1234 543 1237 556
rect 1234 526 1237 536
rect 1250 526 1253 556
rect 1234 523 1253 526
rect 1258 523 1261 706
rect 1266 613 1269 713
rect 1274 613 1277 816
rect 1298 743 1301 796
rect 1314 736 1317 746
rect 1282 683 1285 736
rect 1298 733 1317 736
rect 1322 733 1325 823
rect 1338 816 1341 836
rect 1330 813 1341 816
rect 1330 766 1333 813
rect 1338 793 1341 806
rect 1346 803 1349 886
rect 1354 853 1357 916
rect 1370 836 1373 1016
rect 1378 973 1381 1043
rect 1386 1023 1389 1203
rect 1386 956 1389 986
rect 1382 953 1389 956
rect 1382 886 1385 953
rect 1382 883 1389 886
rect 1370 833 1381 836
rect 1354 803 1357 816
rect 1362 773 1365 826
rect 1370 783 1373 826
rect 1378 806 1381 833
rect 1386 813 1389 883
rect 1394 853 1397 1176
rect 1402 916 1405 1196
rect 1410 1193 1413 1336
rect 1418 1166 1421 1336
rect 1426 1283 1429 1476
rect 1434 1226 1437 1493
rect 1442 1463 1445 1516
rect 1454 1456 1457 1553
rect 1450 1453 1457 1456
rect 1410 1163 1421 1166
rect 1426 1223 1437 1226
rect 1410 933 1413 1163
rect 1426 1156 1429 1223
rect 1434 1173 1437 1216
rect 1418 1153 1429 1156
rect 1418 1093 1421 1153
rect 1426 1133 1429 1146
rect 1418 943 1421 1046
rect 1426 926 1429 1126
rect 1434 1093 1437 1136
rect 1442 1066 1445 1406
rect 1450 1176 1453 1453
rect 1458 1393 1461 1406
rect 1458 1323 1461 1376
rect 1466 1316 1469 1856
rect 1474 1813 1477 1896
rect 1482 1806 1485 1906
rect 1490 1893 1493 1926
rect 1502 1886 1505 1973
rect 1530 1933 1533 2033
rect 1538 2013 1549 2016
rect 1498 1883 1505 1886
rect 1498 1816 1501 1883
rect 1474 1803 1485 1806
rect 1490 1813 1501 1816
rect 1474 1603 1477 1803
rect 1490 1753 1493 1813
rect 1498 1793 1501 1806
rect 1506 1803 1509 1846
rect 1482 1656 1485 1736
rect 1490 1713 1493 1726
rect 1498 1666 1501 1726
rect 1506 1723 1509 1736
rect 1514 1716 1517 1926
rect 1538 1923 1541 2013
rect 1546 1983 1549 1996
rect 1554 1926 1557 2026
rect 1562 2013 1565 2033
rect 1554 1923 1565 1926
rect 1522 1913 1557 1916
rect 1562 1906 1565 1923
rect 1558 1903 1565 1906
rect 1522 1763 1525 1856
rect 1546 1846 1549 1866
rect 1558 1846 1561 1903
rect 1570 1853 1573 2103
rect 1594 2033 1597 2136
rect 1602 2103 1605 2126
rect 1610 2016 1613 2126
rect 1618 2116 1621 2283
rect 1626 2143 1629 2166
rect 1634 2133 1637 2336
rect 1642 2313 1645 2336
rect 1650 2323 1653 2336
rect 1642 2213 1653 2216
rect 1658 2196 1661 2343
rect 1666 2303 1669 2353
rect 1682 2296 1685 2363
rect 1674 2293 1685 2296
rect 1650 2193 1661 2196
rect 1666 2193 1669 2206
rect 1618 2113 1629 2116
rect 1626 2046 1629 2113
rect 1602 2013 1613 2016
rect 1618 2043 1629 2046
rect 1618 2026 1621 2043
rect 1618 2023 1637 2026
rect 1610 1943 1613 2006
rect 1578 1923 1581 1936
rect 1586 1903 1589 1936
rect 1594 1933 1605 1936
rect 1618 1916 1621 2023
rect 1626 1963 1629 2006
rect 1634 2003 1637 2016
rect 1610 1913 1621 1916
rect 1538 1843 1549 1846
rect 1554 1843 1561 1846
rect 1610 1846 1613 1913
rect 1610 1843 1621 1846
rect 1538 1796 1541 1843
rect 1554 1806 1557 1843
rect 1562 1823 1605 1826
rect 1562 1813 1565 1823
rect 1570 1806 1573 1816
rect 1554 1803 1573 1806
rect 1538 1793 1549 1796
rect 1506 1713 1517 1716
rect 1522 1713 1525 1736
rect 1530 1733 1533 1776
rect 1546 1756 1549 1793
rect 1538 1753 1549 1756
rect 1506 1683 1509 1713
rect 1538 1706 1541 1753
rect 1522 1703 1541 1706
rect 1490 1663 1501 1666
rect 1482 1653 1493 1656
rect 1474 1493 1477 1596
rect 1474 1383 1477 1396
rect 1474 1333 1477 1366
rect 1458 1203 1461 1316
rect 1466 1313 1473 1316
rect 1470 1236 1473 1313
rect 1466 1233 1473 1236
rect 1450 1173 1461 1176
rect 1450 1133 1453 1166
rect 1458 1086 1461 1173
rect 1466 1103 1469 1233
rect 1434 1063 1445 1066
rect 1434 1043 1437 1063
rect 1434 993 1437 1006
rect 1418 923 1429 926
rect 1402 913 1421 916
rect 1402 903 1413 906
rect 1402 813 1405 896
rect 1378 803 1405 806
rect 1370 773 1389 776
rect 1370 766 1373 773
rect 1394 766 1397 796
rect 1330 763 1349 766
rect 1290 693 1293 726
rect 1266 573 1269 606
rect 1274 593 1277 606
rect 1282 546 1285 636
rect 1274 543 1285 546
rect 1210 513 1229 516
rect 1202 493 1221 496
rect 1178 396 1181 436
rect 1186 433 1197 436
rect 1186 413 1189 426
rect 1202 413 1205 466
rect 1170 393 1181 396
rect 1138 336 1141 346
rect 1130 333 1141 336
rect 1138 323 1141 333
rect 1170 326 1173 393
rect 1146 316 1149 326
rect 1170 323 1181 326
rect 1122 313 1149 316
rect 1178 303 1181 323
rect 1194 313 1197 406
rect 1210 366 1213 436
rect 1218 423 1221 493
rect 1226 413 1229 513
rect 1250 496 1253 516
rect 1258 503 1269 506
rect 1250 493 1261 496
rect 1210 363 1221 366
rect 1202 333 1205 346
rect 1218 303 1221 363
rect 1234 336 1237 436
rect 1250 416 1253 436
rect 1246 413 1253 416
rect 1246 356 1249 413
rect 1246 353 1253 356
rect 1234 333 1245 336
rect 1226 316 1229 326
rect 1242 323 1245 333
rect 1250 316 1253 353
rect 1226 313 1253 316
rect 1258 313 1261 493
rect 1266 446 1269 503
rect 1274 456 1277 543
rect 1282 463 1285 536
rect 1290 533 1293 616
rect 1298 613 1301 733
rect 1298 593 1301 606
rect 1290 473 1293 526
rect 1298 513 1301 586
rect 1306 536 1309 726
rect 1314 723 1325 726
rect 1314 643 1317 723
rect 1330 713 1333 756
rect 1314 543 1317 586
rect 1306 533 1317 536
rect 1314 523 1317 533
rect 1322 503 1325 656
rect 1330 613 1333 706
rect 1338 693 1341 746
rect 1346 653 1349 763
rect 1362 763 1373 766
rect 1386 763 1397 766
rect 1354 723 1357 746
rect 1362 726 1365 763
rect 1370 733 1373 756
rect 1362 723 1381 726
rect 1362 666 1365 723
rect 1354 663 1365 666
rect 1330 583 1341 586
rect 1346 583 1349 606
rect 1338 533 1341 583
rect 1354 576 1357 663
rect 1346 573 1357 576
rect 1330 513 1333 526
rect 1274 453 1285 456
rect 1266 443 1301 446
rect 1266 413 1269 443
rect 1282 423 1285 436
rect 1290 403 1293 426
rect 1298 413 1301 443
rect 1306 403 1309 486
rect 1314 393 1317 406
rect 1322 373 1325 456
rect 1346 413 1349 573
rect 1354 533 1357 566
rect 1362 553 1365 606
rect 1370 603 1373 616
rect 1378 603 1381 636
rect 1386 443 1389 763
rect 1394 703 1397 736
rect 1402 733 1405 803
rect 1410 793 1413 903
rect 1418 726 1421 913
rect 1426 876 1429 923
rect 1434 893 1437 916
rect 1426 873 1437 876
rect 1426 813 1429 826
rect 1426 743 1429 756
rect 1434 743 1437 873
rect 1442 833 1445 1056
rect 1450 923 1453 1086
rect 1458 1083 1465 1086
rect 1462 1026 1465 1083
rect 1458 1023 1465 1026
rect 1458 986 1461 1023
rect 1474 1013 1477 1216
rect 1482 1193 1485 1646
rect 1490 1603 1493 1653
rect 1522 1636 1525 1703
rect 1490 1583 1493 1596
rect 1490 1313 1493 1576
rect 1498 1403 1501 1626
rect 1506 1396 1509 1636
rect 1514 1633 1525 1636
rect 1514 1596 1517 1633
rect 1546 1616 1549 1726
rect 1554 1723 1557 1796
rect 1578 1783 1581 1806
rect 1562 1706 1565 1766
rect 1586 1746 1589 1816
rect 1602 1813 1605 1823
rect 1594 1753 1597 1806
rect 1618 1786 1621 1843
rect 1626 1803 1629 1926
rect 1634 1886 1637 1976
rect 1650 1956 1653 2193
rect 1674 2186 1677 2293
rect 1694 2246 1697 2393
rect 1694 2243 1701 2246
rect 1698 2223 1701 2243
rect 1666 2183 1677 2186
rect 1666 1966 1669 2183
rect 1690 2143 1701 2146
rect 1682 2023 1685 2126
rect 1690 2083 1693 2136
rect 1698 2023 1701 2143
rect 1706 2016 1709 2446
rect 1714 2383 1717 2426
rect 1722 2323 1725 2426
rect 1730 2356 1733 2493
rect 1738 2413 1741 2436
rect 1738 2373 1741 2406
rect 1730 2353 1737 2356
rect 1734 2296 1737 2353
rect 1746 2313 1749 2366
rect 1754 2353 1757 2416
rect 1762 2313 1765 2533
rect 1778 2516 1781 2716
rect 1794 2546 1797 2793
rect 1810 2733 1813 2746
rect 1818 2706 1821 2726
rect 1810 2703 1821 2706
rect 1810 2636 1813 2703
rect 1810 2633 1821 2636
rect 1818 2613 1821 2633
rect 1826 2593 1829 2803
rect 1842 2746 1845 2893
rect 1850 2883 1869 2886
rect 1858 2823 1861 2846
rect 1866 2813 1869 2883
rect 1838 2743 1845 2746
rect 1838 2666 1841 2743
rect 1850 2673 1853 2736
rect 1838 2663 1845 2666
rect 1834 2603 1837 2636
rect 1794 2543 1801 2546
rect 1774 2513 1781 2516
rect 1774 2456 1777 2513
rect 1786 2463 1789 2536
rect 1798 2456 1801 2543
rect 1810 2523 1813 2536
rect 1818 2533 1821 2546
rect 1774 2453 1781 2456
rect 1770 2333 1773 2386
rect 1734 2293 1749 2296
rect 1714 2213 1717 2246
rect 1722 2213 1725 2226
rect 1746 2156 1749 2293
rect 1770 2223 1773 2256
rect 1770 2203 1773 2216
rect 1730 2153 1749 2156
rect 1730 2136 1733 2153
rect 1714 2033 1717 2136
rect 1722 2103 1725 2136
rect 1730 2133 1741 2136
rect 1730 2113 1733 2126
rect 1722 2023 1725 2046
rect 1682 2013 1709 2016
rect 1674 2003 1685 2006
rect 1682 1983 1685 2003
rect 1666 1963 1677 1966
rect 1650 1953 1661 1956
rect 1642 1913 1645 1926
rect 1650 1903 1653 1936
rect 1658 1886 1661 1953
rect 1674 1896 1677 1963
rect 1722 1946 1725 2006
rect 1722 1943 1729 1946
rect 1706 1933 1717 1936
rect 1634 1883 1645 1886
rect 1642 1786 1645 1883
rect 1654 1883 1661 1886
rect 1666 1893 1677 1896
rect 1698 1893 1701 1926
rect 1654 1796 1657 1883
rect 1666 1873 1669 1893
rect 1714 1843 1717 1916
rect 1726 1856 1729 1943
rect 1722 1853 1729 1856
rect 1722 1836 1725 1853
rect 1714 1833 1725 1836
rect 1666 1806 1669 1826
rect 1666 1803 1677 1806
rect 1654 1793 1661 1796
rect 1602 1783 1621 1786
rect 1626 1783 1645 1786
rect 1602 1746 1605 1783
rect 1586 1743 1605 1746
rect 1570 1713 1573 1726
rect 1578 1716 1581 1736
rect 1578 1713 1597 1716
rect 1562 1703 1573 1706
rect 1570 1646 1573 1703
rect 1570 1643 1581 1646
rect 1522 1613 1549 1616
rect 1522 1603 1525 1613
rect 1514 1593 1525 1596
rect 1514 1523 1517 1536
rect 1498 1393 1509 1396
rect 1498 1286 1501 1393
rect 1514 1386 1517 1516
rect 1522 1473 1525 1593
rect 1530 1523 1533 1546
rect 1490 1283 1501 1286
rect 1506 1383 1517 1386
rect 1490 1196 1493 1283
rect 1506 1276 1509 1383
rect 1522 1333 1525 1406
rect 1530 1386 1533 1416
rect 1538 1413 1541 1606
rect 1554 1513 1557 1626
rect 1570 1583 1573 1606
rect 1562 1523 1565 1536
rect 1546 1403 1549 1416
rect 1562 1403 1565 1476
rect 1530 1383 1541 1386
rect 1522 1313 1525 1326
rect 1530 1283 1533 1356
rect 1498 1273 1509 1276
rect 1498 1203 1501 1273
rect 1538 1266 1541 1383
rect 1546 1276 1549 1376
rect 1570 1356 1573 1416
rect 1578 1413 1581 1643
rect 1586 1433 1589 1713
rect 1602 1696 1605 1743
rect 1610 1703 1613 1776
rect 1594 1693 1605 1696
rect 1594 1593 1597 1606
rect 1602 1526 1605 1693
rect 1626 1623 1629 1783
rect 1650 1716 1653 1736
rect 1642 1713 1653 1716
rect 1642 1626 1645 1713
rect 1642 1623 1653 1626
rect 1610 1573 1613 1606
rect 1626 1543 1629 1606
rect 1650 1603 1653 1623
rect 1658 1536 1661 1793
rect 1674 1746 1677 1803
rect 1698 1763 1701 1806
rect 1666 1743 1677 1746
rect 1706 1743 1709 1806
rect 1666 1713 1669 1743
rect 1690 1693 1693 1726
rect 1698 1713 1701 1726
rect 1674 1606 1677 1626
rect 1682 1613 1685 1636
rect 1594 1523 1605 1526
rect 1554 1333 1557 1356
rect 1562 1353 1573 1356
rect 1546 1273 1557 1276
rect 1506 1263 1549 1266
rect 1490 1193 1501 1196
rect 1482 1053 1485 1136
rect 1490 1013 1493 1106
rect 1498 1083 1501 1193
rect 1506 1123 1509 1263
rect 1514 1163 1517 1196
rect 1522 1193 1525 1256
rect 1506 1016 1509 1096
rect 1514 1063 1517 1136
rect 1522 1103 1525 1126
rect 1506 1013 1513 1016
rect 1466 1001 1477 1004
rect 1458 983 1465 986
rect 1462 916 1465 983
rect 1474 953 1477 1001
rect 1458 913 1465 916
rect 1402 723 1421 726
rect 1394 603 1397 656
rect 1394 583 1397 596
rect 1402 556 1405 616
rect 1410 603 1413 723
rect 1426 613 1429 726
rect 1434 693 1437 726
rect 1442 696 1445 806
rect 1450 753 1453 866
rect 1458 816 1461 913
rect 1458 813 1469 816
rect 1458 793 1461 806
rect 1458 766 1461 786
rect 1466 773 1469 813
rect 1458 763 1469 766
rect 1450 733 1453 746
rect 1466 733 1469 763
rect 1474 716 1477 946
rect 1482 933 1485 1006
rect 1482 813 1485 836
rect 1490 813 1493 956
rect 1498 806 1501 1006
rect 1510 936 1513 1013
rect 1522 943 1525 1086
rect 1530 1053 1533 1136
rect 1538 1123 1541 1216
rect 1546 1133 1549 1263
rect 1554 1126 1557 1273
rect 1546 1123 1557 1126
rect 1510 933 1517 936
rect 1506 913 1509 926
rect 1514 906 1517 933
rect 1470 713 1477 716
rect 1482 803 1501 806
rect 1506 903 1517 906
rect 1442 693 1461 696
rect 1442 623 1445 686
rect 1434 603 1445 606
rect 1394 553 1405 556
rect 1394 523 1397 553
rect 1410 483 1413 536
rect 1418 513 1421 576
rect 1450 566 1453 606
rect 1458 573 1461 693
rect 1470 566 1473 713
rect 1442 563 1453 566
rect 1458 563 1473 566
rect 1426 523 1429 556
rect 1434 533 1445 536
rect 1354 403 1365 406
rect 1354 383 1357 403
rect 1362 393 1373 396
rect 1314 353 1333 356
rect 1314 343 1317 353
rect 1330 333 1333 353
rect 1378 336 1381 406
rect 1370 333 1381 336
rect 1266 303 1269 326
rect 1098 253 1141 256
rect 1034 163 1045 166
rect 930 93 933 126
rect 1010 113 1013 126
rect 1042 86 1045 163
rect 1066 123 1069 236
rect 1098 213 1101 253
rect 1138 213 1141 253
rect 1114 186 1117 206
rect 1242 203 1245 226
rect 1266 216 1269 286
rect 1258 213 1269 216
rect 1234 193 1245 196
rect 1106 183 1117 186
rect 1106 133 1109 183
rect 1218 133 1221 146
rect 1034 83 1045 86
rect 1090 86 1093 126
rect 1130 86 1133 126
rect 1218 96 1221 126
rect 1226 113 1229 126
rect 1234 106 1237 136
rect 1242 123 1245 193
rect 1258 133 1261 146
rect 1266 136 1269 213
rect 1274 203 1277 216
rect 1282 203 1285 256
rect 1290 213 1293 296
rect 1370 283 1373 333
rect 1378 273 1381 326
rect 1410 323 1413 426
rect 1426 423 1429 516
rect 1426 386 1429 416
rect 1434 413 1437 526
rect 1442 403 1445 533
rect 1450 453 1453 536
rect 1458 436 1461 563
rect 1482 546 1485 803
rect 1490 733 1493 786
rect 1498 726 1501 736
rect 1490 723 1501 726
rect 1490 666 1493 706
rect 1498 683 1501 723
rect 1506 686 1509 903
rect 1522 883 1525 936
rect 1530 933 1533 956
rect 1538 876 1541 1106
rect 1522 873 1541 876
rect 1514 803 1517 846
rect 1522 813 1525 873
rect 1514 743 1517 756
rect 1530 736 1533 836
rect 1538 813 1541 866
rect 1546 833 1549 1123
rect 1562 1103 1565 1353
rect 1578 1346 1581 1406
rect 1586 1373 1589 1416
rect 1594 1383 1597 1523
rect 1602 1503 1605 1516
rect 1610 1493 1613 1536
rect 1618 1533 1661 1536
rect 1666 1603 1677 1606
rect 1602 1403 1605 1416
rect 1570 1343 1581 1346
rect 1570 1313 1573 1343
rect 1578 1236 1581 1336
rect 1594 1323 1597 1346
rect 1610 1343 1613 1406
rect 1578 1233 1589 1236
rect 1570 1093 1573 1216
rect 1578 1203 1581 1226
rect 1578 1183 1581 1196
rect 1554 803 1557 1056
rect 1562 896 1565 1086
rect 1570 993 1573 1026
rect 1578 1013 1581 1126
rect 1586 1083 1589 1233
rect 1602 1223 1605 1236
rect 1618 1216 1621 1533
rect 1642 1506 1645 1526
rect 1650 1523 1661 1526
rect 1666 1513 1669 1603
rect 1682 1573 1685 1606
rect 1698 1593 1701 1626
rect 1706 1573 1709 1706
rect 1674 1543 1685 1546
rect 1674 1506 1677 1543
rect 1682 1533 1701 1536
rect 1682 1523 1685 1533
rect 1642 1503 1677 1506
rect 1698 1473 1701 1516
rect 1714 1506 1717 1833
rect 1722 1783 1725 1826
rect 1738 1803 1741 2133
rect 1778 2056 1781 2453
rect 1794 2453 1801 2456
rect 1794 2376 1797 2453
rect 1810 2413 1813 2486
rect 1818 2393 1821 2526
rect 1826 2453 1829 2526
rect 1842 2516 1845 2663
rect 1858 2616 1861 2786
rect 1882 2776 1885 2893
rect 1898 2876 1901 2933
rect 1894 2873 1901 2876
rect 1894 2796 1897 2873
rect 1894 2793 1901 2796
rect 1882 2773 1893 2776
rect 1874 2716 1877 2736
rect 1882 2723 1885 2756
rect 1890 2716 1893 2773
rect 1870 2713 1877 2716
rect 1882 2713 1893 2716
rect 1870 2636 1873 2713
rect 1882 2703 1885 2713
rect 1870 2633 1877 2636
rect 1858 2613 1865 2616
rect 1850 2533 1853 2606
rect 1862 2556 1865 2613
rect 1858 2553 1865 2556
rect 1874 2553 1877 2633
rect 1858 2533 1861 2553
rect 1882 2523 1885 2666
rect 1890 2603 1893 2626
rect 1842 2513 1853 2516
rect 1794 2373 1805 2376
rect 1786 2333 1789 2346
rect 1802 2226 1805 2373
rect 1834 2313 1837 2476
rect 1850 2446 1853 2513
rect 1890 2506 1893 2526
rect 1898 2513 1901 2793
rect 1906 2776 1909 2926
rect 1914 2923 1917 2996
rect 1922 2803 1925 2926
rect 1930 2873 1933 3026
rect 1970 3016 1973 3113
rect 1938 3003 1941 3016
rect 1946 2996 1949 3016
rect 1970 3013 1981 3016
rect 1946 2993 1957 2996
rect 1954 2946 1957 2993
rect 1978 2946 1981 3013
rect 1986 3003 1989 3036
rect 1994 2993 1997 3133
rect 2010 3013 2013 3086
rect 2026 3053 2029 3223
rect 2042 3196 2045 3206
rect 2058 3203 2061 3216
rect 2074 3196 2077 3206
rect 2042 3193 2077 3196
rect 2082 3163 2085 3216
rect 2090 3183 2093 3216
rect 2102 3156 2105 3233
rect 2058 3143 2061 3156
rect 2098 3153 2105 3156
rect 2002 2983 2005 3006
rect 1946 2943 1957 2946
rect 1970 2943 1981 2946
rect 1906 2773 1933 2776
rect 1914 2726 1917 2736
rect 1906 2723 1917 2726
rect 1922 2723 1925 2736
rect 1906 2713 1909 2723
rect 1914 2703 1917 2716
rect 1930 2656 1933 2773
rect 1906 2653 1933 2656
rect 1906 2613 1909 2653
rect 1922 2613 1925 2636
rect 1842 2443 1853 2446
rect 1882 2503 1893 2506
rect 1882 2446 1885 2503
rect 1882 2443 1893 2446
rect 1842 2296 1845 2443
rect 1890 2426 1893 2443
rect 1850 2403 1853 2426
rect 1890 2423 1901 2426
rect 1858 2413 1893 2416
rect 1838 2293 1845 2296
rect 1802 2223 1829 2226
rect 1794 2213 1813 2216
rect 1786 2193 1789 2206
rect 1802 2203 1813 2206
rect 1826 2186 1829 2223
rect 1838 2196 1841 2293
rect 1838 2193 1845 2196
rect 1810 2183 1829 2186
rect 1810 2086 1813 2183
rect 1834 2133 1837 2176
rect 1842 2143 1845 2193
rect 1850 2176 1853 2396
rect 1858 2333 1861 2413
rect 1898 2406 1901 2423
rect 1866 2383 1869 2406
rect 1874 2403 1901 2406
rect 1874 2393 1877 2403
rect 1858 2223 1861 2306
rect 1866 2223 1877 2226
rect 1882 2206 1885 2336
rect 1898 2323 1901 2336
rect 1858 2196 1861 2206
rect 1878 2203 1885 2206
rect 1858 2193 1869 2196
rect 1850 2173 1857 2176
rect 1834 2093 1837 2116
rect 1810 2083 1829 2086
rect 1826 2066 1829 2083
rect 1826 2063 1833 2066
rect 1770 2053 1781 2056
rect 1754 1936 1757 2036
rect 1770 1966 1773 2053
rect 1770 1963 1781 1966
rect 1786 1963 1789 2046
rect 1818 2023 1821 2056
rect 1830 2016 1833 2063
rect 1842 2043 1845 2126
rect 1854 2116 1857 2173
rect 1866 2133 1869 2186
rect 1878 2146 1881 2203
rect 1874 2143 1881 2146
rect 1854 2113 1861 2116
rect 1826 2013 1833 2016
rect 1746 1933 1757 1936
rect 1746 1913 1749 1933
rect 1754 1923 1765 1926
rect 1770 1923 1773 1946
rect 1778 1906 1781 1963
rect 1826 1936 1829 2013
rect 1850 1973 1853 2026
rect 1858 2016 1861 2113
rect 1858 2013 1865 2016
rect 1794 1923 1797 1936
rect 1818 1933 1829 1936
rect 1770 1903 1781 1906
rect 1746 1746 1749 1856
rect 1770 1836 1773 1903
rect 1770 1833 1781 1836
rect 1762 1793 1765 1816
rect 1778 1806 1781 1833
rect 1786 1823 1789 1906
rect 1818 1846 1821 1933
rect 1850 1926 1853 1956
rect 1834 1863 1837 1926
rect 1842 1923 1853 1926
rect 1794 1826 1797 1846
rect 1818 1843 1829 1846
rect 1794 1823 1805 1826
rect 1742 1743 1749 1746
rect 1722 1696 1725 1716
rect 1722 1693 1733 1696
rect 1730 1646 1733 1693
rect 1742 1686 1745 1743
rect 1754 1693 1757 1736
rect 1762 1713 1765 1766
rect 1770 1723 1773 1806
rect 1778 1803 1785 1806
rect 1782 1736 1785 1803
rect 1802 1776 1805 1823
rect 1778 1733 1785 1736
rect 1794 1773 1805 1776
rect 1778 1713 1781 1733
rect 1794 1716 1797 1773
rect 1802 1723 1805 1756
rect 1818 1726 1821 1746
rect 1810 1723 1821 1726
rect 1794 1713 1805 1716
rect 1742 1683 1749 1686
rect 1722 1643 1733 1646
rect 1722 1596 1725 1643
rect 1738 1613 1741 1626
rect 1722 1593 1733 1596
rect 1714 1503 1721 1506
rect 1626 1363 1629 1466
rect 1674 1403 1677 1436
rect 1706 1423 1709 1496
rect 1718 1416 1721 1503
rect 1682 1413 1701 1416
rect 1626 1313 1629 1326
rect 1634 1233 1637 1336
rect 1642 1323 1645 1336
rect 1650 1323 1653 1386
rect 1642 1216 1645 1286
rect 1650 1223 1661 1226
rect 1666 1223 1669 1266
rect 1674 1226 1677 1336
rect 1690 1333 1693 1356
rect 1698 1333 1701 1413
rect 1714 1413 1721 1416
rect 1714 1353 1717 1413
rect 1730 1346 1733 1593
rect 1746 1576 1749 1683
rect 1762 1583 1765 1626
rect 1770 1603 1773 1636
rect 1778 1613 1781 1656
rect 1786 1613 1797 1616
rect 1742 1573 1749 1576
rect 1742 1516 1745 1573
rect 1754 1563 1765 1566
rect 1754 1523 1757 1563
rect 1802 1543 1805 1713
rect 1826 1583 1829 1843
rect 1834 1816 1837 1826
rect 1834 1813 1845 1816
rect 1850 1796 1853 1906
rect 1842 1793 1853 1796
rect 1842 1636 1845 1793
rect 1862 1786 1865 2013
rect 1874 1793 1877 2143
rect 1882 2123 1885 2136
rect 1890 2123 1893 2206
rect 1890 2033 1901 2036
rect 1890 2013 1893 2033
rect 1906 2016 1909 2566
rect 1914 2323 1917 2606
rect 1930 2603 1933 2626
rect 1938 2613 1941 2926
rect 1946 2923 1949 2943
rect 1954 2816 1957 2926
rect 1970 2836 1973 2943
rect 1986 2933 1997 2936
rect 1970 2833 1977 2836
rect 1954 2813 1965 2816
rect 1946 2683 1949 2806
rect 1962 2736 1965 2813
rect 1974 2756 1977 2833
rect 1974 2753 1981 2756
rect 1954 2733 1965 2736
rect 1978 2733 1981 2753
rect 1954 2666 1957 2733
rect 1950 2663 1957 2666
rect 1950 2576 1953 2663
rect 1962 2586 1965 2716
rect 1978 2706 1981 2726
rect 1974 2703 1981 2706
rect 1974 2616 1977 2703
rect 1986 2686 1989 2933
rect 2010 2923 2013 3006
rect 2050 2936 2053 3116
rect 2074 3103 2077 3126
rect 2082 2996 2085 3026
rect 2074 2993 2085 2996
rect 1994 2823 1997 2866
rect 2026 2843 2029 2926
rect 2010 2803 2013 2826
rect 2002 2733 2005 2766
rect 1994 2713 1997 2726
rect 2010 2703 2013 2726
rect 2026 2723 2029 2756
rect 1986 2683 1997 2686
rect 1974 2613 1981 2616
rect 1978 2596 1981 2613
rect 1986 2603 1989 2676
rect 1978 2593 1989 2596
rect 1962 2583 1973 2586
rect 1950 2573 1957 2576
rect 1922 2333 1925 2536
rect 1930 2413 1933 2536
rect 1946 2403 1949 2456
rect 1930 2326 1933 2346
rect 1954 2326 1957 2573
rect 1970 2446 1973 2583
rect 1970 2443 1981 2446
rect 1970 2413 1973 2426
rect 1962 2343 1965 2406
rect 1978 2396 1981 2443
rect 1974 2393 1981 2396
rect 1974 2326 1977 2393
rect 1930 2323 1937 2326
rect 1922 2213 1925 2296
rect 1934 2236 1937 2323
rect 1930 2233 1937 2236
rect 1930 2206 1933 2233
rect 1922 2203 1933 2206
rect 1922 2086 1925 2203
rect 1938 2193 1941 2216
rect 1946 2186 1949 2326
rect 1954 2323 1965 2326
rect 1974 2323 1981 2326
rect 1962 2236 1965 2323
rect 1978 2303 1981 2323
rect 1986 2293 1989 2593
rect 1994 2506 1997 2683
rect 2002 2643 2029 2646
rect 2002 2613 2005 2643
rect 2018 2623 2021 2636
rect 2026 2613 2029 2643
rect 2018 2583 2021 2606
rect 2026 2566 2029 2606
rect 2002 2563 2029 2566
rect 2002 2523 2005 2563
rect 2010 2533 2013 2546
rect 2034 2523 2037 2936
rect 2042 2933 2053 2936
rect 2042 2516 2045 2933
rect 2050 2903 2053 2926
rect 2058 2923 2061 2946
rect 2074 2906 2077 2993
rect 2074 2903 2085 2906
rect 2050 2813 2053 2826
rect 2018 2513 2045 2516
rect 1994 2503 2009 2506
rect 2006 2446 2009 2503
rect 2018 2456 2021 2513
rect 2018 2453 2025 2456
rect 1994 2403 1997 2446
rect 2006 2443 2013 2446
rect 2002 2403 2005 2426
rect 2010 2396 2013 2443
rect 1994 2393 2013 2396
rect 1994 2343 1997 2393
rect 2022 2386 2025 2453
rect 2018 2383 2025 2386
rect 2018 2336 2021 2383
rect 2002 2333 2021 2336
rect 1938 2183 1949 2186
rect 1954 2233 1965 2236
rect 1938 2113 1941 2183
rect 1946 2123 1949 2166
rect 1946 2103 1949 2116
rect 1954 2086 1957 2233
rect 1922 2083 1933 2086
rect 1898 2013 1909 2016
rect 1890 1816 1893 2006
rect 1906 1913 1909 1976
rect 1914 1836 1917 2046
rect 1930 1966 1933 2083
rect 1946 2083 1957 2086
rect 1962 2083 1965 2206
rect 1970 2183 1973 2216
rect 1986 2193 1989 2266
rect 1970 2096 1973 2116
rect 1986 2113 1989 2136
rect 1970 2093 1981 2096
rect 1946 1996 1949 2083
rect 1962 2003 1965 2046
rect 1978 2036 1981 2093
rect 1970 2033 1981 2036
rect 1970 2013 1973 2033
rect 1994 2023 1997 2316
rect 1946 1993 1957 1996
rect 1922 1963 1933 1966
rect 1922 1943 1925 1963
rect 1954 1946 1957 1993
rect 1954 1943 1961 1946
rect 1922 1926 1925 1936
rect 1922 1923 1941 1926
rect 1946 1906 1949 1936
rect 1938 1903 1949 1906
rect 1914 1833 1925 1836
rect 1886 1813 1893 1816
rect 1858 1783 1865 1786
rect 1858 1756 1861 1783
rect 1854 1753 1861 1756
rect 1854 1696 1857 1753
rect 1866 1733 1869 1746
rect 1866 1703 1869 1716
rect 1854 1693 1861 1696
rect 1834 1633 1845 1636
rect 1762 1523 1765 1536
rect 1742 1513 1749 1516
rect 1722 1343 1733 1346
rect 1682 1313 1685 1326
rect 1698 1293 1701 1326
rect 1674 1223 1717 1226
rect 1658 1216 1661 1223
rect 1722 1216 1725 1343
rect 1614 1213 1621 1216
rect 1614 1146 1617 1213
rect 1626 1193 1629 1206
rect 1634 1196 1637 1216
rect 1642 1213 1653 1216
rect 1658 1213 1677 1216
rect 1634 1193 1641 1196
rect 1614 1143 1621 1146
rect 1594 1123 1597 1136
rect 1570 913 1573 936
rect 1562 893 1569 896
rect 1566 806 1569 893
rect 1578 823 1581 936
rect 1586 863 1589 1046
rect 1594 1023 1597 1116
rect 1602 1103 1605 1126
rect 1610 1093 1613 1126
rect 1618 1076 1621 1143
rect 1614 1073 1621 1076
rect 1602 983 1605 1006
rect 1614 976 1617 1073
rect 1602 973 1617 976
rect 1594 923 1597 936
rect 1566 803 1581 806
rect 1562 793 1573 796
rect 1578 786 1581 803
rect 1570 783 1581 786
rect 1514 733 1533 736
rect 1514 693 1517 733
rect 1522 696 1525 726
rect 1530 703 1533 726
rect 1522 693 1533 696
rect 1506 683 1525 686
rect 1490 663 1517 666
rect 1490 613 1493 656
rect 1490 553 1493 606
rect 1466 543 1477 546
rect 1482 543 1493 546
rect 1466 443 1469 536
rect 1490 523 1493 543
rect 1498 506 1501 616
rect 1506 583 1509 606
rect 1514 556 1517 663
rect 1522 603 1525 683
rect 1458 433 1469 436
rect 1458 393 1461 406
rect 1466 396 1469 433
rect 1474 403 1477 506
rect 1494 503 1501 506
rect 1506 553 1517 556
rect 1482 413 1485 446
rect 1494 436 1497 503
rect 1494 433 1501 436
rect 1498 413 1501 433
rect 1506 423 1509 553
rect 1530 546 1533 686
rect 1538 603 1541 736
rect 1546 723 1549 766
rect 1546 693 1549 716
rect 1554 676 1557 756
rect 1550 673 1557 676
rect 1550 616 1553 673
rect 1546 613 1553 616
rect 1514 543 1533 546
rect 1514 473 1517 543
rect 1522 523 1525 536
rect 1530 506 1533 536
rect 1546 526 1549 613
rect 1554 583 1557 596
rect 1554 533 1557 566
rect 1562 536 1565 766
rect 1570 563 1573 783
rect 1586 743 1589 826
rect 1594 813 1597 826
rect 1602 793 1605 973
rect 1626 966 1629 1176
rect 1638 1026 1641 1193
rect 1650 1106 1653 1213
rect 1674 1203 1677 1213
rect 1698 1213 1725 1216
rect 1658 1116 1661 1126
rect 1666 1123 1669 1166
rect 1674 1143 1693 1146
rect 1690 1133 1693 1143
rect 1658 1113 1669 1116
rect 1690 1106 1693 1116
rect 1650 1103 1693 1106
rect 1650 1053 1653 1103
rect 1698 1046 1701 1213
rect 1746 1206 1749 1513
rect 1794 1446 1797 1516
rect 1834 1466 1837 1633
rect 1842 1573 1845 1626
rect 1850 1596 1853 1616
rect 1858 1613 1861 1693
rect 1874 1643 1877 1736
rect 1886 1716 1889 1813
rect 1886 1713 1893 1716
rect 1898 1713 1901 1806
rect 1906 1783 1909 1826
rect 1922 1716 1925 1833
rect 1938 1786 1941 1903
rect 1958 1896 1961 1943
rect 1954 1893 1961 1896
rect 1938 1783 1949 1786
rect 1946 1763 1949 1783
rect 1914 1713 1925 1716
rect 1890 1693 1893 1713
rect 1874 1616 1877 1636
rect 1874 1613 1885 1616
rect 1890 1613 1901 1616
rect 1850 1593 1857 1596
rect 1866 1593 1869 1606
rect 1854 1546 1857 1593
rect 1874 1586 1877 1606
rect 1866 1583 1877 1586
rect 1890 1556 1893 1606
rect 1850 1543 1857 1546
rect 1874 1553 1893 1556
rect 1850 1466 1853 1543
rect 1834 1463 1845 1466
rect 1850 1463 1861 1466
rect 1786 1443 1797 1446
rect 1762 1413 1765 1426
rect 1786 1396 1789 1443
rect 1810 1423 1813 1436
rect 1786 1393 1797 1396
rect 1794 1373 1797 1393
rect 1802 1353 1805 1416
rect 1810 1383 1813 1406
rect 1802 1323 1805 1336
rect 1810 1333 1813 1346
rect 1818 1333 1821 1446
rect 1842 1423 1845 1463
rect 1826 1396 1829 1416
rect 1850 1403 1853 1456
rect 1826 1393 1845 1396
rect 1794 1293 1797 1316
rect 1770 1253 1781 1256
rect 1770 1213 1773 1253
rect 1778 1213 1797 1216
rect 1706 1203 1749 1206
rect 1706 1106 1709 1203
rect 1714 1123 1717 1176
rect 1738 1136 1741 1186
rect 1722 1133 1741 1136
rect 1706 1103 1717 1106
rect 1694 1043 1701 1046
rect 1618 963 1629 966
rect 1634 1023 1641 1026
rect 1658 1026 1661 1036
rect 1658 1023 1685 1026
rect 1578 733 1605 736
rect 1578 606 1581 666
rect 1594 663 1597 726
rect 1602 723 1605 733
rect 1602 653 1605 716
rect 1594 623 1597 636
rect 1586 613 1597 616
rect 1602 613 1605 636
rect 1610 606 1613 926
rect 1618 923 1621 963
rect 1634 923 1637 1023
rect 1666 1013 1685 1016
rect 1642 916 1645 1006
rect 1658 996 1661 1006
rect 1682 1003 1685 1013
rect 1658 993 1677 996
rect 1650 923 1653 986
rect 1642 913 1653 916
rect 1618 753 1621 866
rect 1626 863 1637 866
rect 1626 823 1629 863
rect 1650 846 1653 913
rect 1658 876 1661 976
rect 1674 913 1677 993
rect 1694 966 1697 1043
rect 1714 1036 1717 1103
rect 1738 1063 1741 1116
rect 1754 1053 1757 1126
rect 1706 1033 1717 1036
rect 1694 963 1701 966
rect 1698 943 1701 963
rect 1658 873 1669 876
rect 1642 843 1653 846
rect 1634 813 1637 826
rect 1634 773 1637 806
rect 1642 766 1645 843
rect 1626 763 1645 766
rect 1618 693 1621 736
rect 1626 733 1629 763
rect 1626 673 1629 726
rect 1634 703 1637 736
rect 1642 633 1645 756
rect 1650 716 1653 836
rect 1658 823 1661 866
rect 1666 856 1669 873
rect 1666 853 1673 856
rect 1658 723 1661 796
rect 1670 766 1673 853
rect 1682 796 1685 916
rect 1706 853 1709 1033
rect 1714 993 1717 1016
rect 1722 1013 1733 1016
rect 1714 923 1717 966
rect 1730 923 1733 946
rect 1738 906 1741 1026
rect 1754 1003 1757 1046
rect 1762 1033 1765 1206
rect 1802 1203 1805 1306
rect 1770 1133 1773 1166
rect 1770 1093 1773 1116
rect 1786 1063 1789 1126
rect 1794 1123 1797 1156
rect 1810 1126 1813 1236
rect 1818 1166 1821 1286
rect 1826 1203 1829 1326
rect 1834 1316 1837 1336
rect 1834 1313 1845 1316
rect 1842 1266 1845 1313
rect 1834 1263 1845 1266
rect 1834 1233 1837 1263
rect 1858 1246 1861 1463
rect 1866 1333 1869 1456
rect 1874 1403 1877 1553
rect 1882 1533 1893 1536
rect 1906 1533 1909 1556
rect 1890 1523 1909 1526
rect 1882 1396 1885 1476
rect 1906 1466 1909 1516
rect 1914 1473 1917 1713
rect 1930 1613 1933 1686
rect 1922 1503 1925 1606
rect 1930 1533 1933 1556
rect 1874 1393 1885 1396
rect 1890 1463 1909 1466
rect 1866 1303 1869 1326
rect 1842 1243 1861 1246
rect 1842 1176 1845 1243
rect 1874 1216 1877 1393
rect 1890 1366 1893 1463
rect 1914 1413 1917 1426
rect 1882 1363 1893 1366
rect 1882 1283 1885 1363
rect 1890 1333 1901 1336
rect 1890 1303 1893 1333
rect 1922 1323 1925 1416
rect 1930 1333 1933 1476
rect 1906 1313 1917 1316
rect 1938 1313 1941 1696
rect 1946 1663 1949 1746
rect 1946 1613 1949 1636
rect 1954 1596 1957 1893
rect 1962 1803 1965 1816
rect 1962 1676 1965 1736
rect 1970 1693 1973 2006
rect 1978 1966 1981 1986
rect 1978 1963 1989 1966
rect 1986 1896 1989 1963
rect 1978 1893 1989 1896
rect 1962 1673 1973 1676
rect 1970 1633 1973 1673
rect 1978 1616 1981 1893
rect 1986 1803 1989 1826
rect 1994 1813 1997 1876
rect 1986 1713 1989 1726
rect 1994 1723 1997 1766
rect 2002 1706 2005 2333
rect 2010 2243 2013 2326
rect 2026 2316 2029 2356
rect 2018 2313 2029 2316
rect 2010 2123 2013 2206
rect 2018 2143 2021 2313
rect 2034 2236 2037 2506
rect 2050 2496 2053 2736
rect 2046 2493 2053 2496
rect 2046 2416 2049 2493
rect 2058 2423 2061 2706
rect 2066 2516 2069 2846
rect 2082 2823 2085 2903
rect 2090 2806 2093 3136
rect 2098 3133 2101 3153
rect 2114 3136 2117 3263
rect 2110 3133 2117 3136
rect 2098 3013 2101 3046
rect 2110 3026 2113 3133
rect 2110 3023 2117 3026
rect 2098 2976 2101 3006
rect 2106 2976 2109 3006
rect 2098 2973 2109 2976
rect 2098 2943 2101 2973
rect 2114 2966 2117 3023
rect 2122 2983 2125 3273
rect 2130 3106 2133 3296
rect 2146 3266 2149 3353
rect 2138 3263 2149 3266
rect 2138 3226 2141 3263
rect 2138 3223 2149 3226
rect 2146 3146 2149 3223
rect 2170 3203 2173 3326
rect 2178 3303 2181 3336
rect 2194 3276 2197 3346
rect 2258 3333 2261 3356
rect 2202 3323 2221 3326
rect 2274 3313 2277 3336
rect 2194 3273 2213 3276
rect 2178 3203 2189 3206
rect 2138 3143 2149 3146
rect 2138 3123 2141 3143
rect 2186 3133 2189 3196
rect 2130 3103 2141 3106
rect 2106 2963 2117 2966
rect 2098 2813 2101 2886
rect 2086 2803 2093 2806
rect 2074 2713 2077 2736
rect 2086 2716 2089 2803
rect 2106 2786 2109 2963
rect 2138 2956 2141 3103
rect 2162 3086 2165 3116
rect 2154 3083 2165 3086
rect 2130 2953 2141 2956
rect 2114 2903 2117 2936
rect 2122 2933 2125 2946
rect 2130 2916 2133 2953
rect 2126 2913 2133 2916
rect 2114 2803 2117 2846
rect 2106 2783 2113 2786
rect 2098 2723 2101 2766
rect 2110 2716 2113 2783
rect 2126 2776 2129 2913
rect 2138 2813 2141 2926
rect 2146 2873 2149 2936
rect 2146 2793 2149 2806
rect 2126 2773 2133 2776
rect 2086 2713 2093 2716
rect 2090 2633 2093 2713
rect 2106 2713 2113 2716
rect 2122 2713 2125 2756
rect 2074 2583 2077 2626
rect 2098 2623 2101 2636
rect 2106 2606 2109 2713
rect 2130 2636 2133 2773
rect 2154 2766 2157 3016
rect 2170 2973 2173 3086
rect 2186 3016 2189 3056
rect 2194 3026 2197 3266
rect 2210 3166 2213 3273
rect 2202 3163 2213 3166
rect 2202 3143 2205 3163
rect 2234 3063 2237 3126
rect 2194 3023 2213 3026
rect 2186 3013 2197 3016
rect 2162 2903 2165 2916
rect 2170 2896 2173 2926
rect 2178 2903 2181 2986
rect 2186 2933 2189 2976
rect 2162 2893 2173 2896
rect 2162 2803 2165 2893
rect 2186 2823 2189 2916
rect 2138 2763 2157 2766
rect 2138 2703 2141 2763
rect 2154 2743 2173 2746
rect 2146 2706 2149 2736
rect 2154 2723 2157 2743
rect 2162 2726 2165 2736
rect 2170 2733 2173 2743
rect 2178 2726 2181 2766
rect 2162 2723 2181 2726
rect 2146 2703 2157 2706
rect 2102 2603 2109 2606
rect 2114 2633 2133 2636
rect 2102 2536 2105 2603
rect 2082 2533 2093 2536
rect 2102 2533 2109 2536
rect 2090 2516 2093 2533
rect 2066 2513 2077 2516
rect 2074 2436 2077 2513
rect 2066 2433 2077 2436
rect 2086 2513 2093 2516
rect 2086 2436 2089 2513
rect 2098 2463 2101 2516
rect 2086 2433 2093 2436
rect 2046 2413 2053 2416
rect 2050 2333 2053 2413
rect 2026 2233 2037 2236
rect 2026 2193 2029 2233
rect 2034 2213 2045 2216
rect 2050 2203 2053 2326
rect 2058 2313 2061 2336
rect 2026 2163 2037 2166
rect 2034 2133 2037 2163
rect 2066 2156 2069 2433
rect 2074 2403 2077 2416
rect 2090 2413 2093 2433
rect 2098 2383 2101 2406
rect 2074 2323 2093 2326
rect 2098 2323 2101 2336
rect 2090 2303 2093 2316
rect 2106 2306 2109 2533
rect 2114 2503 2117 2633
rect 2154 2626 2157 2703
rect 2122 2623 2133 2626
rect 2154 2623 2165 2626
rect 2122 2613 2157 2616
rect 2146 2563 2149 2606
rect 2102 2303 2109 2306
rect 2066 2153 2077 2156
rect 2042 2106 2045 2126
rect 2034 2103 2045 2106
rect 2010 2023 2013 2046
rect 2034 2036 2037 2103
rect 2034 2033 2045 2036
rect 2010 1823 2013 1906
rect 2010 1713 2013 1726
rect 1998 1703 2005 1706
rect 1998 1636 2001 1703
rect 2018 1696 2021 1946
rect 2026 1896 2029 2016
rect 2042 1933 2045 2033
rect 2050 2013 2053 2036
rect 2058 2023 2061 2146
rect 2074 2046 2077 2153
rect 2090 2123 2093 2246
rect 2102 2176 2105 2303
rect 2114 2183 2117 2426
rect 2122 2413 2125 2526
rect 2130 2486 2133 2536
rect 2138 2503 2141 2526
rect 2154 2523 2157 2613
rect 2162 2523 2165 2623
rect 2178 2583 2181 2706
rect 2186 2603 2189 2796
rect 2194 2583 2197 3013
rect 2202 2816 2205 3016
rect 2210 2906 2213 3023
rect 2218 3003 2221 3026
rect 2218 2926 2221 2946
rect 2226 2933 2237 2936
rect 2218 2923 2229 2926
rect 2210 2903 2221 2906
rect 2202 2813 2209 2816
rect 2206 2746 2209 2813
rect 2202 2743 2209 2746
rect 2202 2566 2205 2743
rect 2170 2523 2173 2546
rect 2130 2483 2149 2486
rect 2102 2173 2109 2176
rect 2106 2106 2109 2173
rect 2122 2166 2125 2406
rect 2146 2356 2149 2483
rect 2170 2403 2173 2426
rect 2130 2353 2149 2356
rect 2130 2316 2133 2353
rect 2138 2333 2149 2336
rect 2130 2313 2137 2316
rect 2134 2186 2137 2313
rect 2146 2213 2149 2333
rect 2154 2323 2157 2336
rect 2186 2333 2189 2566
rect 2198 2563 2205 2566
rect 2198 2496 2201 2563
rect 2210 2533 2213 2716
rect 2218 2706 2221 2903
rect 2234 2796 2237 2816
rect 2230 2793 2237 2796
rect 2230 2726 2233 2793
rect 2242 2733 2245 3306
rect 2306 3276 2309 3326
rect 2298 3273 2309 3276
rect 2298 3226 2301 3273
rect 2314 3246 2317 3266
rect 2314 3243 2325 3246
rect 2298 3223 2309 3226
rect 2258 3213 2277 3216
rect 2250 3023 2253 3126
rect 2298 3123 2301 3206
rect 2306 3133 2309 3223
rect 2322 3196 2325 3243
rect 2338 3226 2341 3366
rect 2346 3303 2349 3326
rect 2354 3283 2357 3393
rect 2474 3356 2477 3406
rect 2314 3193 2325 3196
rect 2334 3223 2341 3226
rect 2314 3123 2317 3193
rect 2322 3133 2325 3176
rect 2334 3146 2337 3223
rect 2334 3143 2341 3146
rect 2346 3143 2349 3216
rect 2370 3203 2373 3306
rect 2418 3303 2421 3336
rect 2434 3333 2437 3356
rect 2466 3353 2477 3356
rect 2442 3333 2445 3346
rect 2426 3313 2437 3316
rect 2258 3083 2261 3116
rect 2330 3106 2333 3126
rect 2322 3103 2333 3106
rect 2282 3003 2285 3026
rect 2298 3013 2301 3086
rect 2322 3026 2325 3103
rect 2306 3023 2325 3026
rect 2306 2963 2309 3023
rect 2314 3003 2317 3016
rect 2322 3003 2325 3016
rect 2330 2976 2333 3016
rect 2322 2973 2333 2976
rect 2250 2923 2253 2946
rect 2250 2813 2253 2866
rect 2258 2803 2261 2926
rect 2322 2916 2325 2973
rect 2330 2923 2333 2966
rect 2314 2913 2325 2916
rect 2230 2723 2237 2726
rect 2218 2703 2225 2706
rect 2222 2646 2225 2703
rect 2218 2643 2225 2646
rect 2218 2563 2221 2643
rect 2226 2613 2229 2626
rect 2226 2583 2229 2606
rect 2210 2523 2221 2526
rect 2210 2503 2213 2523
rect 2226 2506 2229 2576
rect 2222 2503 2229 2506
rect 2198 2493 2205 2496
rect 2194 2393 2197 2406
rect 2202 2376 2205 2493
rect 2222 2426 2225 2503
rect 2198 2373 2205 2376
rect 2154 2303 2157 2316
rect 2178 2246 2181 2296
rect 2198 2266 2201 2373
rect 2210 2293 2213 2426
rect 2222 2423 2229 2426
rect 2226 2386 2229 2423
rect 2222 2383 2229 2386
rect 2198 2263 2205 2266
rect 2174 2243 2181 2246
rect 2154 2203 2157 2236
rect 2118 2163 2125 2166
rect 2130 2183 2137 2186
rect 2162 2183 2165 2216
rect 2130 2163 2133 2183
rect 2118 2106 2121 2163
rect 2174 2156 2177 2243
rect 2174 2153 2181 2156
rect 2130 2143 2149 2146
rect 2130 2133 2133 2143
rect 2146 2136 2149 2143
rect 2066 2043 2077 2046
rect 2098 2103 2109 2106
rect 2114 2103 2121 2106
rect 2050 1933 2053 1956
rect 2066 1946 2069 2043
rect 2098 2026 2101 2103
rect 2058 1943 2069 1946
rect 2042 1923 2053 1926
rect 2026 1893 2053 1896
rect 2026 1823 2029 1856
rect 2026 1783 2029 1816
rect 2034 1803 2037 1886
rect 2026 1713 2029 1736
rect 1950 1593 1957 1596
rect 1950 1446 1953 1593
rect 1962 1453 1965 1616
rect 1974 1613 1981 1616
rect 1974 1536 1977 1613
rect 1974 1533 1981 1536
rect 1970 1493 1973 1516
rect 1950 1443 1957 1446
rect 1946 1403 1949 1426
rect 1890 1283 1901 1286
rect 1882 1223 1885 1246
rect 1874 1213 1885 1216
rect 1890 1213 1893 1283
rect 1834 1173 1845 1176
rect 1818 1163 1829 1166
rect 1818 1133 1821 1146
rect 1810 1123 1821 1126
rect 1826 1086 1829 1163
rect 1834 1093 1837 1173
rect 1858 1156 1861 1206
rect 1858 1153 1877 1156
rect 1842 1133 1869 1136
rect 1794 1016 1797 1086
rect 1790 1013 1797 1016
rect 1810 1083 1829 1086
rect 1762 976 1765 1006
rect 1770 986 1773 996
rect 1770 983 1781 986
rect 1762 973 1773 976
rect 1746 913 1749 926
rect 1754 913 1757 936
rect 1762 933 1765 956
rect 1770 936 1773 973
rect 1778 963 1781 983
rect 1790 956 1793 1013
rect 1802 973 1805 1006
rect 1810 996 1813 1083
rect 1818 1016 1821 1076
rect 1826 1023 1829 1083
rect 1818 1013 1829 1016
rect 1834 1013 1837 1026
rect 1826 1003 1829 1013
rect 1810 993 1829 996
rect 1834 993 1837 1006
rect 1790 953 1797 956
rect 1770 933 1781 936
rect 1770 916 1773 926
rect 1786 923 1789 936
rect 1770 913 1789 916
rect 1738 903 1781 906
rect 1690 803 1693 836
rect 1706 823 1717 826
rect 1738 823 1741 846
rect 1682 793 1693 796
rect 1666 763 1673 766
rect 1666 743 1669 763
rect 1650 713 1661 716
rect 1658 646 1661 713
rect 1674 653 1677 736
rect 1682 723 1685 756
rect 1658 643 1669 646
rect 1618 623 1653 626
rect 1618 613 1629 616
rect 1578 603 1597 606
rect 1562 533 1589 536
rect 1546 523 1557 526
rect 1526 503 1533 506
rect 1538 513 1549 516
rect 1526 436 1529 503
rect 1514 433 1529 436
rect 1498 396 1501 406
rect 1466 393 1501 396
rect 1426 383 1437 386
rect 1418 316 1421 366
rect 1410 313 1421 316
rect 1314 223 1317 266
rect 1410 236 1413 313
rect 1434 266 1437 383
rect 1514 373 1517 433
rect 1522 396 1525 416
rect 1530 403 1533 426
rect 1538 413 1541 513
rect 1554 413 1557 523
rect 1562 413 1565 526
rect 1578 473 1581 526
rect 1522 393 1533 396
rect 1466 333 1469 356
rect 1458 323 1477 326
rect 1490 323 1493 336
rect 1498 333 1517 336
rect 1514 326 1517 333
rect 1514 323 1525 326
rect 1530 323 1533 393
rect 1562 376 1565 406
rect 1554 373 1573 376
rect 1570 356 1573 373
rect 1578 363 1581 406
rect 1594 383 1597 603
rect 1610 603 1629 606
rect 1610 573 1613 603
rect 1618 523 1621 556
rect 1634 533 1637 586
rect 1626 513 1629 526
rect 1642 523 1645 576
rect 1650 533 1653 566
rect 1658 503 1661 616
rect 1666 443 1669 643
rect 1674 603 1677 616
rect 1682 593 1685 606
rect 1690 513 1693 793
rect 1698 773 1701 806
rect 1706 746 1709 823
rect 1714 793 1717 816
rect 1746 813 1749 826
rect 1722 803 1741 806
rect 1698 743 1709 746
rect 1698 723 1701 743
rect 1698 583 1701 626
rect 1706 533 1709 736
rect 1714 703 1717 786
rect 1722 723 1725 776
rect 1746 733 1749 756
rect 1722 713 1741 716
rect 1714 616 1717 656
rect 1722 623 1725 713
rect 1730 693 1733 706
rect 1714 613 1725 616
rect 1722 546 1725 613
rect 1730 566 1733 636
rect 1746 623 1749 636
rect 1746 593 1749 606
rect 1730 563 1741 566
rect 1714 543 1725 546
rect 1618 413 1621 426
rect 1642 413 1653 416
rect 1618 393 1621 406
rect 1666 396 1669 406
rect 1674 403 1677 456
rect 1682 413 1685 426
rect 1714 423 1717 543
rect 1722 523 1725 536
rect 1738 533 1741 563
rect 1754 546 1757 896
rect 1762 823 1765 836
rect 1762 793 1765 806
rect 1762 653 1765 736
rect 1762 613 1765 626
rect 1754 543 1765 546
rect 1730 523 1741 526
rect 1754 516 1757 536
rect 1698 413 1717 416
rect 1682 403 1693 406
rect 1682 396 1685 403
rect 1666 393 1685 396
rect 1570 353 1581 356
rect 1602 346 1605 366
rect 1474 316 1477 323
rect 1474 313 1517 316
rect 1498 303 1509 306
rect 1426 263 1437 266
rect 1426 243 1429 263
rect 1370 223 1373 236
rect 1410 233 1437 236
rect 1378 213 1381 226
rect 1266 133 1277 136
rect 1258 113 1261 126
rect 1266 106 1269 126
rect 1234 103 1269 106
rect 1234 96 1237 103
rect 1218 93 1237 96
rect 1090 83 1133 86
rect 682 0 685 26
rect 1034 23 1037 83
rect 1106 0 1109 76
rect 1274 73 1277 133
rect 1290 123 1293 136
rect 1298 113 1301 206
rect 1338 186 1341 206
rect 1330 183 1341 186
rect 1306 113 1309 136
rect 1330 126 1333 183
rect 1354 173 1357 206
rect 1386 203 1389 216
rect 1394 193 1397 206
rect 1410 203 1413 233
rect 1418 156 1421 216
rect 1426 203 1429 226
rect 1434 203 1437 233
rect 1522 226 1525 323
rect 1442 203 1445 216
rect 1458 193 1461 216
rect 1466 203 1469 226
rect 1522 223 1541 226
rect 1514 203 1517 216
rect 1522 203 1525 223
rect 1530 156 1533 216
rect 1538 196 1541 223
rect 1546 203 1549 216
rect 1554 203 1557 226
rect 1578 216 1581 346
rect 1602 343 1613 346
rect 1610 296 1613 343
rect 1602 293 1613 296
rect 1626 293 1629 326
rect 1578 213 1589 216
rect 1538 193 1549 196
rect 1346 133 1349 156
rect 1418 153 1429 156
rect 1330 123 1349 126
rect 1346 96 1349 123
rect 1354 106 1357 126
rect 1354 103 1365 106
rect 1370 96 1373 116
rect 1346 93 1373 96
rect 1378 93 1381 126
rect 1386 113 1389 136
rect 1418 133 1421 146
rect 1426 126 1429 153
rect 1490 153 1533 156
rect 1466 126 1469 136
rect 1490 126 1493 153
rect 1370 86 1373 93
rect 1394 86 1397 126
rect 1418 123 1429 126
rect 1410 103 1413 116
rect 1418 113 1421 123
rect 1370 83 1397 86
rect 1434 83 1437 126
rect 1466 123 1493 126
rect 1498 116 1501 136
rect 1514 133 1517 146
rect 1514 116 1517 126
rect 1490 93 1493 116
rect 1498 113 1517 116
rect 1538 113 1541 176
rect 1570 93 1573 136
rect 1586 133 1589 213
rect 1602 203 1605 293
rect 1610 213 1621 216
rect 1634 206 1637 256
rect 1642 213 1645 236
rect 1634 203 1645 206
rect 1650 173 1653 216
rect 1634 123 1637 136
rect 1666 123 1669 326
rect 1674 323 1677 386
rect 1714 363 1717 406
rect 1722 403 1725 426
rect 1738 423 1741 516
rect 1750 513 1757 516
rect 1690 236 1693 346
rect 1730 303 1733 416
rect 1750 406 1753 513
rect 1750 403 1757 406
rect 1754 383 1757 403
rect 1762 376 1765 543
rect 1770 393 1773 896
rect 1778 706 1781 903
rect 1786 713 1789 913
rect 1794 756 1797 953
rect 1802 893 1805 936
rect 1810 933 1813 986
rect 1802 773 1805 816
rect 1810 813 1813 906
rect 1818 873 1821 926
rect 1826 903 1829 993
rect 1834 863 1837 896
rect 1826 823 1829 846
rect 1834 813 1837 836
rect 1818 803 1829 806
rect 1834 793 1837 806
rect 1794 753 1801 756
rect 1778 703 1785 706
rect 1782 636 1785 703
rect 1798 696 1801 753
rect 1834 743 1837 766
rect 1826 733 1837 736
rect 1794 693 1801 696
rect 1782 633 1789 636
rect 1778 596 1781 616
rect 1786 613 1789 633
rect 1778 593 1785 596
rect 1782 496 1785 593
rect 1794 543 1797 693
rect 1810 653 1813 726
rect 1834 683 1837 726
rect 1842 703 1845 1133
rect 1850 1023 1853 1116
rect 1866 1016 1869 1126
rect 1874 1123 1877 1153
rect 1882 1106 1885 1213
rect 1854 1013 1869 1016
rect 1878 1103 1885 1106
rect 1854 956 1857 1013
rect 1850 953 1857 956
rect 1850 923 1853 953
rect 1850 873 1853 916
rect 1858 853 1861 936
rect 1866 933 1869 956
rect 1866 826 1869 926
rect 1878 916 1881 1103
rect 1890 973 1893 1186
rect 1898 1163 1901 1206
rect 1898 1083 1901 1136
rect 1898 1013 1901 1026
rect 1850 823 1869 826
rect 1874 913 1881 916
rect 1890 913 1893 946
rect 1906 933 1909 1306
rect 1914 1213 1917 1313
rect 1922 1303 1941 1306
rect 1946 1246 1949 1326
rect 1922 1243 1949 1246
rect 1922 1213 1925 1243
rect 1954 1236 1957 1443
rect 1962 1393 1965 1416
rect 1962 1303 1965 1366
rect 1922 1136 1925 1206
rect 1914 1133 1925 1136
rect 1914 1123 1917 1133
rect 1930 1126 1933 1236
rect 1938 1233 1957 1236
rect 1938 1176 1941 1233
rect 1962 1216 1965 1286
rect 1970 1233 1973 1426
rect 1978 1316 1981 1533
rect 1986 1453 1989 1636
rect 1998 1633 2005 1636
rect 1986 1413 1989 1446
rect 1986 1333 1989 1366
rect 1978 1313 1989 1316
rect 1978 1283 1981 1306
rect 1954 1213 1965 1216
rect 1946 1186 1949 1206
rect 1970 1193 1973 1216
rect 1946 1183 1965 1186
rect 1938 1173 1949 1176
rect 1946 1133 1949 1173
rect 1954 1133 1957 1176
rect 1922 1106 1925 1126
rect 1930 1123 1957 1126
rect 1922 1103 1933 1106
rect 1914 1003 1917 1096
rect 1930 1026 1933 1103
rect 1922 1023 1933 1026
rect 1922 933 1925 1023
rect 1930 933 1933 956
rect 1850 733 1853 823
rect 1858 803 1861 816
rect 1858 793 1869 796
rect 1866 733 1869 793
rect 1802 603 1805 626
rect 1810 613 1821 616
rect 1826 613 1829 666
rect 1810 586 1813 613
rect 1818 593 1821 606
rect 1834 603 1837 676
rect 1850 636 1853 726
rect 1866 683 1869 716
rect 1842 633 1853 636
rect 1842 613 1845 633
rect 1850 613 1853 626
rect 1842 603 1853 606
rect 1858 603 1861 646
rect 1866 613 1869 656
rect 1810 583 1821 586
rect 1850 583 1853 603
rect 1810 533 1813 546
rect 1810 513 1813 526
rect 1778 493 1785 496
rect 1754 373 1765 376
rect 1754 346 1757 373
rect 1762 353 1773 356
rect 1754 343 1765 346
rect 1738 323 1741 336
rect 1762 276 1765 343
rect 1770 323 1773 353
rect 1778 283 1781 493
rect 1786 436 1789 476
rect 1818 473 1821 583
rect 1850 523 1853 576
rect 1866 526 1869 536
rect 1858 523 1869 526
rect 1826 513 1837 516
rect 1858 493 1861 523
rect 1786 433 1813 436
rect 1786 423 1789 433
rect 1794 416 1797 426
rect 1794 413 1805 416
rect 1810 413 1813 433
rect 1826 413 1829 466
rect 1874 456 1877 913
rect 1914 906 1917 926
rect 1882 813 1885 906
rect 1906 903 1917 906
rect 1906 836 1909 903
rect 1906 833 1917 836
rect 1882 723 1885 786
rect 1890 733 1893 806
rect 1898 716 1901 816
rect 1914 813 1917 833
rect 1906 766 1909 806
rect 1922 803 1925 926
rect 1930 803 1933 906
rect 1938 803 1941 1006
rect 1946 793 1949 1086
rect 1954 863 1957 1123
rect 1906 763 1917 766
rect 1890 713 1901 716
rect 1890 693 1893 713
rect 1882 613 1885 626
rect 1890 583 1893 606
rect 1898 603 1901 706
rect 1906 626 1909 736
rect 1914 723 1917 763
rect 1922 653 1925 766
rect 1954 746 1957 826
rect 1962 806 1965 1183
rect 1970 1123 1973 1136
rect 1978 1083 1981 1226
rect 1986 1026 1989 1313
rect 1970 1023 1989 1026
rect 1970 986 1973 1016
rect 1978 993 1981 1006
rect 1970 983 1981 986
rect 1970 833 1973 936
rect 1978 906 1981 983
rect 1986 923 1989 1023
rect 1994 933 1997 1616
rect 2002 1423 2005 1633
rect 2010 1623 2013 1696
rect 2018 1693 2025 1696
rect 2022 1626 2025 1693
rect 2018 1623 2025 1626
rect 2010 1586 2013 1616
rect 2018 1593 2021 1623
rect 2026 1593 2029 1606
rect 2010 1583 2029 1586
rect 2034 1583 2037 1736
rect 2010 1523 2013 1556
rect 2018 1533 2021 1546
rect 2026 1526 2029 1583
rect 2018 1523 2029 1526
rect 2018 1403 2021 1523
rect 2034 1473 2037 1556
rect 2026 1423 2037 1426
rect 2002 1343 2021 1346
rect 2002 1323 2005 1343
rect 2010 1323 2013 1336
rect 2018 1333 2021 1343
rect 2042 1336 2045 1856
rect 2050 1836 2053 1893
rect 2058 1853 2061 1943
rect 2050 1833 2057 1836
rect 2054 1746 2057 1833
rect 2050 1743 2057 1746
rect 2050 1593 2053 1743
rect 2058 1683 2061 1726
rect 2066 1706 2069 1936
rect 2074 1813 2077 1956
rect 2082 1873 2085 2026
rect 2098 2023 2105 2026
rect 2090 1883 2093 2006
rect 2102 1956 2105 2023
rect 2102 1953 2109 1956
rect 2098 1923 2101 1936
rect 2106 1906 2109 1953
rect 2114 1943 2117 2103
rect 2138 2096 2141 2136
rect 2146 2133 2157 2136
rect 2154 2123 2165 2126
rect 2122 2093 2141 2096
rect 2102 1903 2109 1906
rect 2102 1826 2105 1903
rect 2102 1823 2109 1826
rect 2082 1733 2085 1766
rect 2074 1723 2085 1726
rect 2066 1703 2073 1706
rect 2058 1586 2061 1646
rect 2050 1583 2061 1586
rect 2050 1413 2053 1583
rect 2058 1473 2061 1576
rect 2070 1566 2073 1703
rect 2082 1613 2085 1636
rect 2082 1593 2085 1606
rect 2066 1563 2073 1566
rect 2026 1326 2029 1336
rect 2042 1333 2049 1336
rect 2018 1323 2029 1326
rect 2018 1316 2021 1323
rect 2002 1313 2021 1316
rect 2002 1123 2005 1313
rect 2010 1233 2013 1306
rect 2034 1276 2037 1326
rect 2026 1273 2037 1276
rect 2026 1213 2029 1273
rect 2010 1193 2013 1206
rect 2010 1133 2013 1156
rect 2010 1093 2013 1116
rect 2018 1096 2021 1136
rect 2026 1123 2029 1206
rect 2034 1106 2037 1236
rect 2046 1226 2049 1333
rect 2042 1223 2049 1226
rect 2042 1113 2045 1223
rect 2050 1163 2053 1206
rect 2034 1103 2045 1106
rect 2018 1093 2037 1096
rect 2002 1023 2005 1076
rect 2018 1046 2021 1086
rect 2010 1043 2021 1046
rect 2002 963 2005 1006
rect 2010 993 2013 1043
rect 2034 1036 2037 1093
rect 2018 1033 2037 1036
rect 2018 993 2021 1033
rect 1978 903 1985 906
rect 2002 903 2005 946
rect 1962 803 1973 806
rect 1946 743 1957 746
rect 1930 626 1933 726
rect 1938 663 1941 736
rect 1946 673 1949 743
rect 1954 643 1957 736
rect 1906 623 1917 626
rect 1906 603 1909 616
rect 1914 566 1917 623
rect 1898 563 1917 566
rect 1922 623 1933 626
rect 1922 563 1925 623
rect 1890 503 1893 536
rect 1898 486 1901 563
rect 1922 536 1925 556
rect 1930 546 1933 616
rect 1946 613 1957 616
rect 1962 613 1965 796
rect 1970 636 1973 803
rect 1982 756 1985 903
rect 1994 823 1997 836
rect 1978 753 1985 756
rect 1978 733 1981 753
rect 1970 633 1981 636
rect 1930 543 1949 546
rect 1866 453 1877 456
rect 1894 483 1901 486
rect 1786 383 1789 406
rect 1794 393 1797 406
rect 1802 343 1805 413
rect 1810 366 1813 406
rect 1810 363 1821 366
rect 1826 363 1829 406
rect 1866 376 1869 453
rect 1866 373 1877 376
rect 1818 353 1821 363
rect 1874 353 1877 373
rect 1802 323 1805 336
rect 1850 303 1853 326
rect 1882 323 1885 446
rect 1894 416 1897 483
rect 1894 413 1901 416
rect 1898 396 1901 413
rect 1906 406 1909 536
rect 1922 533 1933 536
rect 1914 513 1917 526
rect 1922 523 1933 526
rect 1930 503 1933 516
rect 1938 483 1941 536
rect 1922 413 1925 426
rect 1930 413 1933 476
rect 1946 463 1949 543
rect 1954 536 1957 606
rect 1970 583 1973 626
rect 1978 576 1981 633
rect 1986 613 1989 646
rect 1994 633 1997 806
rect 2002 803 2005 846
rect 2018 806 2021 946
rect 2026 933 2029 1006
rect 2034 933 2037 1016
rect 2042 1003 2045 1103
rect 2050 936 2053 1136
rect 2058 1083 2061 1406
rect 2066 1316 2069 1563
rect 2090 1556 2093 1806
rect 2098 1723 2101 1806
rect 2098 1603 2101 1686
rect 2090 1553 2101 1556
rect 2074 1543 2101 1546
rect 2074 1413 2077 1456
rect 2074 1383 2077 1406
rect 2074 1333 2077 1366
rect 2066 1313 2073 1316
rect 2070 1246 2073 1313
rect 2082 1283 2085 1536
rect 2098 1523 2101 1543
rect 2090 1383 2093 1506
rect 2098 1393 2101 1516
rect 2098 1323 2101 1336
rect 2098 1303 2101 1316
rect 2106 1296 2109 1823
rect 2114 1803 2117 1936
rect 2122 1803 2125 2093
rect 2130 1933 2133 2086
rect 2114 1713 2117 1766
rect 2122 1693 2125 1726
rect 2130 1646 2133 1876
rect 2138 1866 2141 2046
rect 2154 2013 2157 2106
rect 2170 2006 2173 2076
rect 2154 2003 2173 2006
rect 2178 1986 2181 2153
rect 2186 2043 2189 2236
rect 2194 2113 2197 2246
rect 2186 2013 2189 2026
rect 2146 1923 2149 1986
rect 2174 1983 2181 1986
rect 2154 1933 2157 1966
rect 2162 1866 2165 1936
rect 2174 1926 2177 1983
rect 2174 1923 2181 1926
rect 2178 1903 2181 1923
rect 2138 1863 2157 1866
rect 2162 1863 2181 1866
rect 2138 1823 2141 1856
rect 2138 1706 2141 1816
rect 2146 1723 2149 1816
rect 2154 1796 2157 1863
rect 2170 1816 2173 1856
rect 2162 1813 2173 1816
rect 2178 1806 2181 1863
rect 2186 1853 2189 2006
rect 2194 1813 2197 2066
rect 2202 1953 2205 2263
rect 2170 1803 2181 1806
rect 2202 1803 2205 1936
rect 2154 1793 2161 1796
rect 2158 1736 2161 1793
rect 2158 1733 2165 1736
rect 2138 1703 2145 1706
rect 2114 1643 2133 1646
rect 2114 1513 2117 1643
rect 2122 1613 2125 1636
rect 2142 1626 2145 1703
rect 2154 1693 2157 1726
rect 2142 1623 2149 1626
rect 2122 1603 2133 1606
rect 2122 1533 2125 1596
rect 2114 1393 2117 1506
rect 2130 1476 2133 1576
rect 2138 1553 2141 1616
rect 2146 1543 2149 1623
rect 2154 1516 2157 1606
rect 2162 1596 2165 1733
rect 2170 1706 2173 1803
rect 2170 1703 2177 1706
rect 2174 1636 2177 1703
rect 2186 1663 2189 1766
rect 2194 1733 2197 1746
rect 2170 1633 2177 1636
rect 2170 1613 2173 1633
rect 2162 1593 2169 1596
rect 2138 1513 2157 1516
rect 2138 1483 2141 1513
rect 2166 1496 2169 1593
rect 2130 1473 2141 1476
rect 2114 1356 2117 1386
rect 2122 1363 2125 1416
rect 2130 1403 2133 1416
rect 2138 1363 2141 1473
rect 2154 1443 2157 1496
rect 2162 1493 2169 1496
rect 2154 1393 2157 1416
rect 2114 1353 2125 1356
rect 2122 1323 2125 1353
rect 2090 1293 2109 1296
rect 2066 1243 2073 1246
rect 2066 1123 2069 1243
rect 2074 1163 2077 1226
rect 2082 1173 2085 1216
rect 2090 1196 2093 1293
rect 2098 1203 2101 1286
rect 2106 1276 2109 1293
rect 2130 1283 2133 1336
rect 2138 1333 2141 1346
rect 2154 1343 2157 1386
rect 2106 1273 2133 1276
rect 2106 1203 2109 1216
rect 2090 1193 2109 1196
rect 2074 1133 2077 1146
rect 2090 1123 2093 1146
rect 2098 1143 2101 1176
rect 2098 1056 2101 1136
rect 2106 1106 2109 1193
rect 2114 1183 2117 1206
rect 2114 1123 2117 1156
rect 2122 1146 2125 1216
rect 2130 1213 2133 1273
rect 2130 1153 2133 1206
rect 2122 1143 2133 1146
rect 2106 1103 2113 1106
rect 2122 1103 2125 1136
rect 2066 1053 2101 1056
rect 2058 1013 2061 1046
rect 2066 946 2069 1053
rect 2082 1013 2093 1016
rect 2098 1013 2101 1046
rect 2110 1036 2113 1103
rect 2106 1033 2113 1036
rect 2074 993 2077 1006
rect 2090 973 2093 1006
rect 2098 946 2101 1006
rect 2106 976 2109 1033
rect 2114 993 2117 1016
rect 2106 973 2117 976
rect 2130 973 2133 1143
rect 2042 933 2053 936
rect 2058 943 2101 946
rect 2042 906 2045 933
rect 2050 916 2053 926
rect 2058 923 2061 943
rect 2066 916 2069 936
rect 2050 913 2069 916
rect 2074 906 2077 926
rect 2082 923 2085 936
rect 2090 913 2093 926
rect 2042 903 2093 906
rect 2098 903 2101 936
rect 2090 896 2093 903
rect 2090 893 2101 896
rect 2042 823 2045 866
rect 2026 813 2045 816
rect 2066 813 2069 856
rect 2018 803 2045 806
rect 2050 793 2061 796
rect 2002 733 2005 766
rect 1970 573 1981 576
rect 1954 533 1965 536
rect 1954 503 1957 526
rect 1970 523 1973 573
rect 1978 523 1981 546
rect 1938 423 1949 426
rect 1954 416 1957 476
rect 1994 443 1997 606
rect 2002 573 2005 626
rect 2010 613 2013 756
rect 2018 743 2029 746
rect 2018 733 2037 736
rect 2018 696 2021 733
rect 2026 716 2029 726
rect 2034 723 2037 733
rect 2066 723 2069 736
rect 2074 716 2077 816
rect 2082 763 2085 856
rect 2098 823 2101 893
rect 2114 846 2117 973
rect 2138 953 2141 1326
rect 2146 1316 2149 1336
rect 2146 1313 2153 1316
rect 2150 1246 2153 1313
rect 2146 1243 2153 1246
rect 2146 1026 2149 1243
rect 2154 1203 2157 1226
rect 2154 1123 2157 1186
rect 2162 1176 2165 1493
rect 2178 1483 2181 1616
rect 2186 1523 2189 1616
rect 2194 1593 2197 1616
rect 2202 1603 2205 1776
rect 2210 1743 2213 2286
rect 2222 2256 2225 2383
rect 2234 2346 2237 2723
rect 2250 2706 2253 2726
rect 2258 2723 2261 2736
rect 2242 2593 2245 2706
rect 2250 2703 2257 2706
rect 2254 2586 2257 2703
rect 2250 2583 2257 2586
rect 2250 2536 2253 2583
rect 2250 2533 2257 2536
rect 2242 2393 2245 2526
rect 2254 2436 2257 2533
rect 2250 2433 2257 2436
rect 2250 2353 2253 2433
rect 2258 2383 2261 2416
rect 2234 2343 2245 2346
rect 2222 2253 2229 2256
rect 2226 2233 2229 2253
rect 2218 2203 2221 2216
rect 2226 2193 2229 2206
rect 2234 2196 2237 2336
rect 2242 2326 2245 2343
rect 2242 2323 2253 2326
rect 2250 2246 2253 2323
rect 2266 2306 2269 2906
rect 2274 2813 2277 2826
rect 2274 2613 2277 2726
rect 2282 2713 2285 2736
rect 2290 2683 2293 2816
rect 2290 2633 2293 2666
rect 2298 2626 2301 2796
rect 2314 2756 2317 2913
rect 2338 2896 2341 3143
rect 2362 3116 2365 3136
rect 2358 3113 2365 3116
rect 2346 2923 2349 3066
rect 2358 3026 2361 3113
rect 2358 3023 2365 3026
rect 2330 2893 2341 2896
rect 2330 2836 2333 2893
rect 2330 2833 2341 2836
rect 2314 2753 2321 2756
rect 2290 2623 2301 2626
rect 2274 2393 2277 2526
rect 2282 2323 2285 2576
rect 2290 2553 2293 2623
rect 2306 2616 2309 2736
rect 2298 2613 2309 2616
rect 2298 2546 2301 2613
rect 2306 2553 2309 2606
rect 2290 2543 2301 2546
rect 2318 2546 2321 2753
rect 2330 2546 2333 2816
rect 2338 2746 2341 2833
rect 2346 2813 2349 2886
rect 2354 2833 2357 3006
rect 2362 2953 2365 3023
rect 2370 2933 2373 3186
rect 2378 2993 2381 3296
rect 2386 3203 2389 3216
rect 2394 3203 2397 3286
rect 2402 3156 2405 3216
rect 2410 3183 2413 3216
rect 2386 3153 2405 3156
rect 2386 3123 2389 3153
rect 2394 3143 2405 3146
rect 2394 3076 2397 3136
rect 2402 3133 2405 3143
rect 2410 3123 2413 3156
rect 2394 3073 2405 3076
rect 2386 2913 2389 3066
rect 2402 3026 2405 3073
rect 2418 3056 2421 3246
rect 2426 3133 2429 3146
rect 2394 3023 2405 3026
rect 2414 3053 2421 3056
rect 2394 3003 2397 3023
rect 2414 2996 2417 3053
rect 2426 3003 2429 3046
rect 2434 3013 2437 3166
rect 2442 3123 2445 3296
rect 2466 3206 2469 3353
rect 2482 3293 2485 3326
rect 2466 3203 2477 3206
rect 2490 3203 2493 3346
rect 2538 3333 2541 3386
rect 2554 3333 2565 3336
rect 2538 3313 2541 3326
rect 2546 3323 2565 3326
rect 2570 3316 2573 3336
rect 2602 3323 2605 3366
rect 2658 3333 2677 3336
rect 2658 3316 2661 3326
rect 2498 3213 2517 3216
rect 2474 3186 2477 3203
rect 2458 3136 2461 3186
rect 2474 3183 2485 3186
rect 2454 3133 2461 3136
rect 2442 3003 2445 3116
rect 2454 3036 2457 3133
rect 2454 3033 2461 3036
rect 2414 2993 2421 2996
rect 2370 2806 2373 2846
rect 2362 2803 2373 2806
rect 2362 2746 2365 2803
rect 2338 2743 2349 2746
rect 2362 2743 2373 2746
rect 2338 2723 2341 2736
rect 2346 2633 2349 2743
rect 2370 2723 2373 2743
rect 2338 2613 2341 2626
rect 2354 2616 2357 2666
rect 2378 2653 2381 2866
rect 2386 2823 2389 2836
rect 2394 2806 2397 2956
rect 2390 2803 2397 2806
rect 2390 2646 2393 2803
rect 2402 2733 2405 2846
rect 2410 2823 2413 2906
rect 2418 2816 2421 2993
rect 2450 2963 2453 3016
rect 2450 2923 2453 2936
rect 2426 2833 2429 2906
rect 2434 2833 2445 2836
rect 2410 2813 2421 2816
rect 2426 2813 2437 2816
rect 2390 2643 2397 2646
rect 2346 2573 2349 2616
rect 2354 2613 2365 2616
rect 2318 2543 2325 2546
rect 2330 2543 2341 2546
rect 2354 2543 2357 2606
rect 2290 2343 2293 2543
rect 2298 2373 2301 2536
rect 2306 2523 2309 2536
rect 2306 2413 2309 2486
rect 2314 2463 2317 2526
rect 2322 2503 2325 2543
rect 2330 2486 2333 2526
rect 2326 2483 2333 2486
rect 2326 2406 2329 2483
rect 2338 2413 2341 2536
rect 2346 2433 2349 2506
rect 2298 2333 2301 2356
rect 2242 2243 2253 2246
rect 2262 2303 2269 2306
rect 2242 2206 2245 2243
rect 2250 2213 2253 2226
rect 2242 2203 2253 2206
rect 2234 2193 2245 2196
rect 2218 1953 2221 2136
rect 2226 1946 2229 2146
rect 2242 2123 2245 2193
rect 2250 2116 2253 2203
rect 2262 2196 2265 2303
rect 2290 2296 2293 2316
rect 2274 2203 2277 2296
rect 2286 2293 2293 2296
rect 2286 2196 2289 2293
rect 2298 2263 2301 2326
rect 2298 2203 2301 2246
rect 2262 2193 2269 2196
rect 2286 2193 2293 2196
rect 2234 2113 2253 2116
rect 2234 2013 2237 2113
rect 2242 2003 2245 2046
rect 2250 2013 2253 2026
rect 2226 1943 2253 1946
rect 2226 1933 2237 1936
rect 2210 1613 2213 1666
rect 2218 1556 2221 1926
rect 2242 1923 2245 1936
rect 2250 1906 2253 1943
rect 2242 1903 2253 1906
rect 2226 1836 2229 1856
rect 2226 1833 2233 1836
rect 2230 1626 2233 1833
rect 2242 1826 2245 1903
rect 2242 1823 2253 1826
rect 2258 1823 2261 2146
rect 2226 1623 2233 1626
rect 2226 1606 2229 1623
rect 2226 1603 2237 1606
rect 2194 1476 2197 1556
rect 2214 1553 2221 1556
rect 2242 1556 2245 1806
rect 2250 1743 2253 1823
rect 2250 1683 2253 1726
rect 2258 1693 2261 1736
rect 2266 1676 2269 2193
rect 2274 2103 2277 2146
rect 2290 2126 2293 2193
rect 2290 2123 2297 2126
rect 2282 2023 2285 2116
rect 2294 2046 2297 2123
rect 2290 2043 2297 2046
rect 2274 1736 2277 2016
rect 2282 1763 2285 1926
rect 2290 1756 2293 2043
rect 2298 1803 2301 2026
rect 2306 2013 2309 2406
rect 2314 2333 2317 2406
rect 2326 2403 2333 2406
rect 2314 2303 2317 2326
rect 2330 2226 2333 2403
rect 2354 2363 2357 2516
rect 2362 2403 2365 2556
rect 2362 2316 2365 2336
rect 2354 2313 2365 2316
rect 2354 2236 2357 2313
rect 2354 2233 2365 2236
rect 2322 2223 2333 2226
rect 2314 2163 2317 2216
rect 2314 2043 2317 2116
rect 2306 1866 2309 1956
rect 2314 1933 2317 1966
rect 2322 1933 2325 2223
rect 2330 2123 2333 2216
rect 2338 2163 2341 2206
rect 2338 2113 2341 2126
rect 2346 2086 2349 2216
rect 2354 2173 2357 2206
rect 2362 2146 2365 2233
rect 2370 2193 2373 2636
rect 2378 2586 2381 2616
rect 2386 2603 2389 2626
rect 2378 2583 2389 2586
rect 2378 2533 2381 2583
rect 2378 2463 2381 2506
rect 2378 2413 2381 2456
rect 2386 2403 2389 2546
rect 2394 2506 2397 2643
rect 2402 2573 2405 2726
rect 2410 2666 2413 2813
rect 2450 2806 2453 2906
rect 2418 2803 2453 2806
rect 2418 2686 2421 2803
rect 2426 2783 2437 2786
rect 2426 2723 2429 2783
rect 2450 2776 2453 2796
rect 2458 2783 2461 3033
rect 2466 3013 2469 3126
rect 2482 3106 2485 3183
rect 2514 3176 2517 3206
rect 2522 3203 2525 3266
rect 2506 3173 2517 3176
rect 2506 3123 2509 3173
rect 2514 3133 2517 3166
rect 2482 3103 2493 3106
rect 2490 3036 2493 3103
rect 2474 3033 2493 3036
rect 2474 3003 2477 3033
rect 2522 3023 2525 3046
rect 2530 3016 2533 3126
rect 2538 3036 2541 3226
rect 2562 3223 2565 3316
rect 2570 3313 2581 3316
rect 2642 3313 2661 3316
rect 2578 3296 2581 3313
rect 2578 3293 2589 3296
rect 2586 3236 2589 3293
rect 2570 3233 2589 3236
rect 2570 3203 2573 3233
rect 2586 3213 2597 3216
rect 2626 3213 2629 3226
rect 2586 3186 2589 3213
rect 2578 3183 2589 3186
rect 2546 3073 2549 3136
rect 2554 3113 2557 3136
rect 2578 3116 2581 3183
rect 2594 3123 2597 3206
rect 2634 3203 2637 3296
rect 2578 3113 2597 3116
rect 2562 3046 2565 3106
rect 2586 3086 2589 3106
rect 2582 3083 2589 3086
rect 2562 3043 2573 3046
rect 2538 3033 2557 3036
rect 2538 3023 2549 3026
rect 2466 2886 2469 2916
rect 2474 2903 2477 2966
rect 2482 2943 2485 3016
rect 2522 3013 2533 3016
rect 2490 2993 2517 2996
rect 2466 2883 2477 2886
rect 2474 2816 2477 2883
rect 2470 2813 2477 2816
rect 2434 2773 2453 2776
rect 2434 2733 2437 2773
rect 2450 2733 2453 2773
rect 2442 2696 2445 2726
rect 2458 2696 2461 2756
rect 2470 2736 2473 2813
rect 2490 2796 2493 2993
rect 2498 2946 2501 2986
rect 2514 2983 2517 2993
rect 2522 2963 2525 3013
rect 2530 2976 2533 3006
rect 2530 2973 2549 2976
rect 2498 2943 2509 2946
rect 2506 2846 2509 2943
rect 2538 2933 2541 2966
rect 2530 2913 2533 2926
rect 2546 2906 2549 2973
rect 2554 2926 2557 3033
rect 2570 2956 2573 3043
rect 2562 2953 2573 2956
rect 2562 2933 2565 2953
rect 2554 2923 2565 2926
rect 2562 2913 2565 2923
rect 2582 2906 2585 3083
rect 2546 2903 2585 2906
rect 2482 2793 2493 2796
rect 2498 2843 2509 2846
rect 2498 2793 2501 2843
rect 2538 2826 2541 2846
rect 2522 2813 2525 2826
rect 2538 2823 2557 2826
rect 2538 2813 2541 2823
rect 2546 2806 2549 2816
rect 2506 2803 2549 2806
rect 2470 2733 2477 2736
rect 2442 2693 2461 2696
rect 2418 2683 2445 2686
rect 2410 2663 2421 2666
rect 2418 2576 2421 2663
rect 2434 2636 2437 2656
rect 2430 2633 2437 2636
rect 2430 2586 2433 2633
rect 2442 2596 2445 2683
rect 2466 2676 2469 2706
rect 2450 2673 2469 2676
rect 2450 2603 2453 2673
rect 2466 2663 2469 2673
rect 2474 2653 2477 2733
rect 2482 2646 2485 2726
rect 2490 2653 2493 2786
rect 2498 2683 2501 2786
rect 2506 2733 2509 2803
rect 2554 2753 2557 2823
rect 2562 2803 2565 2826
rect 2570 2756 2573 2866
rect 2578 2806 2581 2903
rect 2594 2896 2597 3113
rect 2602 2923 2605 3096
rect 2610 3003 2613 3066
rect 2618 2936 2621 3126
rect 2642 3113 2645 3286
rect 2626 3016 2629 3046
rect 2650 3043 2653 3226
rect 2658 3093 2661 3216
rect 2666 3073 2669 3326
rect 2674 3263 2677 3333
rect 2682 3323 2685 3396
rect 2730 3343 2757 3346
rect 2730 3333 2733 3343
rect 2674 3133 2677 3206
rect 2706 3203 2709 3226
rect 2714 3213 2717 3326
rect 2738 3323 2741 3336
rect 2746 3323 2749 3336
rect 2754 3333 2757 3343
rect 2762 3266 2765 3326
rect 2794 3293 2797 3336
rect 2818 3323 2821 3336
rect 2722 3213 2733 3216
rect 2738 3203 2741 3266
rect 2746 3263 2765 3266
rect 2746 3186 2749 3263
rect 2754 3236 2757 3256
rect 2754 3233 2765 3236
rect 2738 3183 2749 3186
rect 2682 3113 2685 3136
rect 2682 3073 2685 3106
rect 2690 3056 2693 3126
rect 2698 3096 2701 3146
rect 2706 3113 2709 3126
rect 2738 3116 2741 3183
rect 2762 3166 2765 3233
rect 2794 3203 2797 3246
rect 2818 3203 2821 3316
rect 2826 3253 2829 3396
rect 2858 3323 2869 3326
rect 2858 3306 2861 3323
rect 2850 3303 2861 3306
rect 2850 3246 2853 3303
rect 2850 3243 2861 3246
rect 2754 3163 2765 3166
rect 2754 3126 2757 3163
rect 2762 3133 2765 3146
rect 2754 3123 2761 3126
rect 2722 3113 2741 3116
rect 2698 3093 2709 3096
rect 2682 3053 2693 3056
rect 2650 3033 2661 3036
rect 2626 3013 2637 3016
rect 2658 3013 2661 3026
rect 2642 2943 2645 3006
rect 2594 2893 2605 2896
rect 2586 2823 2589 2856
rect 2578 2803 2585 2806
rect 2562 2753 2573 2756
rect 2562 2746 2565 2753
rect 2522 2743 2565 2746
rect 2474 2643 2485 2646
rect 2458 2603 2461 2616
rect 2442 2593 2469 2596
rect 2430 2583 2437 2586
rect 2410 2573 2421 2576
rect 2410 2523 2413 2573
rect 2418 2523 2429 2526
rect 2426 2513 2429 2523
rect 2394 2503 2405 2506
rect 2402 2426 2405 2503
rect 2394 2423 2405 2426
rect 2394 2396 2397 2423
rect 2410 2403 2421 2406
rect 2378 2393 2397 2396
rect 2378 2196 2381 2393
rect 2386 2353 2421 2356
rect 2386 2303 2389 2346
rect 2386 2213 2397 2216
rect 2378 2193 2397 2196
rect 2354 2143 2365 2146
rect 2370 2113 2373 2126
rect 2378 2103 2381 2146
rect 2386 2123 2389 2186
rect 2394 2096 2397 2193
rect 2402 2183 2405 2256
rect 2410 2213 2413 2266
rect 2418 2233 2421 2353
rect 2426 2316 2429 2446
rect 2434 2333 2437 2583
rect 2458 2556 2461 2576
rect 2454 2553 2461 2556
rect 2442 2503 2445 2516
rect 2454 2466 2457 2553
rect 2466 2526 2469 2593
rect 2474 2536 2477 2643
rect 2498 2556 2501 2606
rect 2506 2603 2509 2696
rect 2498 2553 2505 2556
rect 2482 2543 2493 2546
rect 2474 2533 2485 2536
rect 2466 2523 2477 2526
rect 2482 2516 2485 2533
rect 2466 2473 2469 2516
rect 2474 2513 2485 2516
rect 2490 2513 2493 2543
rect 2454 2463 2461 2466
rect 2458 2416 2461 2463
rect 2442 2333 2445 2416
rect 2458 2413 2465 2416
rect 2450 2343 2453 2406
rect 2462 2326 2465 2413
rect 2462 2323 2469 2326
rect 2426 2313 2437 2316
rect 2434 2226 2437 2313
rect 2458 2293 2461 2316
rect 2426 2223 2437 2226
rect 2426 2186 2429 2223
rect 2450 2203 2453 2266
rect 2458 2213 2461 2226
rect 2466 2206 2469 2323
rect 2474 2213 2477 2513
rect 2502 2506 2505 2553
rect 2498 2503 2505 2506
rect 2482 2386 2485 2456
rect 2498 2403 2501 2503
rect 2514 2416 2517 2736
rect 2522 2596 2525 2743
rect 2530 2733 2557 2736
rect 2530 2683 2533 2733
rect 2546 2706 2549 2726
rect 2562 2723 2565 2736
rect 2570 2723 2573 2746
rect 2582 2716 2585 2803
rect 2578 2713 2585 2716
rect 2546 2703 2565 2706
rect 2530 2623 2533 2646
rect 2538 2613 2541 2636
rect 2554 2623 2557 2696
rect 2562 2683 2565 2703
rect 2578 2613 2581 2713
rect 2594 2696 2597 2886
rect 2602 2836 2605 2893
rect 2610 2843 2613 2936
rect 2618 2933 2637 2936
rect 2618 2923 2629 2926
rect 2602 2833 2629 2836
rect 2602 2813 2605 2826
rect 2590 2693 2597 2696
rect 2590 2616 2593 2693
rect 2602 2686 2605 2736
rect 2610 2693 2613 2826
rect 2602 2683 2613 2686
rect 2602 2623 2605 2666
rect 2590 2613 2597 2616
rect 2610 2613 2613 2683
rect 2618 2623 2621 2826
rect 2626 2723 2629 2833
rect 2634 2646 2637 2933
rect 2642 2823 2645 2926
rect 2650 2813 2653 2936
rect 2666 2923 2669 3016
rect 2682 2916 2685 3053
rect 2706 3046 2709 3093
rect 2698 3043 2709 3046
rect 2698 2926 2701 3043
rect 2722 3036 2725 3113
rect 2722 3033 2733 3036
rect 2730 3016 2733 3033
rect 2722 3013 2733 3016
rect 2738 3013 2741 3106
rect 2758 3046 2761 3123
rect 2770 3113 2773 3136
rect 2770 3053 2773 3076
rect 2758 3043 2765 3046
rect 2698 2923 2709 2926
rect 2658 2883 2661 2916
rect 2682 2913 2693 2916
rect 2666 2893 2669 2906
rect 2642 2663 2645 2736
rect 2650 2733 2653 2786
rect 2658 2773 2661 2826
rect 2666 2766 2669 2816
rect 2674 2803 2677 2846
rect 2682 2796 2685 2856
rect 2690 2823 2693 2913
rect 2714 2843 2717 2916
rect 2722 2903 2725 2936
rect 2746 2933 2749 3016
rect 2754 2926 2757 3026
rect 2746 2923 2757 2926
rect 2682 2793 2693 2796
rect 2658 2763 2669 2766
rect 2650 2713 2653 2726
rect 2522 2593 2533 2596
rect 2530 2466 2533 2593
rect 2546 2516 2549 2586
rect 2578 2553 2581 2606
rect 2522 2463 2533 2466
rect 2542 2513 2549 2516
rect 2554 2543 2589 2546
rect 2522 2443 2525 2463
rect 2542 2446 2545 2513
rect 2542 2443 2549 2446
rect 2506 2413 2517 2416
rect 2530 2406 2533 2416
rect 2538 2413 2541 2426
rect 2522 2403 2533 2406
rect 2482 2383 2493 2386
rect 2490 2276 2493 2383
rect 2482 2273 2493 2276
rect 2458 2203 2469 2206
rect 2426 2183 2437 2186
rect 2402 2113 2405 2136
rect 2418 2123 2421 2176
rect 2434 2136 2437 2183
rect 2458 2146 2461 2203
rect 2426 2133 2437 2136
rect 2454 2143 2461 2146
rect 2426 2113 2429 2133
rect 2454 2096 2457 2143
rect 2466 2123 2469 2136
rect 2466 2103 2469 2116
rect 2394 2093 2405 2096
rect 2342 2083 2349 2086
rect 2362 2083 2373 2086
rect 2342 2026 2345 2083
rect 2314 1883 2317 1916
rect 2306 1863 2317 1866
rect 2314 1796 2317 1863
rect 2330 1846 2333 2026
rect 2342 2023 2349 2026
rect 2346 2003 2349 2023
rect 2354 2016 2357 2076
rect 2354 2013 2365 2016
rect 2370 2003 2373 2083
rect 2386 2023 2389 2056
rect 2402 2016 2405 2093
rect 2394 2013 2405 2016
rect 2434 2013 2437 2056
rect 2338 1953 2341 1996
rect 2346 1923 2349 1936
rect 2346 1903 2349 1916
rect 2354 1913 2357 1936
rect 2306 1793 2317 1796
rect 2326 1843 2333 1846
rect 2306 1773 2309 1793
rect 2290 1753 2301 1756
rect 2274 1733 2285 1736
rect 2282 1676 2285 1733
rect 2262 1673 2269 1676
rect 2274 1673 2285 1676
rect 2250 1603 2253 1636
rect 2262 1576 2265 1673
rect 2262 1573 2269 1576
rect 2274 1573 2277 1673
rect 2298 1656 2301 1753
rect 2326 1736 2329 1843
rect 2338 1776 2341 1836
rect 2346 1796 2349 1816
rect 2354 1803 2357 1816
rect 2362 1813 2365 1926
rect 2378 1816 2381 1906
rect 2378 1813 2389 1816
rect 2378 1796 2381 1806
rect 2346 1793 2381 1796
rect 2338 1773 2373 1776
rect 2326 1733 2333 1736
rect 2322 1693 2325 1716
rect 2290 1653 2301 1656
rect 2242 1553 2261 1556
rect 2170 1473 2197 1476
rect 2170 1383 2173 1473
rect 2178 1413 2181 1446
rect 2194 1436 2197 1446
rect 2186 1433 2197 1436
rect 2186 1413 2189 1433
rect 2194 1406 2197 1416
rect 2186 1403 2197 1406
rect 2170 1183 2173 1346
rect 2162 1173 2169 1176
rect 2166 1106 2169 1173
rect 2178 1143 2181 1366
rect 2186 1133 2189 1403
rect 2202 1363 2205 1536
rect 2214 1476 2217 1553
rect 2214 1473 2221 1476
rect 2210 1336 2213 1456
rect 2218 1343 2221 1473
rect 2226 1403 2229 1546
rect 2250 1533 2253 1546
rect 2234 1443 2237 1516
rect 2242 1506 2245 1526
rect 2258 1523 2261 1553
rect 2242 1503 2249 1506
rect 2246 1436 2249 1503
rect 2242 1433 2249 1436
rect 2234 1373 2237 1406
rect 2242 1346 2245 1433
rect 2234 1343 2245 1346
rect 2194 1283 2197 1326
rect 2202 1323 2205 1336
rect 2210 1333 2221 1336
rect 2194 1183 2197 1236
rect 2202 1223 2205 1266
rect 2218 1246 2221 1333
rect 2218 1243 2229 1246
rect 2226 1223 2229 1243
rect 2234 1216 2237 1343
rect 2250 1336 2253 1346
rect 2242 1333 2253 1336
rect 2258 1333 2261 1456
rect 2250 1283 2253 1326
rect 2210 1206 2213 1216
rect 2234 1213 2245 1216
rect 2210 1203 2237 1206
rect 2242 1196 2245 1213
rect 2266 1206 2269 1573
rect 2274 1503 2277 1526
rect 2274 1363 2277 1426
rect 2274 1313 2277 1326
rect 2274 1223 2277 1256
rect 2282 1213 2285 1546
rect 2290 1443 2293 1653
rect 2306 1613 2309 1626
rect 2314 1603 2317 1636
rect 2298 1543 2301 1596
rect 2322 1593 2325 1626
rect 2330 1576 2333 1733
rect 2338 1676 2341 1746
rect 2346 1683 2349 1736
rect 2338 1673 2349 1676
rect 2306 1573 2333 1576
rect 2306 1553 2309 1573
rect 2306 1473 2309 1536
rect 2322 1513 2325 1566
rect 2330 1466 2333 1536
rect 2338 1513 2341 1606
rect 2298 1463 2333 1466
rect 2298 1436 2301 1463
rect 2290 1433 2301 1436
rect 2290 1206 2293 1433
rect 2306 1426 2309 1446
rect 2298 1423 2309 1426
rect 2298 1283 2301 1423
rect 2314 1413 2317 1426
rect 2306 1376 2309 1406
rect 2322 1376 2325 1446
rect 2330 1403 2333 1456
rect 2338 1403 2341 1416
rect 2306 1373 2325 1376
rect 2322 1356 2325 1373
rect 2322 1353 2341 1356
rect 2314 1283 2317 1336
rect 2330 1333 2333 1346
rect 2338 1333 2341 1353
rect 2322 1303 2325 1326
rect 2346 1276 2349 1673
rect 2354 1533 2357 1746
rect 2354 1453 2357 1526
rect 2362 1486 2365 1736
rect 2370 1733 2373 1773
rect 2386 1726 2389 1813
rect 2370 1723 2389 1726
rect 2370 1623 2373 1723
rect 2378 1583 2381 1716
rect 2386 1603 2389 1706
rect 2370 1533 2373 1546
rect 2378 1493 2381 1526
rect 2362 1483 2381 1486
rect 2354 1393 2357 1416
rect 2306 1273 2349 1276
rect 2306 1216 2309 1273
rect 2306 1213 2313 1216
rect 2330 1213 2333 1246
rect 2266 1203 2277 1206
rect 2282 1203 2293 1206
rect 2226 1193 2245 1196
rect 2194 1143 2205 1146
rect 2162 1103 2169 1106
rect 2162 1036 2165 1103
rect 2178 1073 2181 1126
rect 2202 1106 2205 1143
rect 2194 1103 2205 1106
rect 2194 1046 2197 1103
rect 2194 1043 2205 1046
rect 2162 1033 2173 1036
rect 2146 1023 2153 1026
rect 2150 946 2153 1023
rect 2162 1003 2165 1016
rect 2146 943 2153 946
rect 2106 843 2117 846
rect 2082 723 2085 736
rect 2098 733 2101 816
rect 2026 713 2053 716
rect 2074 713 2085 716
rect 2018 693 2029 696
rect 2026 626 2029 693
rect 2018 623 2029 626
rect 2042 623 2053 626
rect 2010 533 2013 606
rect 2018 516 2021 623
rect 2042 613 2053 616
rect 2010 513 2021 516
rect 2010 436 2013 513
rect 2026 493 2029 606
rect 2042 596 2045 613
rect 2038 593 2045 596
rect 2038 536 2041 593
rect 2050 573 2053 606
rect 2038 533 2045 536
rect 2034 503 2037 516
rect 2042 453 2045 533
rect 2050 493 2053 526
rect 2058 523 2061 606
rect 2066 533 2069 586
rect 2074 533 2077 713
rect 2098 706 2101 726
rect 2094 703 2101 706
rect 2094 626 2097 703
rect 2106 636 2109 843
rect 2130 826 2133 936
rect 2114 823 2133 826
rect 2114 693 2117 823
rect 2122 806 2125 816
rect 2130 813 2133 823
rect 2122 803 2133 806
rect 2122 726 2125 766
rect 2138 746 2141 936
rect 2146 903 2149 943
rect 2170 933 2173 1033
rect 2178 1023 2197 1026
rect 2178 933 2181 1006
rect 2194 1003 2197 1023
rect 2202 996 2205 1043
rect 2210 1016 2213 1166
rect 2226 1106 2229 1193
rect 2258 1163 2277 1166
rect 2234 1133 2237 1146
rect 2258 1133 2261 1163
rect 2266 1133 2269 1156
rect 2242 1123 2261 1126
rect 2226 1103 2237 1106
rect 2210 1013 2221 1016
rect 2194 993 2205 996
rect 2210 993 2213 1006
rect 2154 923 2181 926
rect 2170 906 2173 923
rect 2186 916 2189 976
rect 2194 933 2197 993
rect 2218 976 2221 1013
rect 2234 986 2237 1103
rect 2258 1003 2261 1096
rect 2266 1083 2269 1116
rect 2274 1113 2277 1163
rect 2266 996 2269 1076
rect 2274 1023 2277 1056
rect 2214 973 2221 976
rect 2226 983 2237 986
rect 2258 993 2269 996
rect 2274 993 2277 1016
rect 2282 1013 2285 1203
rect 2298 1146 2301 1206
rect 2290 1143 2301 1146
rect 2310 1146 2313 1213
rect 2322 1163 2325 1206
rect 2338 1203 2341 1266
rect 2346 1223 2349 1246
rect 2354 1153 2357 1296
rect 2362 1146 2365 1426
rect 2310 1143 2317 1146
rect 2290 1106 2293 1143
rect 2298 1113 2301 1136
rect 2290 1103 2301 1106
rect 2162 903 2173 906
rect 2178 913 2189 916
rect 2162 836 2165 903
rect 2162 833 2173 836
rect 2146 813 2165 816
rect 2154 783 2157 806
rect 2162 803 2165 813
rect 2170 756 2173 833
rect 2154 753 2173 756
rect 2138 743 2149 746
rect 2122 723 2133 726
rect 2138 703 2141 736
rect 2146 723 2149 743
rect 2154 686 2157 753
rect 2178 746 2181 913
rect 2194 896 2197 926
rect 2190 893 2197 896
rect 2190 836 2193 893
rect 2202 846 2205 936
rect 2214 876 2217 973
rect 2226 933 2229 983
rect 2226 893 2229 916
rect 2214 873 2221 876
rect 2218 856 2221 873
rect 2218 853 2229 856
rect 2242 853 2245 926
rect 2250 923 2253 966
rect 2202 843 2221 846
rect 2190 833 2197 836
rect 2194 816 2197 833
rect 2210 823 2213 836
rect 2162 743 2181 746
rect 2162 723 2165 743
rect 2178 723 2181 736
rect 2186 723 2189 816
rect 2194 813 2213 816
rect 2202 803 2213 806
rect 2218 796 2221 843
rect 2226 813 2229 853
rect 2234 813 2237 846
rect 2250 806 2253 846
rect 2234 803 2253 806
rect 2210 793 2221 796
rect 2202 726 2205 736
rect 2210 733 2213 793
rect 2218 783 2221 793
rect 2258 786 2261 993
rect 2282 963 2285 1006
rect 2266 933 2269 946
rect 2290 926 2293 1096
rect 2298 1073 2301 1103
rect 2314 1066 2317 1143
rect 2330 1143 2349 1146
rect 2330 1133 2333 1143
rect 2306 1063 2317 1066
rect 2298 1003 2301 1016
rect 2274 923 2293 926
rect 2274 836 2277 923
rect 2298 913 2301 936
rect 2306 923 2309 1063
rect 2322 1013 2325 1026
rect 2314 933 2317 1006
rect 2322 923 2325 946
rect 2314 876 2317 916
rect 2254 783 2261 786
rect 2270 833 2277 836
rect 2298 873 2317 876
rect 2226 733 2237 736
rect 2242 733 2245 766
rect 2194 723 2205 726
rect 2194 713 2197 723
rect 2154 683 2165 686
rect 2106 633 2113 636
rect 2082 613 2085 626
rect 2094 623 2101 626
rect 2090 573 2093 606
rect 2026 443 2061 446
rect 2010 433 2021 436
rect 1938 413 1957 416
rect 1938 406 1941 413
rect 1906 403 1917 406
rect 1922 403 1941 406
rect 1914 396 1917 403
rect 1946 396 1949 406
rect 1962 403 1965 416
rect 1898 393 1909 396
rect 1914 393 1949 396
rect 1762 273 1797 276
rect 1690 233 1717 236
rect 1714 203 1717 233
rect 1674 133 1677 176
rect 1714 143 1733 146
rect 1698 133 1709 136
rect 1690 113 1693 126
rect 1706 93 1709 116
rect 1722 103 1725 136
rect 1730 0 1733 143
rect 1746 53 1749 216
rect 1794 213 1797 273
rect 1802 213 1805 276
rect 1754 143 1789 146
rect 1754 123 1757 143
rect 1802 136 1805 146
rect 1770 133 1805 136
rect 1810 133 1837 136
rect 1842 133 1845 156
rect 1866 143 1869 316
rect 1890 223 1893 316
rect 1882 196 1885 206
rect 1890 203 1893 216
rect 1898 203 1901 366
rect 1922 323 1925 346
rect 1946 333 1949 356
rect 1954 323 1957 396
rect 2010 353 2013 416
rect 2018 413 2021 433
rect 2026 423 2029 443
rect 2026 336 2029 406
rect 2034 363 2037 436
rect 2042 423 2045 436
rect 2058 423 2061 443
rect 2066 433 2069 516
rect 2098 503 2101 623
rect 2110 556 2113 633
rect 2106 553 2113 556
rect 2122 556 2125 616
rect 2130 583 2133 616
rect 2146 606 2149 626
rect 2154 613 2157 676
rect 2146 603 2157 606
rect 2122 553 2141 556
rect 2042 356 2045 416
rect 2066 413 2069 426
rect 2106 413 2109 553
rect 2114 533 2125 536
rect 2138 533 2141 553
rect 2114 523 2117 533
rect 2146 523 2149 556
rect 2154 516 2157 603
rect 2162 523 2165 683
rect 2170 613 2173 626
rect 2178 613 2181 646
rect 2186 613 2189 696
rect 2202 653 2205 716
rect 2218 713 2221 726
rect 2186 536 2189 606
rect 2202 603 2205 626
rect 2210 593 2213 606
rect 2218 546 2221 616
rect 2234 573 2237 626
rect 2242 603 2245 716
rect 2254 656 2257 783
rect 2270 776 2273 833
rect 2298 816 2301 873
rect 2290 813 2301 816
rect 2282 803 2301 806
rect 2306 803 2309 856
rect 2330 826 2333 1126
rect 2338 1123 2341 1136
rect 2346 1123 2349 1143
rect 2354 1143 2365 1146
rect 2338 1033 2341 1066
rect 2354 1056 2357 1143
rect 2362 1123 2365 1143
rect 2370 1116 2373 1476
rect 2378 1446 2381 1483
rect 2386 1453 2389 1536
rect 2378 1443 2389 1446
rect 2378 1163 2381 1416
rect 2386 1393 2389 1443
rect 2394 1336 2397 2013
rect 2402 1986 2405 1996
rect 2402 1983 2421 1986
rect 2418 1933 2421 1983
rect 2426 1933 2429 1986
rect 2442 1956 2445 2096
rect 2454 2093 2461 2096
rect 2450 2026 2453 2076
rect 2458 2033 2461 2093
rect 2450 2023 2461 2026
rect 2466 2023 2469 2086
rect 2450 1993 2453 2016
rect 2442 1953 2449 1956
rect 2402 1923 2421 1926
rect 2418 1903 2421 1916
rect 2434 1903 2437 1946
rect 2402 1803 2405 1816
rect 2426 1813 2429 1866
rect 2434 1796 2437 1856
rect 2402 1786 2405 1796
rect 2410 1793 2437 1796
rect 2402 1783 2429 1786
rect 2402 1613 2405 1736
rect 2402 1533 2405 1606
rect 2410 1593 2413 1626
rect 2418 1613 2421 1766
rect 2426 1723 2429 1783
rect 2434 1743 2437 1776
rect 2446 1756 2449 1953
rect 2442 1753 2449 1756
rect 2442 1666 2445 1753
rect 2458 1673 2461 2023
rect 2474 2006 2477 2166
rect 2482 2083 2485 2273
rect 2490 2076 2493 2216
rect 2498 2096 2501 2256
rect 2506 2213 2509 2316
rect 2514 2286 2517 2326
rect 2522 2303 2525 2403
rect 2538 2393 2541 2406
rect 2530 2303 2533 2316
rect 2538 2293 2541 2336
rect 2546 2303 2549 2443
rect 2514 2283 2521 2286
rect 2554 2283 2557 2543
rect 2578 2533 2581 2543
rect 2586 2533 2589 2543
rect 2562 2523 2573 2526
rect 2578 2503 2581 2526
rect 2594 2496 2597 2613
rect 2626 2603 2629 2646
rect 2634 2643 2645 2646
rect 2602 2503 2605 2536
rect 2610 2523 2613 2546
rect 2618 2496 2621 2566
rect 2642 2536 2645 2643
rect 2658 2636 2661 2763
rect 2674 2733 2677 2766
rect 2666 2716 2669 2726
rect 2682 2723 2685 2786
rect 2690 2723 2693 2793
rect 2698 2776 2701 2806
rect 2722 2803 2725 2816
rect 2730 2806 2733 2826
rect 2746 2813 2749 2923
rect 2730 2803 2749 2806
rect 2706 2793 2733 2796
rect 2698 2773 2705 2776
rect 2702 2716 2705 2773
rect 2666 2713 2693 2716
rect 2698 2713 2705 2716
rect 2698 2696 2701 2713
rect 2682 2693 2701 2696
rect 2682 2676 2685 2693
rect 2678 2673 2685 2676
rect 2658 2633 2669 2636
rect 2666 2613 2669 2633
rect 2666 2573 2669 2606
rect 2678 2566 2681 2673
rect 2690 2623 2693 2686
rect 2714 2626 2717 2726
rect 2722 2703 2725 2726
rect 2730 2713 2733 2793
rect 2746 2753 2749 2803
rect 2754 2776 2757 2846
rect 2762 2823 2765 3043
rect 2770 2843 2773 3046
rect 2770 2813 2773 2826
rect 2770 2783 2773 2796
rect 2754 2773 2773 2776
rect 2738 2706 2741 2736
rect 2762 2713 2765 2726
rect 2770 2723 2773 2773
rect 2730 2703 2741 2706
rect 2698 2623 2717 2626
rect 2582 2493 2597 2496
rect 2614 2493 2621 2496
rect 2638 2533 2645 2536
rect 2666 2563 2681 2566
rect 2518 2206 2521 2283
rect 2562 2273 2565 2436
rect 2570 2403 2573 2446
rect 2582 2436 2585 2493
rect 2578 2433 2585 2436
rect 2614 2436 2617 2493
rect 2614 2433 2621 2436
rect 2578 2413 2581 2433
rect 2578 2346 2581 2366
rect 2594 2353 2597 2426
rect 2578 2343 2585 2346
rect 2570 2246 2573 2336
rect 2582 2246 2585 2343
rect 2594 2323 2597 2346
rect 2538 2243 2573 2246
rect 2578 2243 2585 2246
rect 2514 2203 2521 2206
rect 2530 2203 2533 2226
rect 2538 2213 2541 2243
rect 2546 2213 2557 2216
rect 2562 2203 2565 2236
rect 2506 2133 2509 2156
rect 2514 2143 2517 2203
rect 2570 2193 2573 2206
rect 2514 2113 2517 2136
rect 2498 2093 2509 2096
rect 2490 2073 2497 2076
rect 2470 2003 2477 2006
rect 2470 1876 2473 2003
rect 2470 1873 2477 1876
rect 2474 1853 2477 1873
rect 2466 1763 2469 1806
rect 2474 1766 2477 1786
rect 2482 1773 2485 2056
rect 2494 1986 2497 2073
rect 2490 1983 2497 1986
rect 2490 1873 2493 1983
rect 2506 1966 2509 2093
rect 2530 2013 2533 2146
rect 2498 1963 2509 1966
rect 2498 1926 2501 1963
rect 2522 1956 2525 2006
rect 2522 1953 2533 1956
rect 2506 1943 2525 1946
rect 2506 1933 2509 1943
rect 2498 1923 2509 1926
rect 2490 1783 2493 1816
rect 2498 1766 2501 1923
rect 2514 1913 2517 1936
rect 2522 1923 2525 1943
rect 2530 1933 2533 1953
rect 2538 1923 2541 2056
rect 2546 2013 2549 2026
rect 2546 1913 2549 1976
rect 2546 1893 2549 1906
rect 2506 1803 2509 1816
rect 2514 1813 2517 1886
rect 2530 1823 2549 1826
rect 2530 1813 2533 1823
rect 2522 1783 2525 1806
rect 2474 1763 2485 1766
rect 2498 1763 2525 1766
rect 2490 1753 2517 1756
rect 2466 1743 2477 1746
rect 2466 1666 2469 1726
rect 2442 1663 2453 1666
rect 2426 1613 2437 1616
rect 2426 1593 2429 1606
rect 2442 1603 2445 1646
rect 2402 1503 2405 1526
rect 2410 1453 2413 1556
rect 2418 1473 2421 1516
rect 2426 1436 2429 1526
rect 2402 1433 2429 1436
rect 2402 1423 2405 1433
rect 2418 1413 2421 1426
rect 2402 1403 2413 1406
rect 2402 1386 2405 1403
rect 2426 1396 2429 1416
rect 2410 1393 2429 1396
rect 2402 1383 2413 1386
rect 2394 1333 2401 1336
rect 2386 1313 2389 1326
rect 2386 1233 2389 1306
rect 2398 1226 2401 1333
rect 2410 1323 2413 1383
rect 2418 1283 2421 1336
rect 2410 1233 2413 1266
rect 2386 1203 2389 1226
rect 2394 1223 2401 1226
rect 2346 1053 2357 1056
rect 2366 1113 2373 1116
rect 2338 913 2341 926
rect 2346 916 2349 1053
rect 2366 1036 2369 1113
rect 2378 1093 2381 1156
rect 2362 1033 2369 1036
rect 2362 1013 2365 1033
rect 2378 963 2381 1026
rect 2354 923 2357 956
rect 2386 933 2389 1126
rect 2346 913 2357 916
rect 2322 823 2333 826
rect 2322 816 2325 823
rect 2314 813 2325 816
rect 2266 773 2273 776
rect 2254 653 2261 656
rect 2218 543 2229 546
rect 2114 503 2117 516
rect 2122 513 2133 516
rect 2154 513 2165 516
rect 2138 413 2141 426
rect 2146 413 2149 426
rect 1986 333 2029 336
rect 2034 353 2045 356
rect 2034 326 2037 353
rect 2066 343 2069 406
rect 2114 403 2133 406
rect 2074 343 2077 366
rect 2050 333 2061 336
rect 1938 313 1973 316
rect 2002 286 2005 326
rect 1994 283 2005 286
rect 1906 196 1909 206
rect 1938 196 1941 216
rect 1954 203 1957 216
rect 1962 213 1981 216
rect 1962 203 1965 213
rect 1970 203 1989 206
rect 1882 193 1909 196
rect 1906 183 1909 193
rect 1930 193 1941 196
rect 1930 146 1933 193
rect 1930 143 1941 146
rect 1850 133 1885 136
rect 1890 133 1901 136
rect 1770 123 1781 126
rect 1786 0 1789 133
rect 1794 123 1829 126
rect 1834 103 1837 133
rect 1850 103 1853 133
rect 1938 126 1941 143
rect 1946 133 1949 156
rect 1970 146 1973 203
rect 1962 143 1973 146
rect 1858 123 1885 126
rect 1938 123 1957 126
rect 1882 116 1885 123
rect 1858 83 1861 116
rect 1874 63 1877 116
rect 1882 113 1917 116
rect 1914 83 1917 106
rect 1946 93 1949 116
rect 1954 83 1957 123
rect 1962 63 1965 143
rect 1970 103 1973 136
rect 1978 123 1981 196
rect 1986 173 1989 203
rect 1994 166 1997 283
rect 2010 276 2013 326
rect 2034 323 2053 326
rect 2090 323 2093 336
rect 2106 306 2109 336
rect 2002 273 2013 276
rect 2002 203 2005 273
rect 2018 243 2021 306
rect 2098 303 2109 306
rect 2098 256 2101 303
rect 2122 263 2125 336
rect 2162 316 2165 513
rect 2170 503 2173 536
rect 2186 533 2213 536
rect 2170 403 2173 416
rect 2186 413 2189 526
rect 2218 523 2221 536
rect 2226 483 2229 543
rect 2250 513 2253 636
rect 2258 593 2261 653
rect 2234 443 2253 446
rect 2194 413 2197 426
rect 2234 413 2237 443
rect 2242 406 2245 436
rect 2250 423 2253 443
rect 2258 413 2261 536
rect 2266 473 2269 773
rect 2274 603 2277 616
rect 2282 613 2285 726
rect 2298 723 2301 803
rect 2306 733 2309 786
rect 2314 726 2317 813
rect 2322 796 2325 806
rect 2330 803 2333 816
rect 2338 813 2341 836
rect 2338 796 2341 806
rect 2346 796 2349 806
rect 2322 793 2349 796
rect 2354 776 2357 913
rect 2370 823 2381 826
rect 2362 786 2365 806
rect 2370 803 2373 816
rect 2378 803 2381 816
rect 2386 786 2389 836
rect 2362 783 2389 786
rect 2354 773 2381 776
rect 2354 733 2357 766
rect 2362 733 2373 736
rect 2314 723 2325 726
rect 2306 686 2309 716
rect 2322 703 2325 723
rect 2330 693 2333 716
rect 2362 686 2365 726
rect 2378 723 2381 773
rect 2306 683 2365 686
rect 2298 586 2301 636
rect 2306 626 2309 656
rect 2306 623 2317 626
rect 2322 613 2325 656
rect 2338 613 2341 676
rect 2386 653 2389 783
rect 2394 646 2397 1223
rect 2402 956 2405 1206
rect 2418 1163 2421 1226
rect 2410 1013 2413 1116
rect 2418 1113 2421 1156
rect 2426 1133 2429 1336
rect 2434 1123 2437 1556
rect 2450 1523 2453 1663
rect 2458 1663 2469 1666
rect 2442 1443 2445 1516
rect 2450 1493 2453 1506
rect 2458 1486 2461 1663
rect 2466 1633 2469 1656
rect 2474 1643 2477 1743
rect 2482 1733 2485 1746
rect 2490 1733 2493 1753
rect 2506 1733 2509 1746
rect 2514 1733 2517 1753
rect 2482 1713 2485 1726
rect 2466 1603 2469 1616
rect 2466 1513 2469 1546
rect 2474 1503 2477 1536
rect 2482 1523 2485 1706
rect 2498 1693 2501 1726
rect 2490 1513 2493 1676
rect 2514 1636 2517 1726
rect 2522 1713 2525 1763
rect 2530 1696 2533 1806
rect 2538 1743 2541 1816
rect 2538 1703 2541 1736
rect 2546 1723 2549 1823
rect 2554 1733 2557 2156
rect 2562 2133 2573 2136
rect 2570 2103 2573 2126
rect 2562 1933 2565 2016
rect 2570 1993 2573 2006
rect 2578 1923 2581 2243
rect 2594 2156 2597 2286
rect 2602 2253 2605 2326
rect 2610 2236 2613 2416
rect 2618 2383 2621 2433
rect 2626 2393 2629 2486
rect 2638 2446 2641 2533
rect 2666 2516 2669 2563
rect 2674 2523 2685 2526
rect 2690 2523 2693 2606
rect 2698 2516 2701 2623
rect 2706 2613 2725 2616
rect 2706 2603 2709 2613
rect 2706 2523 2709 2596
rect 2714 2533 2717 2586
rect 2634 2443 2641 2446
rect 2618 2323 2621 2336
rect 2626 2306 2629 2336
rect 2634 2316 2637 2443
rect 2642 2353 2645 2426
rect 2642 2323 2645 2346
rect 2650 2316 2653 2476
rect 2658 2333 2661 2516
rect 2666 2513 2677 2516
rect 2666 2413 2669 2466
rect 2674 2406 2677 2513
rect 2682 2476 2685 2516
rect 2690 2503 2693 2516
rect 2698 2513 2709 2516
rect 2682 2473 2701 2476
rect 2666 2403 2677 2406
rect 2634 2313 2645 2316
rect 2650 2313 2657 2316
rect 2622 2303 2629 2306
rect 2622 2246 2625 2303
rect 2606 2233 2613 2236
rect 2618 2243 2625 2246
rect 2606 2176 2609 2233
rect 2606 2173 2613 2176
rect 2594 2153 2605 2156
rect 2586 2053 2589 2126
rect 2594 2046 2597 2136
rect 2602 2103 2605 2153
rect 2602 2083 2605 2096
rect 2586 2043 2597 2046
rect 2586 2023 2589 2043
rect 2602 2023 2605 2036
rect 2578 1883 2581 1916
rect 2570 1813 2581 1816
rect 2586 1806 2589 1986
rect 2594 1813 2597 1916
rect 2602 1836 2605 1996
rect 2610 1883 2613 2173
rect 2618 1843 2621 2243
rect 2626 2203 2629 2236
rect 2626 2053 2629 2126
rect 2634 2116 2637 2306
rect 2642 2153 2645 2313
rect 2654 2246 2657 2313
rect 2650 2243 2657 2246
rect 2634 2113 2641 2116
rect 2602 1833 2621 1836
rect 2578 1803 2589 1806
rect 2554 1706 2557 1726
rect 2550 1703 2557 1706
rect 2506 1633 2517 1636
rect 2526 1693 2533 1696
rect 2498 1613 2501 1626
rect 2506 1603 2509 1633
rect 2526 1626 2529 1693
rect 2514 1596 2517 1626
rect 2526 1623 2533 1626
rect 2530 1603 2533 1623
rect 2514 1593 2533 1596
rect 2450 1483 2461 1486
rect 2442 1403 2445 1436
rect 2442 1343 2445 1396
rect 2450 1353 2453 1483
rect 2458 1346 2461 1466
rect 2466 1463 2477 1466
rect 2482 1463 2501 1466
rect 2466 1415 2469 1463
rect 2482 1423 2485 1463
rect 2466 1412 2484 1415
rect 2466 1403 2485 1406
rect 2466 1383 2469 1403
rect 2450 1343 2461 1346
rect 2442 1323 2445 1336
rect 2442 1136 2445 1316
rect 2450 1286 2453 1343
rect 2458 1293 2461 1336
rect 2466 1306 2469 1376
rect 2474 1323 2477 1396
rect 2466 1303 2473 1306
rect 2450 1283 2461 1286
rect 2450 1256 2453 1276
rect 2458 1263 2461 1283
rect 2450 1253 2461 1256
rect 2458 1213 2461 1253
rect 2470 1226 2473 1303
rect 2466 1223 2473 1226
rect 2450 1156 2453 1206
rect 2450 1153 2461 1156
rect 2442 1133 2461 1136
rect 2442 1116 2445 1133
rect 2426 1113 2445 1116
rect 2418 1093 2421 1106
rect 2418 1003 2421 1026
rect 2426 1013 2429 1113
rect 2442 1093 2445 1106
rect 2434 1023 2445 1026
rect 2402 953 2421 956
rect 2402 933 2405 946
rect 2410 913 2413 926
rect 2418 896 2421 953
rect 2426 933 2429 966
rect 2450 943 2453 1126
rect 2458 1003 2461 1056
rect 2434 916 2437 936
rect 2414 893 2421 896
rect 2426 913 2437 916
rect 2442 913 2445 936
rect 2450 913 2453 926
rect 2466 923 2469 1223
rect 2482 1213 2485 1403
rect 2490 1333 2493 1456
rect 2498 1446 2501 1463
rect 2506 1453 2509 1526
rect 2514 1523 2517 1546
rect 2522 1533 2525 1586
rect 2530 1523 2533 1593
rect 2498 1443 2509 1446
rect 2498 1416 2501 1426
rect 2506 1423 2509 1443
rect 2498 1413 2509 1416
rect 2474 1093 2477 1206
rect 2482 1153 2485 1206
rect 2490 1196 2493 1316
rect 2498 1313 2501 1396
rect 2506 1256 2509 1336
rect 2498 1253 2509 1256
rect 2498 1203 2501 1253
rect 2506 1223 2509 1246
rect 2514 1223 2517 1516
rect 2522 1413 2525 1446
rect 2522 1296 2525 1336
rect 2530 1333 2533 1396
rect 2538 1326 2541 1696
rect 2550 1636 2553 1703
rect 2550 1633 2557 1636
rect 2554 1613 2557 1633
rect 2546 1593 2549 1606
rect 2546 1523 2549 1576
rect 2554 1533 2557 1606
rect 2562 1526 2565 1786
rect 2570 1713 2573 1766
rect 2570 1673 2573 1706
rect 2570 1543 2573 1626
rect 2546 1426 2549 1436
rect 2554 1433 2557 1526
rect 2562 1523 2569 1526
rect 2566 1446 2569 1523
rect 2562 1443 2569 1446
rect 2546 1423 2557 1426
rect 2562 1423 2565 1443
rect 2546 1373 2549 1416
rect 2554 1406 2557 1423
rect 2554 1403 2561 1406
rect 2558 1336 2561 1403
rect 2570 1363 2573 1406
rect 2554 1333 2561 1336
rect 2530 1313 2533 1326
rect 2538 1323 2549 1326
rect 2522 1293 2529 1296
rect 2538 1293 2541 1316
rect 2526 1216 2529 1293
rect 2538 1223 2541 1246
rect 2546 1216 2549 1323
rect 2554 1313 2557 1333
rect 2522 1213 2529 1216
rect 2538 1213 2549 1216
rect 2490 1193 2501 1196
rect 2490 1123 2493 1166
rect 2498 1136 2501 1193
rect 2498 1133 2517 1136
rect 2522 1133 2525 1213
rect 2538 1196 2541 1213
rect 2534 1193 2541 1196
rect 2534 1136 2537 1193
rect 2546 1153 2549 1206
rect 2534 1133 2541 1136
rect 2498 1113 2501 1133
rect 2506 1123 2517 1126
rect 2514 1066 2517 1123
rect 2538 1116 2541 1133
rect 2554 1123 2557 1306
rect 2562 1293 2565 1306
rect 2562 1203 2565 1276
rect 2570 1206 2573 1316
rect 2578 1213 2581 1803
rect 2602 1793 2605 1826
rect 2586 1703 2589 1756
rect 2594 1703 2597 1716
rect 2586 1523 2589 1606
rect 2594 1603 2597 1616
rect 2594 1533 2597 1566
rect 2586 1436 2589 1516
rect 2586 1433 2593 1436
rect 2590 1336 2593 1433
rect 2602 1416 2605 1786
rect 2610 1506 2613 1806
rect 2618 1783 2621 1833
rect 2618 1596 2621 1766
rect 2626 1606 2629 2036
rect 2638 2026 2641 2113
rect 2650 2076 2653 2243
rect 2658 2173 2661 2226
rect 2650 2073 2661 2076
rect 2634 2023 2641 2026
rect 2634 1903 2637 2023
rect 2650 2013 2653 2026
rect 2642 1903 2645 2006
rect 2658 1946 2661 2073
rect 2666 2033 2669 2403
rect 2674 2243 2677 2336
rect 2682 2283 2685 2416
rect 2690 2413 2693 2456
rect 2698 2423 2701 2473
rect 2706 2416 2709 2513
rect 2698 2413 2709 2416
rect 2698 2323 2701 2413
rect 2674 2213 2677 2226
rect 2682 2203 2685 2216
rect 2690 2133 2693 2206
rect 2706 2126 2709 2376
rect 2714 2323 2717 2486
rect 2714 2213 2717 2226
rect 2682 2103 2685 2126
rect 2698 2123 2709 2126
rect 2674 2006 2677 2096
rect 2682 2013 2685 2046
rect 2674 2003 2685 2006
rect 2650 1943 2661 1946
rect 2650 1923 2653 1943
rect 2682 1933 2685 2003
rect 2690 1953 2693 2026
rect 2698 2006 2701 2123
rect 2714 2116 2717 2126
rect 2706 2113 2717 2116
rect 2706 2093 2709 2113
rect 2714 2086 2717 2106
rect 2722 2103 2725 2546
rect 2730 2326 2733 2703
rect 2738 2543 2741 2626
rect 2746 2603 2749 2706
rect 2778 2696 2781 3126
rect 2794 3113 2797 3176
rect 2842 3146 2845 3226
rect 2858 3203 2861 3243
rect 2874 3223 2877 3336
rect 2882 3323 2885 3366
rect 2914 3323 2917 3376
rect 2938 3326 2941 3396
rect 2922 3323 2941 3326
rect 2922 3316 2925 3323
rect 2890 3243 2893 3316
rect 2914 3313 2925 3316
rect 2914 3293 2917 3313
rect 2866 3186 2869 3216
rect 2874 3203 2885 3206
rect 2906 3186 2909 3216
rect 2866 3183 2877 3186
rect 2826 3143 2845 3146
rect 2826 3133 2829 3143
rect 2802 3106 2805 3126
rect 2834 3113 2837 3136
rect 2858 3113 2861 3176
rect 2874 3106 2877 3183
rect 2802 3103 2813 3106
rect 2786 3063 2797 3066
rect 2786 2813 2789 3036
rect 2794 3013 2797 3063
rect 2810 3036 2813 3103
rect 2858 3103 2877 3106
rect 2898 3183 2909 3186
rect 2850 3076 2853 3096
rect 2802 3033 2813 3036
rect 2842 3073 2853 3076
rect 2794 2913 2797 2946
rect 2794 2803 2797 2846
rect 2786 2726 2789 2796
rect 2794 2733 2797 2796
rect 2802 2793 2805 3033
rect 2842 3016 2845 3073
rect 2810 3003 2813 3016
rect 2826 3013 2845 3016
rect 2810 2933 2813 2986
rect 2810 2913 2813 2926
rect 2818 2886 2821 2936
rect 2826 2906 2829 3013
rect 2858 3006 2861 3103
rect 2898 3086 2901 3183
rect 2914 3166 2917 3236
rect 2910 3163 2917 3166
rect 2910 3106 2913 3163
rect 2922 3133 2925 3306
rect 2930 3223 2933 3316
rect 2938 3313 2941 3323
rect 2930 3133 2933 3176
rect 2938 3143 2941 3306
rect 2946 3203 2949 3286
rect 2962 3273 2965 3326
rect 2978 3313 2981 3336
rect 2986 3323 2989 3356
rect 2994 3333 2997 3376
rect 3050 3353 3077 3356
rect 3010 3303 3013 3336
rect 2954 3226 2957 3246
rect 3034 3236 3037 3346
rect 3050 3323 3053 3353
rect 3034 3233 3045 3236
rect 3050 3233 3053 3266
rect 2954 3223 2965 3226
rect 2962 3176 2965 3223
rect 2958 3173 2965 3176
rect 2910 3103 2917 3106
rect 2898 3083 2909 3086
rect 2866 3013 2869 3046
rect 2858 3003 2869 3006
rect 2866 2993 2869 3003
rect 2834 2946 2837 2986
rect 2834 2943 2869 2946
rect 2850 2933 2869 2936
rect 2842 2923 2861 2926
rect 2834 2913 2853 2916
rect 2826 2903 2845 2906
rect 2818 2883 2829 2886
rect 2810 2783 2813 2816
rect 2826 2813 2829 2883
rect 2818 2766 2821 2806
rect 2834 2803 2837 2826
rect 2842 2813 2845 2903
rect 2858 2896 2861 2923
rect 2866 2913 2869 2926
rect 2854 2893 2861 2896
rect 2854 2816 2857 2893
rect 2850 2813 2857 2816
rect 2850 2806 2853 2813
rect 2866 2806 2869 2906
rect 2842 2803 2853 2806
rect 2858 2803 2869 2806
rect 2818 2763 2829 2766
rect 2786 2723 2797 2726
rect 2802 2723 2813 2726
rect 2818 2723 2821 2736
rect 2794 2716 2797 2723
rect 2770 2693 2781 2696
rect 2754 2603 2757 2666
rect 2770 2556 2773 2693
rect 2786 2623 2789 2716
rect 2794 2713 2805 2716
rect 2794 2623 2797 2706
rect 2778 2613 2797 2616
rect 2778 2563 2781 2613
rect 2786 2603 2797 2606
rect 2770 2553 2781 2556
rect 2738 2533 2749 2536
rect 2770 2533 2773 2546
rect 2738 2513 2741 2533
rect 2746 2503 2749 2526
rect 2762 2523 2773 2526
rect 2738 2343 2741 2476
rect 2746 2463 2757 2466
rect 2746 2373 2749 2463
rect 2754 2383 2757 2406
rect 2730 2323 2737 2326
rect 2734 2256 2737 2323
rect 2730 2253 2737 2256
rect 2730 2203 2733 2253
rect 2706 2083 2717 2086
rect 2706 2073 2709 2083
rect 2698 2003 2705 2006
rect 2714 2003 2717 2016
rect 2702 1936 2705 2003
rect 2702 1933 2709 1936
rect 2658 1913 2669 1916
rect 2634 1806 2637 1886
rect 2666 1856 2669 1913
rect 2682 1903 2685 1926
rect 2706 1916 2709 1933
rect 2714 1923 2717 1996
rect 2706 1913 2717 1916
rect 2658 1853 2669 1856
rect 2642 1813 2653 1816
rect 2658 1813 2661 1853
rect 2634 1803 2645 1806
rect 2634 1613 2637 1746
rect 2642 1673 2645 1803
rect 2650 1773 2653 1806
rect 2658 1723 2661 1736
rect 2642 1613 2645 1646
rect 2658 1613 2661 1646
rect 2626 1603 2645 1606
rect 2618 1593 2629 1596
rect 2618 1533 2621 1576
rect 2618 1516 2621 1526
rect 2626 1523 2629 1593
rect 2634 1523 2637 1536
rect 2618 1513 2637 1516
rect 2610 1503 2621 1506
rect 2610 1416 2613 1426
rect 2602 1413 2613 1416
rect 2586 1333 2593 1336
rect 2602 1333 2605 1396
rect 2618 1336 2621 1503
rect 2642 1496 2645 1603
rect 2634 1493 2645 1496
rect 2634 1426 2637 1493
rect 2650 1436 2653 1596
rect 2658 1513 2661 1596
rect 2650 1433 2657 1436
rect 2634 1423 2645 1426
rect 2614 1333 2621 1336
rect 2586 1313 2589 1333
rect 2586 1216 2589 1306
rect 2594 1283 2597 1316
rect 2602 1223 2605 1326
rect 2614 1276 2617 1333
rect 2626 1286 2629 1326
rect 2634 1303 2637 1406
rect 2626 1283 2633 1286
rect 2614 1273 2621 1276
rect 2586 1213 2597 1216
rect 2570 1203 2581 1206
rect 2594 1203 2597 1213
rect 2538 1113 2549 1116
rect 2514 1063 2525 1066
rect 2402 813 2405 856
rect 2414 806 2417 893
rect 2426 813 2429 913
rect 2442 813 2445 846
rect 2414 803 2421 806
rect 2402 673 2405 786
rect 2418 733 2421 803
rect 2418 673 2421 726
rect 2434 713 2437 806
rect 2290 583 2301 586
rect 2274 493 2277 536
rect 2290 533 2293 583
rect 2298 526 2301 536
rect 2282 523 2301 526
rect 2266 463 2293 466
rect 2266 453 2269 463
rect 2274 413 2277 426
rect 2234 403 2253 406
rect 2170 323 2173 346
rect 2202 336 2205 356
rect 2194 333 2205 336
rect 2162 313 2173 316
rect 2098 253 2109 256
rect 2018 223 2021 236
rect 2042 203 2045 226
rect 2050 216 2053 246
rect 2058 223 2077 226
rect 2106 223 2109 253
rect 2050 213 2069 216
rect 1994 163 2005 166
rect 1986 83 1989 116
rect 2002 63 2005 163
rect 2034 133 2037 186
rect 2010 103 2013 126
rect 2026 96 2029 126
rect 2042 123 2045 156
rect 2050 133 2053 196
rect 2066 173 2069 206
rect 2050 103 2053 126
rect 2074 113 2077 223
rect 2130 213 2133 276
rect 2146 223 2149 246
rect 2154 243 2165 246
rect 2154 213 2157 243
rect 2170 223 2173 313
rect 2194 216 2197 333
rect 2162 206 2165 216
rect 2194 213 2205 216
rect 2210 213 2213 366
rect 2218 333 2221 356
rect 2250 333 2253 376
rect 2226 323 2237 326
rect 2226 253 2229 323
rect 2250 306 2253 326
rect 2242 303 2253 306
rect 2242 246 2245 303
rect 2242 243 2253 246
rect 2226 213 2245 216
rect 2122 196 2125 206
rect 2154 196 2157 206
rect 2162 203 2181 206
rect 2114 186 2117 196
rect 2122 193 2157 196
rect 2114 183 2125 186
rect 2122 136 2125 183
rect 2122 133 2157 136
rect 2170 133 2173 156
rect 2066 96 2069 106
rect 2026 93 2069 96
rect 2082 96 2085 126
rect 2106 96 2109 106
rect 2082 93 2109 96
rect 2114 93 2117 116
rect 2122 113 2125 133
rect 2130 83 2133 126
rect 2138 123 2157 126
rect 2178 123 2181 203
rect 2202 193 2205 213
rect 2186 133 2189 176
rect 2138 63 2141 123
rect 2146 106 2149 116
rect 2146 103 2165 106
rect 2162 96 2165 103
rect 2194 96 2197 136
rect 2218 123 2221 206
rect 2226 173 2229 213
rect 2234 196 2237 206
rect 2250 203 2253 243
rect 2258 213 2261 366
rect 2266 333 2269 346
rect 2282 333 2285 456
rect 2290 413 2293 463
rect 2298 413 2301 516
rect 2306 463 2309 606
rect 2314 543 2317 606
rect 2330 586 2333 606
rect 2346 603 2349 636
rect 2354 596 2357 646
rect 2378 643 2397 646
rect 2326 583 2333 586
rect 2346 593 2357 596
rect 2314 503 2317 536
rect 2326 506 2329 583
rect 2338 533 2341 556
rect 2346 523 2349 593
rect 2354 533 2357 586
rect 2362 573 2365 636
rect 2362 526 2365 536
rect 2354 523 2365 526
rect 2326 503 2333 506
rect 2330 483 2333 503
rect 2322 413 2325 426
rect 2354 413 2357 523
rect 2370 503 2373 606
rect 2378 576 2381 643
rect 2402 613 2405 656
rect 2410 616 2413 626
rect 2426 623 2429 706
rect 2442 696 2445 736
rect 2450 723 2453 856
rect 2474 846 2477 1026
rect 2498 1013 2501 1026
rect 2522 1023 2525 1063
rect 2546 1036 2549 1113
rect 2546 1033 2557 1036
rect 2506 1013 2517 1016
rect 2530 1013 2549 1016
rect 2482 923 2485 956
rect 2458 843 2477 846
rect 2458 823 2461 843
rect 2466 813 2469 826
rect 2474 773 2477 836
rect 2482 803 2485 826
rect 2490 783 2493 916
rect 2498 873 2501 1006
rect 2530 1003 2533 1013
rect 2554 1003 2557 1033
rect 2458 713 2485 716
rect 2438 693 2445 696
rect 2438 616 2441 693
rect 2410 613 2421 616
rect 2386 603 2397 606
rect 2386 583 2389 603
rect 2378 573 2397 576
rect 2394 526 2397 573
rect 2378 513 2381 526
rect 2386 523 2397 526
rect 2362 423 2365 456
rect 2362 406 2365 416
rect 2274 263 2277 326
rect 2298 296 2301 406
rect 2346 403 2365 406
rect 2306 303 2309 336
rect 2354 333 2357 356
rect 2362 333 2365 346
rect 2370 326 2373 466
rect 2378 376 2381 436
rect 2386 396 2389 416
rect 2394 403 2397 416
rect 2402 413 2405 586
rect 2410 523 2413 606
rect 2418 553 2421 613
rect 2434 613 2441 616
rect 2426 546 2429 596
rect 2418 543 2429 546
rect 2434 543 2437 613
rect 2442 593 2445 606
rect 2450 576 2453 706
rect 2458 696 2461 713
rect 2458 693 2465 696
rect 2482 693 2485 713
rect 2462 606 2465 693
rect 2458 603 2465 606
rect 2458 583 2461 603
rect 2474 576 2477 616
rect 2482 603 2485 616
rect 2450 573 2477 576
rect 2474 563 2477 573
rect 2410 483 2413 516
rect 2418 493 2421 543
rect 2426 533 2469 536
rect 2442 433 2445 526
rect 2450 493 2453 526
rect 2466 513 2469 533
rect 2474 523 2477 556
rect 2482 523 2485 576
rect 2490 533 2493 736
rect 2498 723 2501 846
rect 2506 803 2509 896
rect 2522 813 2525 936
rect 2530 933 2533 996
rect 2562 973 2565 1136
rect 2570 1123 2573 1136
rect 2578 1053 2581 1203
rect 2602 1176 2605 1196
rect 2594 1173 2605 1176
rect 2594 1086 2597 1173
rect 2610 1133 2613 1256
rect 2618 1173 2621 1273
rect 2630 1176 2633 1283
rect 2642 1203 2645 1423
rect 2654 1386 2657 1433
rect 2666 1426 2669 1816
rect 2674 1803 2677 1846
rect 2674 1733 2677 1746
rect 2674 1696 2677 1726
rect 2682 1713 2685 1816
rect 2690 1733 2693 1876
rect 2698 1736 2701 1856
rect 2706 1743 2709 1906
rect 2714 1813 2717 1913
rect 2714 1793 2717 1806
rect 2698 1733 2709 1736
rect 2674 1693 2681 1696
rect 2678 1606 2681 1693
rect 2690 1613 2693 1726
rect 2714 1723 2717 1736
rect 2722 1723 2725 1996
rect 2730 1853 2733 2136
rect 2738 2133 2741 2236
rect 2746 2123 2749 2276
rect 2754 2183 2757 2316
rect 2762 2233 2765 2406
rect 2770 2403 2773 2506
rect 2770 2293 2773 2306
rect 2778 2273 2781 2553
rect 2786 2543 2789 2586
rect 2786 2523 2789 2536
rect 2786 2473 2789 2516
rect 2794 2483 2797 2556
rect 2802 2426 2805 2713
rect 2810 2703 2813 2723
rect 2826 2713 2829 2763
rect 2842 2746 2845 2803
rect 2850 2776 2853 2796
rect 2858 2783 2861 2803
rect 2850 2773 2861 2776
rect 2834 2743 2845 2746
rect 2834 2733 2837 2743
rect 2818 2703 2829 2706
rect 2810 2613 2813 2686
rect 2810 2543 2813 2606
rect 2818 2583 2821 2703
rect 2834 2646 2837 2726
rect 2842 2723 2845 2736
rect 2858 2733 2861 2773
rect 2850 2703 2853 2726
rect 2874 2716 2877 3016
rect 2882 3003 2885 3036
rect 2898 3013 2901 3066
rect 2882 2786 2885 2936
rect 2890 2923 2893 2976
rect 2906 2946 2909 3083
rect 2914 3003 2917 3103
rect 2922 3096 2925 3126
rect 2922 3093 2929 3096
rect 2926 2996 2929 3093
rect 2938 3003 2941 3126
rect 2946 3123 2949 3136
rect 2958 3116 2961 3173
rect 2954 3113 2961 3116
rect 2898 2943 2909 2946
rect 2922 2993 2929 2996
rect 2922 2946 2925 2993
rect 2922 2943 2933 2946
rect 2890 2796 2893 2826
rect 2898 2813 2901 2943
rect 2906 2933 2925 2936
rect 2930 2926 2933 2943
rect 2890 2793 2901 2796
rect 2882 2783 2893 2786
rect 2866 2713 2877 2716
rect 2866 2666 2869 2713
rect 2866 2663 2877 2666
rect 2834 2643 2845 2646
rect 2874 2643 2877 2663
rect 2842 2616 2845 2643
rect 2834 2613 2845 2616
rect 2858 2623 2877 2626
rect 2858 2613 2861 2623
rect 2834 2536 2837 2613
rect 2850 2593 2853 2606
rect 2810 2473 2813 2536
rect 2834 2533 2845 2536
rect 2786 2423 2805 2426
rect 2786 2403 2789 2423
rect 2810 2416 2813 2426
rect 2794 2413 2813 2416
rect 2786 2383 2789 2396
rect 2794 2373 2797 2406
rect 2786 2333 2789 2346
rect 2786 2253 2789 2316
rect 2802 2306 2805 2406
rect 2810 2323 2813 2406
rect 2818 2396 2821 2496
rect 2826 2433 2829 2506
rect 2834 2503 2837 2516
rect 2826 2413 2829 2426
rect 2818 2393 2825 2396
rect 2822 2326 2825 2393
rect 2834 2363 2837 2476
rect 2818 2323 2825 2326
rect 2802 2303 2809 2306
rect 2762 2146 2765 2206
rect 2770 2186 2773 2216
rect 2770 2183 2781 2186
rect 2754 2143 2765 2146
rect 2754 2116 2757 2143
rect 2746 2113 2757 2116
rect 2738 1933 2741 2046
rect 2746 1983 2749 2113
rect 2762 2026 2765 2136
rect 2770 2113 2773 2146
rect 2778 2123 2781 2183
rect 2786 2173 2789 2226
rect 2794 2203 2797 2296
rect 2806 2226 2809 2303
rect 2802 2223 2809 2226
rect 2770 2086 2773 2106
rect 2770 2083 2781 2086
rect 2778 2036 2781 2083
rect 2754 2023 2765 2026
rect 2770 2033 2781 2036
rect 2754 1933 2757 1996
rect 2762 1953 2765 2006
rect 2698 1686 2701 1706
rect 2730 1703 2733 1816
rect 2738 1793 2741 1906
rect 2746 1776 2749 1926
rect 2754 1843 2757 1926
rect 2770 1903 2773 2033
rect 2786 2013 2797 2016
rect 2778 1876 2781 2006
rect 2770 1873 2781 1876
rect 2770 1856 2773 1873
rect 2786 1866 2789 1996
rect 2802 1913 2805 2223
rect 2810 2183 2813 2206
rect 2818 2166 2821 2323
rect 2826 2286 2829 2306
rect 2826 2283 2833 2286
rect 2830 2166 2833 2283
rect 2814 2163 2821 2166
rect 2826 2163 2833 2166
rect 2814 2076 2817 2163
rect 2814 2073 2821 2076
rect 2810 1996 2813 2056
rect 2818 2013 2821 2073
rect 2810 1993 2817 1996
rect 2826 1993 2829 2163
rect 2834 2113 2837 2146
rect 2814 1906 2817 1993
rect 2826 1923 2829 1946
rect 2794 1893 2797 1906
rect 2814 1903 2829 1906
rect 2834 1903 2837 2076
rect 2778 1863 2805 1866
rect 2770 1853 2789 1856
rect 2786 1836 2789 1853
rect 2802 1836 2805 1863
rect 2754 1833 2773 1836
rect 2754 1813 2757 1833
rect 2770 1816 2773 1833
rect 2778 1823 2781 1836
rect 2786 1833 2793 1836
rect 2802 1833 2813 1836
rect 2754 1783 2757 1806
rect 2762 1793 2765 1816
rect 2770 1813 2781 1816
rect 2742 1773 2749 1776
rect 2742 1716 2745 1773
rect 2754 1726 2757 1736
rect 2762 1733 2765 1746
rect 2754 1723 2761 1726
rect 2742 1713 2749 1716
rect 2698 1683 2709 1686
rect 2706 1636 2709 1683
rect 2698 1633 2709 1636
rect 2698 1613 2701 1633
rect 2706 1613 2717 1616
rect 2678 1603 2693 1606
rect 2690 1556 2693 1603
rect 2686 1553 2693 1556
rect 2674 1463 2677 1536
rect 2686 1496 2689 1553
rect 2706 1546 2709 1613
rect 2722 1573 2725 1616
rect 2698 1543 2709 1546
rect 2686 1493 2693 1496
rect 2666 1423 2677 1426
rect 2682 1423 2685 1476
rect 2650 1383 2657 1386
rect 2666 1386 2669 1416
rect 2674 1393 2677 1423
rect 2690 1413 2693 1493
rect 2698 1386 2701 1543
rect 2706 1513 2709 1536
rect 2666 1383 2701 1386
rect 2626 1173 2633 1176
rect 2618 1106 2621 1126
rect 2626 1113 2629 1173
rect 2634 1133 2637 1156
rect 2650 1136 2653 1383
rect 2658 1203 2661 1366
rect 2666 1253 2669 1336
rect 2674 1293 2677 1326
rect 2698 1323 2701 1383
rect 2690 1303 2693 1316
rect 2666 1243 2693 1246
rect 2666 1213 2669 1243
rect 2642 1133 2653 1136
rect 2642 1106 2645 1133
rect 2610 1096 2613 1106
rect 2618 1103 2645 1106
rect 2610 1093 2629 1096
rect 2594 1083 2605 1086
rect 2602 1013 2605 1083
rect 2594 1003 2605 1006
rect 2538 943 2581 946
rect 2538 933 2541 943
rect 2546 933 2557 936
rect 2530 796 2533 836
rect 2522 793 2533 796
rect 2506 713 2509 756
rect 2514 703 2517 736
rect 2498 603 2501 646
rect 2522 636 2525 793
rect 2530 646 2533 786
rect 2538 656 2541 816
rect 2546 803 2549 846
rect 2554 813 2557 916
rect 2562 913 2565 926
rect 2578 923 2581 943
rect 2586 933 2589 946
rect 2594 916 2597 996
rect 2602 923 2605 966
rect 2594 913 2605 916
rect 2602 896 2605 913
rect 2594 893 2605 896
rect 2562 803 2565 856
rect 2594 836 2597 893
rect 2594 833 2605 836
rect 2570 803 2573 816
rect 2578 803 2581 816
rect 2546 663 2549 736
rect 2554 716 2557 726
rect 2570 723 2573 736
rect 2554 713 2565 716
rect 2578 683 2581 736
rect 2586 723 2589 816
rect 2594 713 2597 746
rect 2538 653 2597 656
rect 2530 643 2549 646
rect 2506 613 2509 636
rect 2514 633 2525 636
rect 2514 543 2517 633
rect 2546 626 2549 643
rect 2546 623 2565 626
rect 2546 603 2549 623
rect 2530 526 2533 586
rect 2562 583 2565 616
rect 2570 556 2573 636
rect 2594 626 2597 653
rect 2602 643 2605 833
rect 2610 733 2613 1026
rect 2618 1013 2621 1026
rect 2626 1003 2629 1093
rect 2642 1043 2645 1103
rect 2634 1003 2637 1016
rect 2618 823 2621 976
rect 2642 926 2645 1006
rect 2650 1003 2653 1126
rect 2666 1073 2669 1206
rect 2674 1203 2677 1216
rect 2682 1133 2685 1236
rect 2690 1203 2693 1243
rect 2674 1106 2677 1126
rect 2690 1123 2693 1136
rect 2698 1126 2701 1216
rect 2706 1183 2709 1416
rect 2714 1356 2717 1556
rect 2722 1533 2725 1566
rect 2730 1443 2733 1676
rect 2738 1476 2741 1626
rect 2746 1486 2749 1713
rect 2758 1606 2761 1723
rect 2758 1603 2765 1606
rect 2754 1543 2757 1586
rect 2762 1543 2765 1603
rect 2754 1523 2757 1536
rect 2754 1493 2757 1506
rect 2746 1483 2757 1486
rect 2738 1473 2749 1476
rect 2722 1423 2733 1426
rect 2722 1366 2725 1406
rect 2730 1403 2733 1423
rect 2746 1403 2749 1473
rect 2754 1396 2757 1483
rect 2746 1393 2757 1396
rect 2722 1363 2733 1366
rect 2714 1353 2725 1356
rect 2722 1246 2725 1353
rect 2746 1346 2749 1393
rect 2738 1343 2749 1346
rect 2754 1343 2757 1366
rect 2738 1266 2741 1343
rect 2738 1263 2749 1266
rect 2722 1243 2733 1246
rect 2714 1173 2717 1206
rect 2698 1123 2709 1126
rect 2674 1103 2685 1106
rect 2658 986 2661 1066
rect 2666 1036 2669 1056
rect 2666 1033 2673 1036
rect 2626 923 2645 926
rect 2654 983 2661 986
rect 2654 926 2657 983
rect 2670 966 2673 1033
rect 2666 963 2673 966
rect 2654 923 2661 926
rect 2594 623 2605 626
rect 2546 553 2573 556
rect 2578 556 2581 616
rect 2578 553 2605 556
rect 2522 523 2533 526
rect 2498 513 2509 516
rect 2458 503 2469 506
rect 2522 466 2525 523
rect 2506 433 2509 466
rect 2522 463 2533 466
rect 2530 443 2533 463
rect 2410 403 2413 426
rect 2514 423 2517 436
rect 2538 413 2541 526
rect 2546 516 2549 553
rect 2554 543 2581 546
rect 2554 533 2557 543
rect 2562 533 2573 536
rect 2578 533 2581 543
rect 2578 523 2589 526
rect 2546 513 2557 516
rect 2594 513 2597 546
rect 2554 446 2557 513
rect 2594 483 2597 506
rect 2602 473 2605 553
rect 2610 523 2613 686
rect 2618 603 2621 736
rect 2626 583 2629 923
rect 2634 913 2645 916
rect 2658 906 2661 923
rect 2634 903 2661 906
rect 2634 686 2637 846
rect 2650 813 2653 876
rect 2642 723 2645 776
rect 2650 733 2653 806
rect 2650 686 2653 726
rect 2634 683 2653 686
rect 2634 643 2637 683
rect 2658 666 2661 856
rect 2666 673 2669 963
rect 2682 946 2685 1103
rect 2698 993 2701 1026
rect 2706 1016 2709 1106
rect 2714 1026 2717 1136
rect 2722 1133 2725 1186
rect 2722 1113 2725 1126
rect 2730 1123 2733 1243
rect 2738 1103 2741 1186
rect 2714 1023 2725 1026
rect 2706 1013 2717 1016
rect 2674 943 2685 946
rect 2698 943 2701 976
rect 2674 843 2677 943
rect 2706 933 2717 936
rect 2722 926 2725 1023
rect 2730 936 2733 1096
rect 2746 1086 2749 1263
rect 2754 1093 2757 1326
rect 2762 1226 2765 1516
rect 2770 1366 2773 1806
rect 2778 1723 2781 1813
rect 2790 1756 2793 1833
rect 2810 1766 2813 1833
rect 2810 1763 2821 1766
rect 2786 1753 2793 1756
rect 2786 1733 2789 1753
rect 2778 1686 2781 1716
rect 2778 1683 2789 1686
rect 2786 1613 2789 1683
rect 2794 1663 2797 1736
rect 2802 1723 2805 1746
rect 2810 1723 2813 1736
rect 2818 1723 2821 1763
rect 2778 1383 2781 1606
rect 2794 1573 2797 1616
rect 2802 1613 2805 1646
rect 2770 1363 2777 1366
rect 2774 1256 2777 1363
rect 2786 1333 2789 1546
rect 2794 1423 2797 1526
rect 2802 1483 2805 1606
rect 2826 1576 2829 1903
rect 2834 1813 2837 1896
rect 2842 1813 2845 2533
rect 2850 2523 2853 2586
rect 2858 2563 2861 2606
rect 2850 2103 2853 2476
rect 2858 2273 2861 2556
rect 2866 2403 2869 2536
rect 2874 2383 2877 2606
rect 2882 2343 2885 2726
rect 2890 2723 2893 2783
rect 2890 2623 2893 2676
rect 2898 2643 2901 2793
rect 2906 2636 2909 2926
rect 2914 2923 2933 2926
rect 2914 2803 2917 2923
rect 2922 2883 2925 2916
rect 2930 2813 2933 2856
rect 2938 2823 2941 2936
rect 2954 2923 2957 3113
rect 2962 2913 2965 3016
rect 2970 3003 2973 3026
rect 2970 2933 2973 2956
rect 2978 2923 2981 3156
rect 2994 2953 2997 3156
rect 3010 3123 3013 3196
rect 3042 3193 3045 3233
rect 3058 3203 3061 3346
rect 3066 3203 3069 3326
rect 3074 3323 3077 3353
rect 3074 3223 3077 3246
rect 3018 3123 3021 3136
rect 3026 3103 3029 3126
rect 3034 3066 3037 3136
rect 3030 3063 3037 3066
rect 3002 3013 3005 3026
rect 3018 3003 3021 3016
rect 3030 2966 3033 3063
rect 3042 3023 3045 3126
rect 3050 3116 3053 3136
rect 3050 3113 3061 3116
rect 3058 3046 3061 3113
rect 3050 3043 3061 3046
rect 3082 3046 3085 3336
rect 3090 3153 3093 3216
rect 3082 3043 3093 3046
rect 3050 3013 3053 3043
rect 3066 3023 3085 3026
rect 3066 3013 3069 3023
rect 3066 2983 3069 3006
rect 3074 2976 3077 3016
rect 3082 3003 3085 3023
rect 3090 2996 3093 3043
rect 3098 3013 3101 3216
rect 3106 3103 3109 3286
rect 3114 3213 3117 3346
rect 3122 3313 3125 3396
rect 3130 3343 3157 3346
rect 3130 3333 3133 3343
rect 3130 3283 3133 3326
rect 3122 3216 3125 3226
rect 3138 3216 3141 3336
rect 3154 3243 3157 3326
rect 3122 3213 3141 3216
rect 3122 3173 3125 3206
rect 3138 3203 3141 3213
rect 3162 3196 3165 3326
rect 3170 3223 3173 3336
rect 3194 3316 3197 3396
rect 3178 3313 3197 3316
rect 3146 3193 3165 3196
rect 3114 3143 3125 3146
rect 3114 3003 3117 3143
rect 3122 3086 3125 3136
rect 3130 3116 3133 3126
rect 3138 3123 3141 3166
rect 3146 3133 3149 3193
rect 3178 3156 3181 3313
rect 3194 3233 3197 3306
rect 3202 3243 3205 3376
rect 3218 3333 3229 3336
rect 3218 3323 3221 3333
rect 3234 3323 3237 3336
rect 3154 3153 3181 3156
rect 3130 3113 3149 3116
rect 3122 3083 3133 3086
rect 3138 3066 3141 3096
rect 3134 3063 3141 3066
rect 3122 3003 3125 3026
rect 3090 2993 3109 2996
rect 3042 2973 3077 2976
rect 3030 2963 3037 2966
rect 3034 2946 3037 2963
rect 3026 2943 3037 2946
rect 3002 2916 3005 2936
rect 3026 2923 3029 2943
rect 3002 2913 3021 2916
rect 2922 2803 2933 2806
rect 2922 2746 2925 2803
rect 2930 2783 2933 2796
rect 2938 2766 2941 2796
rect 2946 2773 2949 2906
rect 2962 2833 2989 2836
rect 2962 2813 2965 2833
rect 2954 2783 2957 2806
rect 2970 2783 2973 2806
rect 2978 2776 2981 2826
rect 2954 2773 2981 2776
rect 2938 2763 2949 2766
rect 2922 2743 2933 2746
rect 2914 2703 2917 2726
rect 2890 2553 2893 2616
rect 2890 2523 2893 2546
rect 2890 2503 2893 2516
rect 2890 2423 2893 2436
rect 2898 2376 2901 2636
rect 2906 2633 2917 2636
rect 2906 2583 2909 2626
rect 2914 2596 2917 2633
rect 2922 2603 2925 2736
rect 2930 2733 2933 2743
rect 2930 2723 2941 2726
rect 2946 2723 2949 2763
rect 2938 2703 2941 2716
rect 2954 2703 2957 2773
rect 2970 2723 2973 2756
rect 2930 2633 2933 2666
rect 2938 2606 2941 2626
rect 2938 2603 2949 2606
rect 2914 2593 2941 2596
rect 2906 2463 2909 2526
rect 2906 2403 2909 2416
rect 2914 2413 2917 2536
rect 2930 2533 2933 2546
rect 2922 2523 2933 2526
rect 2930 2423 2933 2436
rect 2930 2406 2933 2416
rect 2914 2403 2933 2406
rect 2938 2403 2941 2593
rect 2946 2443 2949 2556
rect 2954 2473 2957 2656
rect 2970 2613 2973 2716
rect 2978 2703 2981 2736
rect 2986 2693 2989 2833
rect 3002 2816 3005 2866
rect 2994 2813 3005 2816
rect 3010 2796 3013 2816
rect 3018 2803 3021 2913
rect 3034 2906 3037 2936
rect 3030 2903 3037 2906
rect 3030 2836 3033 2903
rect 3042 2863 3045 2973
rect 3058 2913 3069 2916
rect 3050 2893 3053 2906
rect 3058 2866 3061 2913
rect 3074 2903 3077 2936
rect 3082 2923 3085 2956
rect 3090 2896 3093 2946
rect 3054 2863 3061 2866
rect 3066 2893 3093 2896
rect 3030 2833 3037 2836
rect 3034 2813 3037 2833
rect 3042 2823 3045 2856
rect 3054 2806 3057 2863
rect 3026 2803 3037 2806
rect 3050 2803 3057 2806
rect 3026 2796 3029 2803
rect 3010 2793 3029 2796
rect 3050 2786 3053 2803
rect 2946 2413 2949 2436
rect 2946 2403 2957 2406
rect 2914 2383 2925 2386
rect 2930 2383 2933 2403
rect 2890 2373 2901 2376
rect 2866 2333 2885 2336
rect 2866 2283 2869 2333
rect 2858 2013 2861 2216
rect 2866 2213 2869 2246
rect 2874 2223 2877 2326
rect 2882 2323 2885 2333
rect 2890 2316 2893 2373
rect 2886 2313 2893 2316
rect 2886 2236 2889 2313
rect 2882 2233 2889 2236
rect 2882 2213 2885 2233
rect 2850 2003 2861 2006
rect 2850 1933 2853 1986
rect 2866 1976 2869 2206
rect 2890 2193 2893 2206
rect 2898 2173 2901 2366
rect 2906 2233 2909 2336
rect 2914 2223 2917 2356
rect 2874 2113 2877 2126
rect 2882 2123 2885 2146
rect 2898 2113 2901 2136
rect 2890 2073 2893 2106
rect 2906 2093 2909 2136
rect 2922 2106 2925 2383
rect 2962 2356 2965 2606
rect 2970 2593 2973 2606
rect 2986 2596 2989 2616
rect 2978 2593 2989 2596
rect 2978 2533 2981 2593
rect 2986 2583 2989 2593
rect 2970 2506 2973 2526
rect 2986 2523 2989 2566
rect 2994 2553 2997 2706
rect 2994 2533 2997 2546
rect 2970 2503 2981 2506
rect 2978 2436 2981 2503
rect 2994 2496 2997 2516
rect 2970 2433 2981 2436
rect 2990 2493 2997 2496
rect 2970 2416 2973 2433
rect 2970 2413 2981 2416
rect 2990 2376 2993 2493
rect 2990 2373 2997 2376
rect 2962 2353 2981 2356
rect 2930 2263 2933 2346
rect 2938 2343 2965 2346
rect 2938 2333 2941 2343
rect 2946 2333 2965 2336
rect 2938 2323 2957 2326
rect 2962 2246 2965 2333
rect 2930 2243 2965 2246
rect 2978 2246 2981 2353
rect 2994 2336 2997 2373
rect 3002 2353 3005 2726
rect 3010 2533 3013 2786
rect 3026 2783 3053 2786
rect 3018 2716 3021 2726
rect 3026 2723 3029 2783
rect 3050 2733 3053 2746
rect 3058 2733 3061 2776
rect 3066 2726 3069 2893
rect 3082 2816 3085 2846
rect 3090 2823 3093 2886
rect 3074 2766 3077 2816
rect 3082 2813 3093 2816
rect 3090 2783 3093 2806
rect 3098 2766 3101 2986
rect 3106 2793 3109 2993
rect 3114 2826 3117 2956
rect 3134 2936 3137 3063
rect 3134 2933 3141 2936
rect 3122 2903 3125 2926
rect 3138 2913 3141 2933
rect 3122 2833 3133 2836
rect 3114 2823 3125 2826
rect 3138 2823 3141 2856
rect 3074 2763 3085 2766
rect 3018 2713 3029 2716
rect 3018 2596 3021 2626
rect 3026 2603 3029 2713
rect 3050 2663 3053 2726
rect 3062 2723 3069 2726
rect 3074 2723 3077 2736
rect 3062 2666 3065 2723
rect 3082 2683 3085 2763
rect 3090 2763 3101 2766
rect 3090 2726 3093 2763
rect 3106 2733 3109 2756
rect 3090 2723 3101 2726
rect 3114 2723 3117 2776
rect 3058 2663 3065 2666
rect 3018 2593 3037 2596
rect 3010 2476 3013 2526
rect 3018 2493 3021 2566
rect 3026 2533 3029 2586
rect 3034 2503 3037 2593
rect 3042 2486 3045 2616
rect 3038 2483 3045 2486
rect 3010 2473 3029 2476
rect 3010 2373 3013 2416
rect 3018 2403 3021 2426
rect 3026 2413 3029 2473
rect 3026 2383 3029 2406
rect 3038 2346 3041 2483
rect 2990 2333 2997 2336
rect 3002 2333 3005 2346
rect 3038 2343 3045 2346
rect 2990 2266 2993 2333
rect 3002 2316 3005 2326
rect 3002 2313 3021 2316
rect 3026 2313 3029 2326
rect 3034 2303 3037 2326
rect 2990 2263 2997 2266
rect 2978 2243 2989 2246
rect 2930 2213 2933 2243
rect 2946 2213 2949 2236
rect 2962 2223 2965 2243
rect 2970 2203 2973 2216
rect 2938 2123 2941 2136
rect 2914 2086 2917 2106
rect 2922 2103 2933 2106
rect 2874 1996 2877 2026
rect 2882 2023 2893 2026
rect 2882 2003 2885 2016
rect 2890 1996 2893 2006
rect 2874 1993 2893 1996
rect 2850 1893 2853 1916
rect 2858 1906 2861 1976
rect 2866 1973 2873 1976
rect 2870 1916 2873 1973
rect 2882 1923 2885 1946
rect 2870 1913 2885 1916
rect 2898 1913 2901 2086
rect 2914 2083 2921 2086
rect 2906 2003 2909 2066
rect 2918 1996 2921 2083
rect 2914 1993 2921 1996
rect 2914 1973 2917 1993
rect 2930 1976 2933 2103
rect 2922 1973 2933 1976
rect 2946 1976 2949 2176
rect 2954 2103 2957 2126
rect 2962 2123 2965 2156
rect 2978 2123 2981 2226
rect 2986 2116 2989 2243
rect 2994 2133 2997 2263
rect 3002 2146 3005 2266
rect 3034 2256 3037 2276
rect 3026 2253 3037 2256
rect 3010 2213 3013 2236
rect 3026 2186 3029 2253
rect 3042 2193 3045 2343
rect 3050 2206 3053 2656
rect 3058 2223 3061 2663
rect 3066 2513 3069 2646
rect 3082 2613 3085 2646
rect 3074 2586 3077 2606
rect 3074 2583 3081 2586
rect 3078 2506 3081 2583
rect 3090 2566 3093 2716
rect 3098 2706 3101 2723
rect 3122 2716 3125 2823
rect 3146 2816 3149 3046
rect 3138 2813 3149 2816
rect 3130 2723 3133 2736
rect 3138 2723 3141 2813
rect 3146 2773 3149 2806
rect 3146 2723 3149 2736
rect 3154 2726 3157 3153
rect 3162 3126 3165 3146
rect 3162 3123 3173 3126
rect 3170 3046 3173 3123
rect 3186 3063 3189 3226
rect 3194 3223 3205 3226
rect 3210 3223 3213 3236
rect 3162 3043 3173 3046
rect 3194 3043 3197 3216
rect 3202 3206 3205 3223
rect 3202 3203 3209 3206
rect 3218 3203 3221 3316
rect 3250 3286 3253 3316
rect 3242 3283 3253 3286
rect 3206 3086 3209 3203
rect 3206 3083 3213 3086
rect 3162 3013 3165 3043
rect 3170 2993 3173 3026
rect 3162 2733 3165 2986
rect 3202 2983 3205 3066
rect 3210 2986 3213 3083
rect 3218 3043 3221 3156
rect 3210 2983 3221 2986
rect 3178 2973 3213 2976
rect 3170 2916 3173 2956
rect 3178 2933 3181 2973
rect 3210 2943 3213 2973
rect 3170 2913 3177 2916
rect 3174 2846 3177 2913
rect 3170 2843 3177 2846
rect 3154 2723 3165 2726
rect 3114 2713 3125 2716
rect 3130 2713 3157 2716
rect 3098 2703 3105 2706
rect 3102 2636 3105 2703
rect 3098 2633 3105 2636
rect 3098 2613 3101 2633
rect 3114 2613 3117 2713
rect 3122 2623 3125 2646
rect 3098 2603 3109 2606
rect 3114 2603 3125 2606
rect 3090 2563 3109 2566
rect 3098 2533 3101 2556
rect 3074 2503 3081 2506
rect 3074 2443 3077 2503
rect 3066 2333 3069 2416
rect 3074 2333 3077 2426
rect 3082 2413 3085 2426
rect 3082 2333 3085 2406
rect 3090 2333 3093 2526
rect 3098 2483 3101 2526
rect 3106 2496 3109 2563
rect 3114 2516 3117 2603
rect 3130 2556 3133 2713
rect 3138 2613 3141 2706
rect 3154 2613 3157 2706
rect 3130 2553 3137 2556
rect 3122 2533 3125 2546
rect 3114 2513 3125 2516
rect 3106 2493 3113 2496
rect 3098 2376 3101 2456
rect 3110 2416 3113 2493
rect 3106 2413 3113 2416
rect 3106 2393 3109 2413
rect 3122 2396 3125 2513
rect 3134 2496 3137 2553
rect 3118 2393 3125 2396
rect 3130 2493 3137 2496
rect 3098 2373 3109 2376
rect 3066 2323 3077 2326
rect 3066 2303 3069 2323
rect 3050 2203 3057 2206
rect 3026 2183 3045 2186
rect 3002 2143 3029 2146
rect 2970 2113 2989 2116
rect 2970 2046 2973 2113
rect 2994 2086 2997 2106
rect 2962 2043 2973 2046
rect 2986 2083 2997 2086
rect 2954 1983 2957 2016
rect 2946 1973 2957 1976
rect 2858 1903 2869 1906
rect 2866 1836 2869 1903
rect 2866 1833 2877 1836
rect 2850 1813 2861 1816
rect 2834 1793 2837 1806
rect 2842 1746 2845 1806
rect 2842 1743 2853 1746
rect 2834 1733 2845 1736
rect 2810 1573 2829 1576
rect 2810 1403 2813 1573
rect 2818 1513 2821 1566
rect 2826 1533 2829 1573
rect 2826 1486 2829 1506
rect 2822 1483 2829 1486
rect 2822 1416 2825 1483
rect 2834 1433 2837 1526
rect 2822 1413 2829 1416
rect 2826 1396 2829 1413
rect 2834 1403 2837 1426
rect 2786 1283 2789 1326
rect 2802 1323 2805 1336
rect 2810 1323 2813 1346
rect 2818 1333 2821 1396
rect 2826 1393 2837 1396
rect 2770 1253 2777 1256
rect 2770 1233 2773 1253
rect 2762 1223 2773 1226
rect 2786 1223 2789 1246
rect 2770 1166 2773 1223
rect 2778 1173 2781 1216
rect 2802 1186 2805 1316
rect 2818 1283 2821 1316
rect 2826 1213 2829 1386
rect 2786 1183 2805 1186
rect 2770 1163 2781 1166
rect 2762 1086 2765 1156
rect 2738 1083 2749 1086
rect 2754 1083 2765 1086
rect 2738 943 2741 1083
rect 2746 1013 2749 1026
rect 2746 973 2749 1006
rect 2730 933 2749 936
rect 2706 916 2709 926
rect 2722 923 2733 926
rect 2706 913 2725 916
rect 2730 906 2733 923
rect 2738 913 2741 926
rect 2722 903 2733 906
rect 2746 903 2749 933
rect 2674 743 2677 806
rect 2682 763 2685 836
rect 2698 813 2701 826
rect 2706 823 2717 826
rect 2674 703 2677 736
rect 2682 716 2685 726
rect 2690 723 2693 736
rect 2682 713 2701 716
rect 2642 663 2661 666
rect 2642 613 2645 663
rect 2658 623 2661 656
rect 2706 653 2709 823
rect 2714 673 2717 816
rect 2722 786 2725 903
rect 2730 853 2733 896
rect 2730 803 2733 826
rect 2738 803 2741 896
rect 2746 796 2749 896
rect 2754 813 2757 1083
rect 2762 1053 2765 1076
rect 2762 796 2765 1046
rect 2770 816 2773 1116
rect 2778 1023 2781 1163
rect 2786 1133 2789 1183
rect 2810 1156 2813 1206
rect 2834 1196 2837 1393
rect 2842 1293 2845 1733
rect 2850 1713 2853 1743
rect 2858 1696 2861 1806
rect 2854 1693 2861 1696
rect 2854 1586 2857 1693
rect 2866 1596 2869 1806
rect 2874 1706 2877 1833
rect 2882 1723 2885 1913
rect 2906 1903 2909 1956
rect 2890 1813 2893 1856
rect 2898 1803 2901 1816
rect 2914 1813 2917 1826
rect 2914 1743 2917 1766
rect 2874 1703 2881 1706
rect 2878 1646 2881 1703
rect 2874 1643 2881 1646
rect 2874 1613 2877 1643
rect 2890 1626 2893 1716
rect 2882 1623 2909 1626
rect 2882 1603 2885 1623
rect 2866 1593 2873 1596
rect 2854 1583 2861 1586
rect 2850 1523 2853 1566
rect 2858 1543 2861 1583
rect 2850 1493 2853 1516
rect 2858 1503 2861 1536
rect 2870 1496 2873 1593
rect 2890 1573 2893 1616
rect 2898 1606 2901 1616
rect 2898 1603 2909 1606
rect 2914 1593 2917 1606
rect 2922 1586 2925 1973
rect 2938 1933 2941 1956
rect 2954 1923 2957 1973
rect 2962 1916 2965 2043
rect 2986 2036 2989 2083
rect 2986 2033 2997 2036
rect 2970 2013 2973 2026
rect 2994 2013 2997 2033
rect 2994 1983 2997 1996
rect 2978 1923 2981 1976
rect 2994 1956 2997 1976
rect 2990 1953 2997 1956
rect 2946 1913 2965 1916
rect 2946 1846 2949 1913
rect 2946 1843 2953 1846
rect 2930 1793 2933 1826
rect 2938 1723 2941 1796
rect 2950 1786 2953 1843
rect 2962 1786 2965 1906
rect 2970 1853 2973 1916
rect 2990 1856 2993 1953
rect 2990 1853 2997 1856
rect 2970 1793 2973 1816
rect 2950 1783 2957 1786
rect 2962 1783 2973 1786
rect 2930 1603 2933 1616
rect 2946 1603 2949 1766
rect 2954 1703 2957 1783
rect 2962 1693 2965 1726
rect 2882 1516 2885 1566
rect 2914 1533 2917 1586
rect 2922 1583 2933 1586
rect 2930 1526 2933 1583
rect 2946 1566 2949 1586
rect 2898 1523 2909 1526
rect 2922 1523 2933 1526
rect 2942 1563 2949 1566
rect 2954 1563 2957 1626
rect 2898 1516 2901 1523
rect 2882 1513 2901 1516
rect 2866 1493 2873 1496
rect 2866 1426 2869 1493
rect 2850 1423 2869 1426
rect 2850 1386 2853 1423
rect 2858 1393 2861 1416
rect 2866 1413 2877 1416
rect 2882 1413 2885 1426
rect 2850 1383 2861 1386
rect 2794 1153 2813 1156
rect 2830 1193 2837 1196
rect 2778 1003 2781 1016
rect 2786 996 2789 1116
rect 2794 1003 2797 1153
rect 2786 993 2797 996
rect 2778 906 2781 946
rect 2786 913 2789 926
rect 2794 913 2797 993
rect 2802 933 2805 1126
rect 2818 1086 2821 1136
rect 2830 1096 2833 1193
rect 2830 1093 2837 1096
rect 2810 1083 2821 1086
rect 2810 1016 2813 1083
rect 2826 1023 2829 1076
rect 2810 1013 2821 1016
rect 2810 953 2813 1006
rect 2818 993 2821 1013
rect 2834 993 2837 1093
rect 2842 1006 2845 1236
rect 2850 1033 2853 1266
rect 2858 1226 2861 1383
rect 2874 1323 2877 1406
rect 2882 1313 2885 1406
rect 2890 1403 2893 1436
rect 2922 1426 2925 1523
rect 2942 1506 2945 1563
rect 2962 1556 2965 1606
rect 2954 1553 2965 1556
rect 2954 1533 2957 1553
rect 2970 1546 2973 1783
rect 2978 1733 2981 1836
rect 2986 1823 2989 1836
rect 2986 1706 2989 1816
rect 2994 1803 2997 1853
rect 2978 1703 2989 1706
rect 2978 1553 2981 1703
rect 2986 1636 2989 1656
rect 2986 1633 2993 1636
rect 2990 1546 2993 1633
rect 2962 1543 2973 1546
rect 2986 1543 2993 1546
rect 2962 1533 2965 1543
rect 2938 1503 2945 1506
rect 2938 1436 2941 1503
rect 2938 1433 2945 1436
rect 2914 1423 2925 1426
rect 2890 1333 2893 1396
rect 2898 1383 2901 1416
rect 2914 1316 2917 1423
rect 2930 1366 2933 1416
rect 2922 1363 2933 1366
rect 2922 1323 2925 1363
rect 2930 1353 2933 1363
rect 2942 1346 2945 1433
rect 2954 1396 2957 1526
rect 2978 1493 2981 1516
rect 2986 1503 2989 1543
rect 2994 1513 2997 1526
rect 2962 1413 2965 1466
rect 2970 1403 2973 1436
rect 2978 1396 2981 1406
rect 2954 1393 2981 1396
rect 2942 1343 2949 1346
rect 2930 1323 2941 1326
rect 2914 1313 2925 1316
rect 2858 1223 2877 1226
rect 2882 1223 2885 1266
rect 2922 1246 2925 1313
rect 2914 1243 2925 1246
rect 2946 1246 2949 1343
rect 2954 1333 2957 1346
rect 2946 1243 2953 1246
rect 2858 1203 2861 1223
rect 2858 1103 2861 1126
rect 2866 1036 2869 1216
rect 2874 1203 2877 1223
rect 2914 1156 2917 1243
rect 2914 1153 2925 1156
rect 2882 1123 2893 1126
rect 2898 1113 2901 1136
rect 2914 1123 2917 1136
rect 2906 1113 2917 1116
rect 2914 1093 2917 1113
rect 2866 1033 2877 1036
rect 2850 1013 2853 1026
rect 2866 1013 2869 1026
rect 2842 1003 2869 1006
rect 2778 903 2785 906
rect 2782 836 2785 903
rect 2782 833 2789 836
rect 2770 813 2781 816
rect 2738 793 2749 796
rect 2754 793 2765 796
rect 2770 793 2773 806
rect 2778 796 2781 813
rect 2786 803 2789 833
rect 2794 803 2797 856
rect 2802 843 2805 926
rect 2818 923 2821 936
rect 2778 793 2797 796
rect 2722 783 2729 786
rect 2726 716 2729 783
rect 2738 733 2741 793
rect 2754 776 2757 793
rect 2754 773 2765 776
rect 2754 726 2757 766
rect 2762 736 2765 773
rect 2762 733 2789 736
rect 2794 733 2797 793
rect 2754 723 2781 726
rect 2726 713 2733 716
rect 2754 713 2757 723
rect 2730 656 2733 713
rect 2762 706 2765 716
rect 2770 706 2773 716
rect 2778 713 2781 723
rect 2762 703 2773 706
rect 2722 653 2733 656
rect 2658 606 2661 616
rect 2682 613 2685 646
rect 2722 633 2725 653
rect 2770 646 2773 703
rect 2786 653 2789 733
rect 2802 716 2805 726
rect 2810 723 2813 916
rect 2826 913 2829 936
rect 2818 903 2845 906
rect 2818 833 2821 903
rect 2850 826 2853 916
rect 2834 786 2837 826
rect 2842 823 2853 826
rect 2842 793 2845 823
rect 2858 816 2861 956
rect 2866 823 2869 1003
rect 2874 973 2877 1033
rect 2882 926 2885 1026
rect 2874 923 2885 926
rect 2890 923 2893 1076
rect 2922 1036 2925 1153
rect 2930 1133 2933 1206
rect 2906 1033 2925 1036
rect 2898 993 2901 1006
rect 2906 953 2909 1033
rect 2930 1026 2933 1116
rect 2938 1083 2941 1236
rect 2950 1186 2953 1243
rect 2946 1183 2953 1186
rect 2914 1023 2941 1026
rect 2914 946 2917 1023
rect 2930 993 2933 1016
rect 2938 1013 2941 1023
rect 2898 943 2917 946
rect 2874 816 2877 916
rect 2882 906 2885 923
rect 2882 903 2889 906
rect 2886 836 2889 903
rect 2850 813 2861 816
rect 2866 813 2877 816
rect 2882 833 2889 836
rect 2850 786 2853 813
rect 2834 783 2853 786
rect 2826 723 2829 736
rect 2802 713 2829 716
rect 2770 643 2781 646
rect 2642 603 2661 606
rect 2634 536 2637 596
rect 2626 533 2637 536
rect 2642 523 2645 603
rect 2666 583 2669 606
rect 2690 603 2693 626
rect 2754 623 2773 626
rect 2754 613 2757 623
rect 2730 583 2733 596
rect 2754 593 2757 606
rect 2778 603 2781 643
rect 2786 613 2789 626
rect 2794 606 2797 616
rect 2786 603 2797 606
rect 2722 563 2757 566
rect 2650 506 2653 546
rect 2682 543 2685 556
rect 2658 533 2669 536
rect 2714 513 2717 526
rect 2642 503 2653 506
rect 2722 496 2725 563
rect 2730 523 2733 536
rect 2746 533 2749 556
rect 2754 536 2757 563
rect 2754 533 2765 536
rect 2770 516 2773 536
rect 2778 523 2781 546
rect 2786 533 2789 603
rect 2714 493 2725 496
rect 2730 513 2773 516
rect 2794 513 2797 536
rect 2802 523 2805 626
rect 2818 613 2821 706
rect 2826 676 2829 713
rect 2834 683 2837 736
rect 2842 676 2845 726
rect 2826 673 2845 676
rect 2826 603 2829 673
rect 2850 663 2853 726
rect 2858 706 2861 736
rect 2866 723 2869 813
rect 2882 766 2885 833
rect 2898 776 2901 943
rect 2922 936 2925 956
rect 2906 933 2925 936
rect 2906 913 2909 933
rect 2930 923 2933 986
rect 2938 973 2941 1006
rect 2946 976 2949 1183
rect 2962 1166 2965 1326
rect 2986 1323 2989 1416
rect 3002 1316 3005 2143
rect 3010 1946 3013 2126
rect 3018 2106 3021 2136
rect 3026 2123 3029 2143
rect 3018 2103 3025 2106
rect 3034 2103 3037 2146
rect 3022 1956 3025 2103
rect 3042 2096 3045 2183
rect 3034 2093 3045 2096
rect 3034 1976 3037 2093
rect 3054 2086 3057 2203
rect 3050 2083 3057 2086
rect 3050 2016 3053 2083
rect 3050 2013 3057 2016
rect 3042 1983 3045 2006
rect 3034 1973 3045 1976
rect 3022 1953 3029 1956
rect 3010 1943 3021 1946
rect 3010 1833 3013 1936
rect 3010 1803 3013 1816
rect 3018 1786 3021 1943
rect 3014 1783 3021 1786
rect 3014 1626 3017 1783
rect 3010 1623 3017 1626
rect 3010 1586 3013 1623
rect 3018 1593 3021 1616
rect 3010 1583 3021 1586
rect 3010 1513 3013 1526
rect 3018 1496 3021 1583
rect 3014 1493 3021 1496
rect 3014 1346 3017 1493
rect 3014 1343 3021 1346
rect 3018 1323 3021 1343
rect 2954 1163 2965 1166
rect 2954 1023 2957 1163
rect 2962 1123 2965 1156
rect 2970 1116 2973 1316
rect 3002 1313 3021 1316
rect 3010 1286 3013 1306
rect 3002 1283 3013 1286
rect 3002 1236 3005 1283
rect 3002 1233 3013 1236
rect 2978 1133 2981 1226
rect 3010 1213 3013 1233
rect 2986 1203 3005 1206
rect 2986 1123 2989 1186
rect 3010 1153 3013 1196
rect 3018 1146 3021 1313
rect 3002 1143 3021 1146
rect 2970 1113 2977 1116
rect 2954 996 2957 1016
rect 2962 1003 2965 1106
rect 2974 1016 2977 1113
rect 2974 1013 2981 1016
rect 2986 1013 2989 1026
rect 2970 996 2973 1006
rect 2954 993 2973 996
rect 2946 973 2957 976
rect 2938 913 2941 926
rect 2954 906 2957 973
rect 2978 933 2981 1013
rect 2994 1006 2997 1136
rect 2986 1003 2997 1006
rect 2986 983 2989 1003
rect 2986 923 2989 936
rect 2970 913 2981 916
rect 2914 813 2917 906
rect 2946 903 2957 906
rect 2906 803 2917 806
rect 2922 803 2925 836
rect 2938 796 2941 816
rect 2946 803 2949 903
rect 2994 896 2997 996
rect 2986 893 2997 896
rect 2930 793 2941 796
rect 2898 773 2905 776
rect 2882 763 2893 766
rect 2874 713 2877 736
rect 2858 703 2865 706
rect 2834 603 2837 656
rect 2862 646 2865 703
rect 2882 683 2885 726
rect 2862 643 2869 646
rect 2858 613 2861 636
rect 2866 613 2869 643
rect 2882 573 2885 676
rect 2890 633 2893 763
rect 2902 696 2905 773
rect 2914 703 2917 736
rect 2930 733 2933 793
rect 2902 693 2917 696
rect 2914 613 2917 693
rect 2922 663 2925 726
rect 2930 626 2933 726
rect 2922 623 2933 626
rect 2922 563 2925 623
rect 2930 593 2933 616
rect 2938 603 2941 726
rect 2946 723 2949 796
rect 2962 746 2965 846
rect 2986 826 2989 893
rect 2986 823 2997 826
rect 2970 796 2973 816
rect 2994 803 2997 823
rect 2970 793 2997 796
rect 2962 743 2969 746
rect 2946 673 2949 716
rect 2954 663 2957 736
rect 2966 676 2969 743
rect 2986 733 2989 746
rect 2978 713 2981 726
rect 2994 723 2997 793
rect 3002 733 3005 1143
rect 3026 1126 3029 1953
rect 3034 1893 3037 1936
rect 3042 1886 3045 1973
rect 3054 1936 3057 2013
rect 3066 2006 3069 2286
rect 3074 2206 3077 2316
rect 3082 2273 3085 2326
rect 3106 2306 3109 2373
rect 3098 2303 3109 2306
rect 3082 2223 3085 2256
rect 3090 2233 3093 2296
rect 3074 2203 3081 2206
rect 3078 2036 3081 2203
rect 3090 2183 3093 2226
rect 3098 2123 3101 2303
rect 3074 2033 3081 2036
rect 3074 2013 3077 2033
rect 3090 2016 3093 2116
rect 3106 2106 3109 2286
rect 3118 2226 3121 2393
rect 3130 2316 3133 2493
rect 3138 2323 3141 2466
rect 3146 2423 3149 2536
rect 3146 2343 3149 2416
rect 3154 2336 3157 2546
rect 3162 2523 3165 2723
rect 3170 2696 3173 2843
rect 3178 2806 3181 2826
rect 3186 2816 3189 2936
rect 3194 2913 3197 2936
rect 3202 2933 3213 2936
rect 3210 2903 3213 2926
rect 3218 2886 3221 2983
rect 3214 2883 3221 2886
rect 3214 2816 3217 2883
rect 3186 2813 3205 2816
rect 3214 2813 3221 2816
rect 3178 2803 3197 2806
rect 3178 2713 3181 2726
rect 3170 2693 3177 2696
rect 3174 2616 3177 2693
rect 3174 2613 3181 2616
rect 3162 2413 3165 2436
rect 3170 2406 3173 2606
rect 3178 2493 3181 2613
rect 3166 2403 3173 2406
rect 3166 2336 3169 2403
rect 3178 2393 3181 2416
rect 3146 2333 3157 2336
rect 3162 2333 3169 2336
rect 3130 2313 3141 2316
rect 3118 2223 3125 2226
rect 3130 2223 3133 2266
rect 3114 2183 3117 2206
rect 3082 2013 3093 2016
rect 3102 2103 3109 2106
rect 3082 2006 3085 2013
rect 3066 2003 3085 2006
rect 3038 1883 3045 1886
rect 3050 1933 3057 1936
rect 3038 1706 3041 1883
rect 3050 1813 3053 1933
rect 3082 1926 3085 2003
rect 3102 1956 3105 2103
rect 3114 2023 3117 2126
rect 3122 2016 3125 2223
rect 3138 2186 3141 2313
rect 3130 2183 3141 2186
rect 3130 2143 3133 2183
rect 3130 2033 3133 2076
rect 3090 1943 3093 1956
rect 3102 1953 3109 1956
rect 3058 1903 3061 1916
rect 3066 1813 3069 1926
rect 3078 1923 3085 1926
rect 3078 1836 3081 1923
rect 3090 1903 3093 1926
rect 3098 1856 3101 1936
rect 3106 1896 3109 1953
rect 3114 1913 3117 2016
rect 3122 2013 3129 2016
rect 3126 1906 3129 2013
rect 3122 1903 3129 1906
rect 3106 1893 3113 1896
rect 3090 1853 3101 1856
rect 3074 1833 3081 1836
rect 3050 1723 3053 1736
rect 3038 1703 3045 1706
rect 3042 1636 3045 1703
rect 3066 1643 3069 1806
rect 3074 1773 3077 1833
rect 3082 1723 3085 1826
rect 3090 1793 3093 1806
rect 3098 1756 3101 1816
rect 3110 1756 3113 1893
rect 3090 1753 3101 1756
rect 3106 1753 3113 1756
rect 3090 1656 3093 1753
rect 3098 1733 3101 1746
rect 3106 1686 3109 1753
rect 3082 1653 3093 1656
rect 3102 1683 3109 1686
rect 3034 1633 3045 1636
rect 3034 1593 3037 1633
rect 3058 1616 3061 1626
rect 3042 1613 3061 1616
rect 3066 1613 3069 1636
rect 3034 1513 3037 1586
rect 3042 1563 3045 1606
rect 3074 1603 3077 1616
rect 3074 1516 3077 1586
rect 3082 1533 3085 1653
rect 3066 1513 3077 1516
rect 3066 1466 3069 1513
rect 3066 1463 3077 1466
rect 3034 1203 3037 1446
rect 3058 1433 3061 1446
rect 3042 1293 3045 1426
rect 3050 1406 3053 1416
rect 3050 1403 3061 1406
rect 3066 1376 3069 1416
rect 3058 1373 3069 1376
rect 3050 1333 3053 1366
rect 3010 1103 3013 1126
rect 3022 1123 3029 1126
rect 3022 1046 3025 1123
rect 3034 1053 3037 1156
rect 3042 1113 3045 1256
rect 3058 1236 3061 1373
rect 3066 1313 3069 1366
rect 3050 1226 3053 1236
rect 3058 1233 3069 1236
rect 3050 1223 3061 1226
rect 3066 1216 3069 1233
rect 3050 1133 3053 1216
rect 3058 1213 3069 1216
rect 3022 1043 3029 1046
rect 3010 1013 3013 1036
rect 3026 996 3029 1043
rect 3050 1023 3053 1036
rect 3042 1003 3045 1016
rect 3026 993 3045 996
rect 3018 933 3021 946
rect 3010 913 3013 926
rect 3018 906 3021 926
rect 3026 923 3029 956
rect 3034 933 3037 976
rect 3042 923 3045 993
rect 3050 943 3053 986
rect 3018 903 3025 906
rect 3010 823 3013 886
rect 3022 836 3025 903
rect 3018 833 3025 836
rect 3018 813 3021 833
rect 3010 793 3013 806
rect 3034 796 3037 866
rect 3042 823 3045 886
rect 3026 793 3037 796
rect 3010 733 3013 756
rect 3026 706 3029 793
rect 3042 753 3045 816
rect 3058 756 3061 1213
rect 3066 1183 3069 1206
rect 3066 1113 3069 1126
rect 3066 973 3069 1016
rect 3066 923 3069 936
rect 3074 896 3077 1463
rect 3082 1186 3085 1526
rect 3090 1423 3093 1646
rect 3102 1636 3105 1683
rect 3102 1633 3109 1636
rect 3114 1633 3117 1676
rect 3098 1603 3101 1616
rect 3098 1523 3101 1596
rect 3106 1533 3109 1633
rect 3106 1513 3109 1526
rect 3114 1466 3117 1536
rect 3122 1526 3125 1903
rect 3138 1886 3141 2176
rect 3146 2006 3149 2333
rect 3154 2263 3157 2326
rect 3162 2256 3165 2333
rect 3170 2303 3173 2316
rect 3154 2253 3165 2256
rect 3154 2013 3157 2253
rect 3162 2223 3165 2246
rect 3170 2176 3173 2276
rect 3162 2173 3173 2176
rect 3162 2013 3165 2173
rect 3178 2166 3181 2366
rect 3170 2163 3181 2166
rect 3170 2083 3173 2163
rect 3178 2143 3181 2156
rect 3186 2126 3189 2766
rect 3194 2753 3197 2803
rect 3194 2716 3197 2736
rect 3202 2723 3205 2813
rect 3210 2783 3213 2796
rect 3218 2766 3221 2813
rect 3214 2763 3221 2766
rect 3214 2716 3217 2763
rect 3226 2726 3229 3246
rect 3234 3213 3237 3256
rect 3242 3223 3245 3283
rect 3258 3273 3261 3326
rect 3274 3233 3277 3366
rect 3282 3343 3309 3346
rect 3282 3333 3285 3343
rect 3290 3283 3293 3336
rect 3250 3223 3277 3226
rect 3250 3213 3253 3223
rect 3250 3203 3261 3206
rect 3234 3193 3261 3196
rect 3234 3133 3237 3193
rect 3242 3133 3245 3156
rect 3258 3133 3261 3193
rect 3234 3056 3237 3126
rect 3242 3123 3253 3126
rect 3242 3083 3245 3123
rect 3234 3053 3253 3056
rect 3234 3023 3237 3046
rect 3234 2923 3237 2966
rect 3242 2953 3245 3006
rect 3250 2943 3253 3053
rect 3234 2903 3237 2916
rect 3242 2873 3245 2936
rect 3258 2926 3261 3126
rect 3266 3103 3269 3206
rect 3274 3133 3277 3223
rect 3266 2996 3269 3026
rect 3274 3006 3277 3126
rect 3282 3023 3285 3256
rect 3290 3183 3293 3236
rect 3298 3213 3301 3226
rect 3306 3206 3309 3316
rect 3314 3296 3317 3336
rect 3322 3316 3325 3326
rect 3330 3323 3333 3386
rect 3346 3333 3373 3336
rect 3322 3313 3341 3316
rect 3314 3293 3325 3296
rect 3322 3236 3325 3293
rect 3346 3256 3349 3326
rect 3314 3233 3325 3236
rect 3338 3253 3349 3256
rect 3314 3213 3317 3233
rect 3322 3213 3333 3216
rect 3298 3203 3309 3206
rect 3322 3203 3325 3213
rect 3338 3206 3341 3253
rect 3354 3246 3357 3316
rect 3362 3293 3365 3316
rect 3370 3303 3373 3333
rect 3330 3203 3341 3206
rect 3346 3243 3357 3246
rect 3346 3203 3349 3243
rect 3354 3213 3357 3226
rect 3362 3223 3365 3266
rect 3370 3213 3373 3236
rect 3378 3206 3381 3326
rect 3386 3263 3389 3316
rect 3362 3203 3381 3206
rect 3290 3123 3293 3156
rect 3274 3003 3285 3006
rect 3266 2993 3281 2996
rect 3254 2923 3261 2926
rect 3254 2846 3257 2923
rect 3254 2843 3261 2846
rect 3250 2816 3253 2826
rect 3234 2813 3253 2816
rect 3234 2793 3237 2806
rect 3234 2743 3237 2776
rect 3258 2766 3261 2843
rect 3266 2813 3269 2976
rect 3278 2876 3281 2993
rect 3278 2873 3285 2876
rect 3250 2763 3261 2766
rect 3226 2723 3237 2726
rect 3194 2713 3205 2716
rect 3214 2713 3221 2716
rect 3194 2573 3197 2646
rect 3194 2513 3197 2536
rect 3202 2523 3205 2713
rect 3210 2603 3213 2626
rect 3218 2613 3221 2713
rect 3234 2656 3237 2723
rect 3250 2703 3253 2763
rect 3258 2733 3261 2756
rect 3258 2706 3261 2726
rect 3266 2723 3269 2746
rect 3274 2733 3277 2856
rect 3274 2706 3277 2716
rect 3258 2703 3277 2706
rect 3282 2696 3285 2873
rect 3290 2823 3293 3016
rect 3298 3003 3301 3203
rect 3306 3073 3309 3136
rect 3314 3093 3317 3126
rect 3322 3123 3325 3136
rect 3330 3123 3333 3203
rect 3362 3196 3365 3203
rect 3346 3193 3365 3196
rect 3346 3133 3349 3193
rect 3298 2923 3301 2946
rect 3298 2893 3301 2916
rect 3298 2816 3301 2876
rect 3306 2853 3309 3016
rect 3314 2933 3317 3016
rect 3322 2963 3325 3056
rect 3330 2956 3333 3026
rect 3338 2973 3341 3126
rect 3354 3123 3357 3146
rect 3362 3133 3365 3186
rect 3386 3173 3389 3216
rect 3394 3146 3397 3226
rect 3402 3203 3405 3216
rect 3378 3143 3397 3146
rect 3362 3123 3373 3126
rect 3378 3116 3381 3143
rect 3386 3133 3397 3136
rect 3418 3133 3421 3146
rect 3370 3113 3381 3116
rect 3354 3056 3357 3106
rect 3350 3053 3357 3056
rect 3350 2986 3353 3053
rect 3370 3046 3373 3113
rect 3394 3093 3397 3126
rect 3410 3086 3413 3126
rect 3434 3113 3437 3136
rect 3362 3043 3373 3046
rect 3402 3083 3413 3086
rect 3362 3003 3365 3043
rect 3386 3013 3389 3026
rect 3402 3023 3405 3083
rect 3370 3003 3381 3006
rect 3370 2986 3373 3003
rect 3394 2996 3397 3016
rect 3410 3013 3413 3026
rect 3418 3013 3421 3036
rect 3442 3026 3445 3126
rect 3378 2993 3397 2996
rect 3350 2983 3357 2986
rect 3370 2983 3381 2986
rect 3330 2953 3341 2956
rect 3322 2923 3325 2936
rect 3330 2933 3333 2946
rect 3338 2893 3341 2953
rect 3346 2886 3349 2966
rect 3354 2913 3357 2983
rect 3322 2883 3349 2886
rect 3306 2823 3309 2836
rect 3290 2813 3301 2816
rect 3314 2813 3317 2826
rect 3290 2803 3293 2813
rect 3298 2803 3309 2806
rect 3306 2733 3309 2803
rect 3226 2653 3237 2656
rect 3274 2693 3285 2696
rect 3210 2516 3213 2576
rect 3218 2533 3221 2546
rect 3226 2523 3229 2653
rect 3234 2613 3237 2636
rect 3242 2556 3245 2626
rect 3234 2553 3245 2556
rect 3234 2516 3237 2553
rect 3210 2513 3237 2516
rect 3210 2506 3213 2513
rect 3194 2503 3213 2506
rect 3194 2393 3197 2406
rect 3202 2403 3205 2426
rect 3194 2216 3197 2336
rect 3202 2333 3205 2376
rect 3202 2236 3205 2326
rect 3210 2246 3213 2503
rect 3218 2253 3221 2426
rect 3226 2333 3229 2496
rect 3226 2263 3229 2316
rect 3210 2243 3221 2246
rect 3202 2233 3213 2236
rect 3194 2213 3201 2216
rect 3198 2146 3201 2213
rect 3198 2143 3205 2146
rect 3182 2123 3189 2126
rect 3182 2056 3185 2123
rect 3182 2053 3189 2056
rect 3146 2003 3157 2006
rect 3134 1883 3141 1886
rect 3134 1816 3137 1883
rect 3134 1813 3141 1816
rect 3130 1783 3133 1796
rect 3130 1633 3133 1756
rect 3138 1616 3141 1813
rect 3146 1676 3149 1996
rect 3154 1686 3157 2003
rect 3162 1943 3165 1996
rect 3162 1803 3165 1896
rect 3170 1786 3173 2026
rect 3178 2013 3181 2036
rect 3178 1896 3181 2006
rect 3186 1906 3189 2053
rect 3194 1973 3197 2136
rect 3202 2023 3205 2143
rect 3194 1913 3197 1936
rect 3186 1903 3197 1906
rect 3202 1903 3205 1926
rect 3178 1893 3185 1896
rect 3182 1826 3185 1893
rect 3182 1823 3189 1826
rect 3166 1783 3173 1786
rect 3166 1726 3169 1783
rect 3178 1733 3181 1806
rect 3186 1796 3189 1823
rect 3194 1813 3197 1903
rect 3210 1803 3213 2233
rect 3186 1793 3213 1796
rect 3166 1723 3173 1726
rect 3154 1683 3165 1686
rect 3146 1673 3157 1676
rect 3130 1613 3141 1616
rect 3146 1613 3149 1626
rect 3130 1533 3141 1536
rect 3146 1533 3149 1546
rect 3122 1523 3133 1526
rect 3114 1463 3121 1466
rect 3090 1253 3093 1356
rect 3098 1263 3101 1436
rect 3106 1353 3109 1456
rect 3118 1346 3121 1463
rect 3114 1343 3121 1346
rect 3106 1273 3109 1316
rect 3082 1183 3101 1186
rect 3082 1133 3085 1176
rect 3098 1146 3101 1183
rect 3106 1153 3109 1206
rect 3082 1023 3085 1126
rect 3090 1123 3093 1146
rect 3098 1143 3105 1146
rect 3090 1013 3093 1036
rect 3070 893 3077 896
rect 3070 776 3073 893
rect 3082 783 3085 926
rect 3090 906 3093 936
rect 3102 926 3105 1143
rect 3102 923 3109 926
rect 3090 903 3097 906
rect 3094 826 3097 903
rect 3090 823 3097 826
rect 3090 806 3093 823
rect 3106 813 3109 923
rect 3114 843 3117 1343
rect 3122 1223 3125 1326
rect 3122 1183 3125 1216
rect 3122 1113 3125 1136
rect 3122 983 3125 996
rect 3122 813 3125 906
rect 3130 806 3133 1523
rect 3138 1453 3141 1533
rect 3146 1503 3149 1516
rect 3138 1413 3149 1416
rect 3154 1413 3157 1673
rect 3162 1453 3165 1683
rect 3170 1523 3173 1723
rect 3186 1706 3189 1776
rect 3202 1713 3205 1736
rect 3186 1703 3193 1706
rect 3178 1506 3181 1676
rect 3190 1636 3193 1703
rect 3186 1633 3193 1636
rect 3186 1573 3189 1633
rect 3194 1553 3197 1614
rect 3174 1503 3181 1506
rect 3162 1413 3165 1436
rect 3138 1306 3141 1356
rect 3146 1343 3149 1413
rect 3174 1406 3177 1503
rect 3154 1403 3165 1406
rect 3170 1403 3177 1406
rect 3154 1323 3157 1336
rect 3162 1323 3165 1386
rect 3138 1303 3149 1306
rect 3146 1226 3149 1303
rect 3138 1223 3149 1226
rect 3138 1166 3141 1223
rect 3162 1213 3165 1296
rect 3170 1283 3173 1403
rect 3178 1333 3181 1396
rect 3186 1346 3189 1526
rect 3202 1513 3205 1656
rect 3210 1576 3213 1793
rect 3218 1583 3221 2243
rect 3226 2183 3229 2196
rect 3226 2143 3229 2156
rect 3226 2026 3229 2136
rect 3234 2093 3237 2416
rect 3242 2266 3245 2546
rect 3250 2523 3253 2606
rect 3250 2283 3253 2516
rect 3258 2456 3261 2616
rect 3266 2533 3269 2556
rect 3266 2473 3269 2526
rect 3274 2466 3277 2693
rect 3290 2613 3293 2696
rect 3298 2606 3301 2716
rect 3306 2633 3309 2716
rect 3282 2603 3301 2606
rect 3282 2523 3285 2603
rect 3290 2513 3293 2546
rect 3298 2533 3301 2556
rect 3306 2523 3309 2606
rect 3306 2496 3309 2516
rect 3302 2493 3309 2496
rect 3274 2463 3285 2466
rect 3258 2453 3277 2456
rect 3258 2413 3261 2426
rect 3258 2323 3261 2356
rect 3242 2263 3249 2266
rect 3246 2156 3249 2263
rect 3258 2213 3261 2236
rect 3246 2153 3253 2156
rect 3242 2133 3245 2146
rect 3242 2103 3245 2126
rect 3226 2023 3233 2026
rect 3230 1956 3233 2023
rect 3242 2003 3245 2016
rect 3250 1996 3253 2153
rect 3258 2133 3261 2206
rect 3258 2103 3261 2116
rect 3242 1993 3253 1996
rect 3230 1953 3237 1956
rect 3226 1923 3229 1936
rect 3226 1903 3229 1916
rect 3226 1766 3229 1816
rect 3234 1813 3237 1953
rect 3242 1926 3245 1993
rect 3258 1986 3261 2096
rect 3250 1983 3261 1986
rect 3250 1933 3253 1983
rect 3242 1923 3249 1926
rect 3246 1806 3249 1923
rect 3234 1776 3237 1806
rect 3246 1803 3253 1806
rect 3258 1803 3261 1926
rect 3266 1906 3269 2446
rect 3274 2203 3277 2453
rect 3282 2376 3285 2463
rect 3302 2426 3305 2493
rect 3314 2453 3317 2806
rect 3322 2506 3325 2883
rect 3330 2823 3333 2836
rect 3330 2796 3333 2816
rect 3338 2813 3341 2826
rect 3330 2793 3341 2796
rect 3330 2613 3333 2786
rect 3338 2723 3341 2793
rect 3346 2773 3349 2856
rect 3362 2846 3365 2976
rect 3370 2933 3373 2966
rect 3378 2923 3381 2983
rect 3426 2966 3429 3026
rect 3394 2963 3429 2966
rect 3438 3023 3445 3026
rect 3370 2913 3381 2916
rect 3354 2843 3365 2846
rect 3354 2803 3357 2843
rect 3362 2823 3373 2826
rect 3362 2793 3365 2816
rect 3370 2803 3373 2823
rect 3354 2723 3357 2766
rect 3378 2763 3381 2913
rect 3386 2833 3389 2936
rect 3386 2803 3389 2816
rect 3362 2743 3389 2746
rect 3362 2733 3365 2743
rect 3370 2723 3373 2736
rect 3378 2723 3381 2736
rect 3386 2733 3389 2743
rect 3346 2683 3349 2716
rect 3338 2556 3341 2606
rect 3330 2553 3341 2556
rect 3346 2553 3349 2626
rect 3330 2533 3333 2553
rect 3354 2536 3357 2616
rect 3362 2613 3365 2706
rect 3386 2696 3389 2726
rect 3378 2693 3389 2696
rect 3370 2593 3373 2606
rect 3378 2563 3381 2693
rect 3394 2653 3397 2963
rect 3402 2933 3405 2956
rect 3438 2946 3441 3023
rect 3434 2943 3441 2946
rect 3402 2823 3405 2926
rect 3410 2906 3413 2926
rect 3410 2903 3421 2906
rect 3418 2856 3421 2903
rect 3410 2853 3421 2856
rect 3434 2856 3437 2943
rect 3434 2853 3445 2856
rect 3402 2783 3405 2816
rect 3410 2813 3413 2853
rect 3346 2533 3357 2536
rect 3386 2533 3389 2606
rect 3338 2513 3341 2526
rect 3322 2503 3329 2506
rect 3326 2436 3329 2503
rect 3346 2496 3349 2533
rect 3322 2433 3329 2436
rect 3342 2493 3349 2496
rect 3302 2423 3309 2426
rect 3290 2393 3293 2416
rect 3282 2373 3289 2376
rect 3286 2306 3289 2373
rect 3298 2333 3301 2406
rect 3282 2303 3289 2306
rect 3282 2183 3285 2303
rect 3290 2203 3293 2286
rect 3298 2203 3301 2216
rect 3274 2013 3277 2136
rect 3282 2113 3285 2126
rect 3282 1923 3285 2026
rect 3290 1933 3293 2196
rect 3298 2013 3301 2066
rect 3298 1993 3301 2006
rect 3266 1903 3277 1906
rect 3274 1836 3277 1903
rect 3266 1833 3277 1836
rect 3250 1786 3253 1803
rect 3250 1783 3257 1786
rect 3234 1773 3245 1776
rect 3226 1763 3237 1766
rect 3226 1593 3229 1716
rect 3234 1633 3237 1763
rect 3242 1733 3245 1773
rect 3254 1726 3257 1783
rect 3250 1723 3257 1726
rect 3242 1633 3245 1646
rect 3234 1613 3245 1616
rect 3210 1573 3221 1576
rect 3218 1506 3221 1573
rect 3234 1533 3237 1613
rect 3218 1503 3229 1506
rect 3202 1416 3205 1426
rect 3194 1413 3205 1416
rect 3194 1383 3197 1413
rect 3186 1343 3197 1346
rect 3178 1276 3181 1326
rect 3186 1323 3189 1336
rect 3170 1273 3181 1276
rect 3146 1203 3165 1206
rect 3162 1183 3165 1196
rect 3138 1163 3149 1166
rect 3146 1026 3149 1163
rect 3138 1023 3149 1026
rect 3138 896 3141 1023
rect 3146 993 3149 1006
rect 3146 923 3149 936
rect 3154 913 3157 996
rect 3138 893 3149 896
rect 3146 826 3149 893
rect 3090 803 3109 806
rect 3114 803 3133 806
rect 3138 823 3149 826
rect 3162 823 3165 926
rect 3170 906 3173 1273
rect 3178 1203 3181 1216
rect 3178 1093 3181 1116
rect 3186 1043 3189 1266
rect 3194 1123 3197 1343
rect 3210 1323 3213 1416
rect 3218 1306 3221 1486
rect 3214 1303 3221 1306
rect 3214 1236 3217 1303
rect 3202 1216 3205 1236
rect 3214 1233 3221 1236
rect 3202 1213 3209 1216
rect 3206 1126 3209 1213
rect 3218 1183 3221 1233
rect 3218 1133 3221 1166
rect 3202 1123 3209 1126
rect 3202 1103 3205 1123
rect 3186 1013 3189 1026
rect 3194 1013 3197 1036
rect 3210 1016 3213 1046
rect 3202 1013 3213 1016
rect 3178 923 3181 936
rect 3170 903 3177 906
rect 3070 773 3077 776
rect 3058 753 3069 756
rect 3042 713 3045 736
rect 3050 723 3053 736
rect 3066 723 3069 753
rect 3026 703 3045 706
rect 2962 673 2969 676
rect 2962 656 2965 673
rect 2954 653 2965 656
rect 2946 613 2949 636
rect 2954 553 2957 653
rect 2994 603 2997 636
rect 3010 563 3013 636
rect 2818 533 2829 536
rect 2866 533 2869 546
rect 2546 443 2557 446
rect 2418 396 2421 406
rect 2386 393 2421 396
rect 2378 373 2385 376
rect 2354 323 2373 326
rect 2382 316 2385 373
rect 2426 366 2429 396
rect 2394 333 2397 366
rect 2402 363 2429 366
rect 2402 336 2405 363
rect 2410 343 2421 346
rect 2402 333 2413 336
rect 2394 323 2405 326
rect 2298 293 2309 296
rect 2306 246 2309 293
rect 2298 243 2309 246
rect 2298 196 2301 243
rect 2322 203 2325 236
rect 2234 193 2269 196
rect 2242 103 2245 136
rect 2266 123 2269 193
rect 2274 163 2277 196
rect 2298 193 2309 196
rect 2306 146 2309 193
rect 2306 143 2325 146
rect 2338 143 2341 216
rect 2346 183 2349 206
rect 2322 123 2325 143
rect 2354 103 2357 306
rect 2362 213 2365 316
rect 2378 313 2385 316
rect 2378 256 2381 313
rect 2378 253 2397 256
rect 2378 223 2381 246
rect 2394 236 2397 253
rect 2394 233 2401 236
rect 2378 123 2381 206
rect 2386 143 2389 206
rect 2398 166 2401 233
rect 2410 213 2413 333
rect 2418 323 2421 343
rect 2426 333 2429 356
rect 2426 273 2429 326
rect 2434 213 2437 386
rect 2442 333 2445 346
rect 2450 336 2453 406
rect 2498 363 2501 406
rect 2546 366 2549 443
rect 2538 363 2549 366
rect 2450 333 2461 336
rect 2450 263 2453 326
rect 2490 253 2493 336
rect 2514 323 2517 346
rect 2522 313 2533 316
rect 2434 193 2437 206
rect 2450 203 2453 236
rect 2398 163 2437 166
rect 2434 123 2437 163
rect 2162 93 2197 96
rect 2442 83 2445 136
rect 2458 113 2461 216
rect 2490 193 2501 196
rect 2490 176 2493 193
rect 2474 173 2493 176
rect 2466 123 2469 166
rect 2474 133 2477 173
rect 2506 166 2509 216
rect 2514 193 2517 206
rect 2522 183 2525 313
rect 2538 283 2541 363
rect 2554 333 2557 416
rect 2562 403 2565 426
rect 2586 366 2589 406
rect 2594 403 2597 416
rect 2618 413 2621 436
rect 2714 406 2717 493
rect 2730 413 2733 513
rect 2746 486 2749 506
rect 2746 483 2757 486
rect 2754 436 2757 483
rect 2750 433 2757 436
rect 2642 386 2645 406
rect 2570 323 2573 366
rect 2582 363 2589 366
rect 2594 383 2645 386
rect 2582 316 2585 363
rect 2594 333 2597 383
rect 2642 373 2645 383
rect 2682 366 2685 406
rect 2714 403 2733 406
rect 2642 363 2685 366
rect 2594 323 2605 326
rect 2582 313 2589 316
rect 2618 313 2621 326
rect 2586 266 2589 313
rect 2578 263 2589 266
rect 2586 203 2589 216
rect 2610 213 2613 226
rect 2530 193 2541 196
rect 2482 163 2509 166
rect 2482 123 2485 163
rect 2618 143 2621 206
rect 2506 93 2509 116
rect 2546 96 2549 126
rect 2554 123 2557 136
rect 2586 106 2589 116
rect 2610 113 2621 116
rect 2626 106 2629 216
rect 2634 213 2637 306
rect 2642 253 2645 363
rect 2690 323 2693 346
rect 2730 333 2733 403
rect 2750 376 2753 433
rect 2746 373 2753 376
rect 2762 373 2765 416
rect 2802 413 2805 456
rect 2810 423 2853 426
rect 2810 413 2821 416
rect 2810 406 2813 413
rect 2794 403 2813 406
rect 2794 386 2797 403
rect 2790 383 2797 386
rect 2722 276 2725 326
rect 2714 273 2725 276
rect 2682 223 2693 226
rect 2682 213 2693 216
rect 2634 163 2637 206
rect 2682 196 2685 213
rect 2674 193 2685 196
rect 2674 146 2677 193
rect 2690 186 2693 206
rect 2698 193 2701 206
rect 2706 186 2709 266
rect 2714 233 2717 273
rect 2730 266 2733 326
rect 2746 303 2749 373
rect 2778 333 2781 346
rect 2722 263 2733 266
rect 2690 183 2709 186
rect 2714 176 2717 216
rect 2722 213 2725 263
rect 2674 143 2685 146
rect 2650 126 2653 136
rect 2642 123 2653 126
rect 2658 113 2661 126
rect 2682 123 2685 143
rect 2698 123 2701 176
rect 2706 173 2717 176
rect 2706 133 2709 173
rect 2722 133 2725 186
rect 2738 173 2741 206
rect 2746 193 2749 206
rect 2762 186 2765 326
rect 2790 306 2793 383
rect 2818 356 2821 406
rect 2802 353 2821 356
rect 2834 353 2837 416
rect 2850 403 2853 416
rect 2858 376 2861 526
rect 2874 523 2877 536
rect 2882 436 2885 526
rect 2906 513 2909 536
rect 2930 443 2933 536
rect 2954 523 2957 546
rect 3018 533 3021 626
rect 3042 623 3045 703
rect 3026 556 3029 616
rect 3074 603 3077 773
rect 3082 703 3085 726
rect 3090 713 3093 803
rect 3114 733 3117 803
rect 3114 696 3117 716
rect 3122 713 3125 726
rect 3106 693 3117 696
rect 3106 646 3109 693
rect 3106 643 3117 646
rect 3114 623 3117 643
rect 3130 623 3133 796
rect 3026 553 3037 556
rect 3010 446 3013 526
rect 3018 513 3021 526
rect 3034 476 3037 553
rect 3058 523 3061 596
rect 3082 533 3085 566
rect 3090 526 3093 596
rect 3122 583 3125 596
rect 3130 593 3133 616
rect 3138 603 3141 823
rect 3174 816 3177 903
rect 3186 893 3189 926
rect 3202 836 3205 1013
rect 3210 983 3213 1006
rect 3218 963 3221 1116
rect 3226 993 3229 1503
rect 3234 1413 3237 1526
rect 3242 1413 3245 1596
rect 3250 1516 3253 1723
rect 3266 1666 3269 1833
rect 3298 1823 3301 1886
rect 3258 1663 3269 1666
rect 3258 1573 3261 1663
rect 3266 1613 3269 1626
rect 3258 1523 3261 1566
rect 3250 1513 3261 1516
rect 3234 1323 3237 1396
rect 3242 1383 3245 1406
rect 3250 1366 3253 1456
rect 3246 1363 3253 1366
rect 3234 1223 3237 1276
rect 3246 1266 3249 1363
rect 3246 1263 3253 1266
rect 3234 973 3237 1206
rect 3242 943 3245 1246
rect 3250 1176 3253 1263
rect 3258 1196 3261 1513
rect 3266 1503 3269 1536
rect 3274 1493 3277 1816
rect 3282 1733 3285 1806
rect 3282 1703 3285 1716
rect 3290 1693 3293 1816
rect 3298 1713 3301 1726
rect 3282 1623 3285 1686
rect 3282 1533 3285 1616
rect 3282 1483 3285 1516
rect 3290 1466 3293 1606
rect 3298 1603 3301 1626
rect 3306 1586 3309 2423
rect 3314 2383 3317 2426
rect 3322 2366 3325 2433
rect 3342 2416 3345 2493
rect 3330 2373 3333 2416
rect 3338 2413 3345 2416
rect 3338 2396 3341 2413
rect 3354 2406 3357 2526
rect 3370 2413 3373 2526
rect 3346 2403 3357 2406
rect 3338 2393 3357 2396
rect 3362 2393 3365 2406
rect 3322 2363 3333 2366
rect 3314 2323 3317 2346
rect 3314 2293 3317 2316
rect 3314 2213 3317 2236
rect 3322 2213 3325 2336
rect 3330 2313 3333 2363
rect 3338 2333 3341 2346
rect 3338 2293 3341 2316
rect 3314 2183 3317 2206
rect 3322 2203 3333 2206
rect 3322 2123 3325 2203
rect 3338 2136 3341 2216
rect 3330 2133 3341 2136
rect 3322 2073 3325 2116
rect 3314 2013 3317 2036
rect 3338 2003 3341 2126
rect 3346 2123 3349 2216
rect 3346 2073 3349 2116
rect 3322 1933 3325 1956
rect 3338 1933 3341 1996
rect 3346 1936 3349 2016
rect 3354 1996 3357 2393
rect 3370 2216 3373 2406
rect 3386 2346 3389 2516
rect 3394 2356 3397 2636
rect 3402 2623 3405 2776
rect 3410 2736 3413 2756
rect 3418 2743 3421 2826
rect 3426 2753 3429 2836
rect 3442 2813 3445 2853
rect 3410 2733 3421 2736
rect 3418 2723 3421 2733
rect 3426 2716 3429 2736
rect 3422 2713 3429 2716
rect 3410 2623 3413 2686
rect 3422 2646 3425 2713
rect 3418 2643 3425 2646
rect 3402 2596 3405 2616
rect 3410 2603 3413 2616
rect 3418 2596 3421 2643
rect 3402 2593 3421 2596
rect 3418 2536 3421 2546
rect 3402 2533 3421 2536
rect 3402 2486 3405 2533
rect 3410 2513 3413 2526
rect 3418 2503 3421 2526
rect 3426 2513 3429 2626
rect 3402 2483 3413 2486
rect 3410 2426 3413 2483
rect 3410 2423 3421 2426
rect 3402 2363 3405 2416
rect 3418 2403 3421 2423
rect 3426 2403 3429 2426
rect 3394 2353 3429 2356
rect 3386 2343 3397 2346
rect 3370 2213 3381 2216
rect 3362 2003 3365 2206
rect 3386 2203 3389 2326
rect 3394 2223 3397 2343
rect 3370 2106 3373 2126
rect 3370 2103 3377 2106
rect 3374 2036 3377 2103
rect 3370 2033 3377 2036
rect 3370 2013 3373 2033
rect 3354 1993 3373 1996
rect 3346 1933 3365 1936
rect 3314 1913 3317 1926
rect 3322 1903 3325 1926
rect 3338 1883 3341 1916
rect 3354 1906 3357 1926
rect 3350 1903 3357 1906
rect 3350 1836 3353 1903
rect 3314 1803 3317 1816
rect 3322 1783 3325 1816
rect 3330 1813 3333 1826
rect 3338 1816 3341 1836
rect 3350 1833 3357 1836
rect 3338 1813 3349 1816
rect 3354 1813 3357 1833
rect 3314 1703 3317 1756
rect 3314 1623 3317 1636
rect 3314 1593 3317 1616
rect 3322 1603 3325 1726
rect 3330 1603 3333 1806
rect 3346 1736 3349 1796
rect 3354 1783 3357 1806
rect 3346 1733 3353 1736
rect 3338 1663 3341 1726
rect 3350 1676 3353 1733
rect 3346 1673 3353 1676
rect 3346 1656 3349 1673
rect 3338 1653 3349 1656
rect 3338 1613 3341 1653
rect 3362 1636 3365 1933
rect 3370 1823 3373 1993
rect 3346 1633 3365 1636
rect 3270 1463 3293 1466
rect 3302 1583 3309 1586
rect 3270 1356 3273 1463
rect 3302 1446 3305 1583
rect 3302 1443 3309 1446
rect 3290 1423 3301 1426
rect 3266 1353 3273 1356
rect 3266 1333 3269 1353
rect 3266 1213 3269 1326
rect 3274 1223 3277 1336
rect 3282 1243 3285 1416
rect 3290 1313 3293 1346
rect 3298 1323 3301 1336
rect 3290 1273 3301 1276
rect 3298 1233 3301 1273
rect 3258 1193 3269 1196
rect 3282 1193 3285 1216
rect 3250 1173 3257 1176
rect 3254 966 3257 1173
rect 3250 963 3257 966
rect 3210 913 3221 916
rect 3170 813 3177 816
rect 3186 833 3205 836
rect 3186 813 3189 833
rect 3194 823 3205 826
rect 3210 813 3213 826
rect 3218 813 3221 836
rect 3146 793 3149 806
rect 3146 573 3149 736
rect 3154 686 3157 716
rect 3162 703 3165 736
rect 3170 723 3173 813
rect 3178 723 3181 746
rect 3194 723 3197 736
rect 3154 683 3165 686
rect 3162 626 3165 683
rect 3154 623 3165 626
rect 3194 626 3197 716
rect 3202 693 3205 706
rect 3210 703 3213 716
rect 3194 623 3213 626
rect 3154 603 3157 623
rect 3186 613 3205 616
rect 3170 593 3181 596
rect 3186 563 3189 613
rect 3082 523 3093 526
rect 3026 473 3037 476
rect 3026 453 3029 473
rect 2962 443 3013 446
rect 2882 433 2933 436
rect 2866 393 2869 416
rect 2882 403 2885 433
rect 2922 413 2925 426
rect 2858 373 2909 376
rect 2802 313 2805 353
rect 2790 303 2797 306
rect 2770 276 2773 296
rect 2770 273 2781 276
rect 2778 226 2781 273
rect 2770 223 2781 226
rect 2770 203 2773 223
rect 2794 206 2797 303
rect 2818 253 2821 336
rect 2866 323 2869 346
rect 2898 243 2901 326
rect 2906 323 2909 373
rect 2922 343 2925 406
rect 2930 403 2933 433
rect 2962 426 2965 443
rect 2962 423 2973 426
rect 2802 233 2853 236
rect 2802 213 2805 233
rect 2786 203 2797 206
rect 2746 183 2765 186
rect 2730 133 2733 166
rect 2714 116 2717 126
rect 2722 123 2733 126
rect 2746 123 2749 183
rect 2786 146 2789 203
rect 2778 143 2789 146
rect 2714 113 2765 116
rect 2770 113 2773 126
rect 2586 103 2629 106
rect 2538 93 2549 96
rect 2778 73 2781 143
rect 2802 136 2805 206
rect 2850 203 2853 233
rect 2858 193 2861 226
rect 2898 213 2901 226
rect 2906 183 2909 206
rect 2914 156 2917 216
rect 2922 193 2925 336
rect 2874 153 2917 156
rect 2930 153 2933 396
rect 2938 376 2941 416
rect 2946 393 2949 406
rect 2954 383 2957 416
rect 2970 376 2973 423
rect 2986 386 2989 436
rect 3010 433 3013 443
rect 2994 403 2997 416
rect 3010 386 3013 406
rect 3034 393 3037 416
rect 3082 413 3085 523
rect 3098 506 3101 526
rect 3098 503 3109 506
rect 3106 446 3109 503
rect 3098 443 3109 446
rect 2986 383 3013 386
rect 2938 373 2945 376
rect 2942 266 2945 373
rect 2962 373 2973 376
rect 2962 333 2965 373
rect 2954 316 2957 326
rect 2962 323 2973 326
rect 2954 313 2973 316
rect 2938 263 2945 266
rect 2938 243 2941 263
rect 2946 213 2965 216
rect 2970 213 2973 313
rect 2986 296 2989 326
rect 2978 293 2989 296
rect 3010 253 3013 383
rect 3034 246 3037 326
rect 3050 253 3053 336
rect 3074 263 3077 326
rect 3034 243 3045 246
rect 2994 223 3005 226
rect 2970 176 2973 206
rect 2978 186 2981 206
rect 3018 203 3021 226
rect 2978 183 3005 186
rect 2970 173 2997 176
rect 2786 103 2789 136
rect 2794 133 2805 136
rect 2826 133 2869 136
rect 2826 113 2829 133
rect 2874 113 2877 153
rect 2930 53 2933 146
rect 2994 133 2997 173
rect 3002 163 3005 183
rect 3010 133 3013 196
rect 2946 113 2949 126
rect 3026 123 3029 216
rect 3042 213 3045 243
rect 3034 203 3045 206
rect 3034 133 3037 186
rect 3042 133 3045 196
rect 3042 113 3045 126
rect 3050 123 3053 156
rect 3066 143 3069 216
rect 3090 203 3093 416
rect 3098 413 3101 443
rect 3130 323 3133 536
rect 3146 496 3149 546
rect 3210 533 3213 623
rect 3218 603 3221 806
rect 3226 793 3229 936
rect 3242 893 3245 916
rect 3250 906 3253 963
rect 3266 946 3269 1193
rect 3282 1166 3285 1186
rect 3258 943 3269 946
rect 3278 1163 3285 1166
rect 3278 946 3281 1163
rect 3290 1136 3293 1226
rect 3298 1143 3301 1156
rect 3290 1133 3301 1136
rect 3298 1123 3301 1133
rect 3290 1013 3293 1096
rect 3298 1003 3301 1016
rect 3298 983 3301 996
rect 3306 976 3309 1443
rect 3314 1123 3317 1576
rect 3338 1533 3341 1606
rect 3330 1523 3341 1526
rect 3346 1516 3349 1633
rect 3370 1626 3373 1736
rect 3378 1733 3381 2016
rect 3386 1823 3389 2196
rect 3394 2163 3397 2216
rect 3402 2203 3405 2336
rect 3410 2283 3413 2326
rect 3418 2313 3421 2336
rect 3426 2306 3429 2353
rect 3418 2303 3429 2306
rect 3410 2203 3413 2216
rect 3418 2196 3421 2303
rect 3434 2286 3437 2766
rect 3442 2613 3445 2806
rect 3442 2486 3445 2556
rect 3450 2533 3453 3016
rect 3450 2503 3453 2526
rect 3442 2483 3449 2486
rect 3402 2193 3421 2196
rect 3430 2283 3437 2286
rect 3394 2023 3397 2036
rect 3394 1833 3397 1936
rect 3402 1803 3405 2193
rect 3410 2123 3413 2146
rect 3418 2133 3421 2156
rect 3430 2146 3433 2283
rect 3446 2276 3449 2483
rect 3426 2143 3433 2146
rect 3442 2273 3449 2276
rect 3418 2013 3421 2026
rect 3410 1933 3413 2006
rect 3410 1913 3413 1926
rect 3418 1846 3421 1936
rect 3426 1893 3429 2143
rect 3442 2076 3445 2273
rect 3438 2073 3445 2076
rect 3414 1843 3421 1846
rect 3386 1733 3389 1786
rect 3414 1756 3417 1843
rect 3414 1753 3421 1756
rect 3378 1683 3381 1726
rect 3394 1716 3397 1736
rect 3390 1713 3397 1716
rect 3354 1613 3357 1626
rect 3362 1623 3373 1626
rect 3362 1603 3365 1623
rect 3370 1603 3373 1616
rect 3378 1596 3381 1666
rect 3338 1513 3349 1516
rect 3354 1593 3381 1596
rect 3390 1596 3393 1713
rect 3402 1603 3405 1726
rect 3410 1723 3413 1736
rect 3418 1733 3421 1753
rect 3426 1696 3429 1836
rect 3438 1776 3441 2073
rect 3438 1773 3445 1776
rect 3434 1743 3437 1756
rect 3390 1593 3397 1596
rect 3322 1313 3325 1476
rect 3330 1403 3333 1446
rect 3338 1386 3341 1513
rect 3334 1383 3341 1386
rect 3334 1306 3337 1383
rect 3346 1323 3349 1496
rect 3334 1303 3341 1306
rect 3322 1223 3325 1246
rect 3330 1193 3333 1286
rect 3322 1143 3333 1146
rect 3314 1013 3317 1036
rect 3322 1013 3325 1136
rect 3330 1133 3333 1143
rect 3338 1123 3341 1303
rect 3346 1106 3349 1316
rect 3338 1103 3349 1106
rect 3338 1036 3341 1103
rect 3338 1033 3349 1036
rect 3346 1013 3349 1033
rect 3330 983 3333 1006
rect 3354 976 3357 1593
rect 3362 1473 3365 1526
rect 3362 1413 3365 1426
rect 3362 1383 3365 1396
rect 3370 1356 3373 1586
rect 3378 1503 3381 1536
rect 3386 1496 3389 1546
rect 3382 1493 3389 1496
rect 3382 1426 3385 1493
rect 3378 1423 3385 1426
rect 3378 1403 3381 1423
rect 3370 1353 3381 1356
rect 3362 1203 3365 1336
rect 3370 1236 3373 1346
rect 3378 1336 3381 1353
rect 3378 1333 3385 1336
rect 3382 1266 3385 1333
rect 3394 1323 3397 1593
rect 3402 1533 3405 1546
rect 3410 1533 3413 1696
rect 3422 1693 3429 1696
rect 3422 1636 3425 1693
rect 3422 1633 3429 1636
rect 3418 1533 3421 1616
rect 3402 1513 3405 1526
rect 3410 1503 3413 1526
rect 3426 1516 3429 1633
rect 3434 1623 3437 1686
rect 3422 1513 3429 1516
rect 3422 1436 3425 1513
rect 3422 1433 3429 1436
rect 3402 1413 3421 1416
rect 3426 1403 3429 1433
rect 3434 1423 3437 1606
rect 3402 1363 3405 1396
rect 3442 1356 3445 1773
rect 3402 1353 3445 1356
rect 3402 1313 3405 1353
rect 3410 1336 3413 1346
rect 3410 1333 3429 1336
rect 3410 1293 3413 1326
rect 3378 1263 3385 1266
rect 3378 1243 3381 1263
rect 3370 1233 3397 1236
rect 3362 1133 3365 1196
rect 3370 1163 3373 1226
rect 3378 1156 3381 1216
rect 3394 1166 3397 1233
rect 3394 1163 3405 1166
rect 3370 1153 3381 1156
rect 3370 1033 3373 1153
rect 3402 1146 3405 1163
rect 3378 1143 3405 1146
rect 3290 973 3309 976
rect 3330 973 3357 976
rect 3278 943 3285 946
rect 3258 913 3261 943
rect 3266 906 3269 926
rect 3250 903 3269 906
rect 3234 723 3237 736
rect 3242 723 3245 816
rect 3258 706 3261 903
rect 3282 886 3285 943
rect 3274 883 3285 886
rect 3274 773 3277 883
rect 3290 813 3293 973
rect 3298 923 3301 946
rect 3306 873 3309 926
rect 3330 923 3333 973
rect 3362 966 3365 1026
rect 3378 1006 3381 1143
rect 3386 1133 3397 1136
rect 3402 1133 3405 1143
rect 3394 1126 3397 1133
rect 3386 1106 3389 1126
rect 3394 1123 3405 1126
rect 3410 1106 3413 1236
rect 3426 1216 3429 1333
rect 3434 1326 3437 1353
rect 3450 1343 3453 2066
rect 3434 1323 3445 1326
rect 3426 1213 3433 1216
rect 3418 1153 3421 1206
rect 3430 1166 3433 1213
rect 3426 1163 3433 1166
rect 3426 1146 3429 1163
rect 3386 1103 3397 1106
rect 3394 1046 3397 1103
rect 3386 1043 3397 1046
rect 3406 1103 3413 1106
rect 3418 1143 3429 1146
rect 3386 1016 3389 1043
rect 3406 1036 3409 1103
rect 3406 1033 3413 1036
rect 3386 1013 3397 1016
rect 3338 926 3341 966
rect 3354 963 3365 966
rect 3370 1003 3389 1006
rect 3354 943 3357 963
rect 3370 946 3373 1003
rect 3394 946 3397 1013
rect 3402 993 3405 1016
rect 3410 963 3413 1033
rect 3418 1013 3421 1143
rect 3426 1096 3429 1116
rect 3426 1093 3433 1096
rect 3430 1036 3433 1093
rect 3426 1033 3433 1036
rect 3362 943 3373 946
rect 3390 943 3397 946
rect 3362 936 3365 943
rect 3354 933 3365 936
rect 3338 923 3357 926
rect 3362 903 3365 933
rect 3314 833 3349 836
rect 3370 833 3373 916
rect 3378 913 3381 926
rect 3390 846 3393 943
rect 3402 876 3405 936
rect 3402 873 3413 876
rect 3390 843 3397 846
rect 3282 793 3285 806
rect 3298 796 3301 826
rect 3290 793 3301 796
rect 3274 723 3285 726
rect 3250 703 3261 706
rect 3250 636 3253 703
rect 3250 633 3261 636
rect 3226 613 3229 626
rect 3258 613 3261 633
rect 3266 613 3269 716
rect 3274 613 3277 723
rect 3290 703 3293 793
rect 3298 736 3301 786
rect 3306 746 3309 816
rect 3314 783 3317 833
rect 3322 793 3325 826
rect 3330 813 3333 826
rect 3306 743 3317 746
rect 3298 733 3309 736
rect 3298 713 3301 726
rect 3282 633 3285 696
rect 3306 666 3309 733
rect 3298 663 3309 666
rect 3290 606 3293 626
rect 3250 603 3293 606
rect 3218 533 3221 546
rect 3242 533 3245 596
rect 3298 583 3301 663
rect 3306 613 3309 626
rect 3314 613 3317 743
rect 3330 713 3333 806
rect 3338 713 3341 726
rect 3346 706 3349 736
rect 3322 703 3349 706
rect 3370 703 3373 826
rect 3394 823 3397 843
rect 3410 823 3413 873
rect 3418 826 3421 936
rect 3426 893 3429 1033
rect 3442 1016 3445 1323
rect 3434 1013 3445 1016
rect 3434 913 3437 1013
rect 3442 976 3445 996
rect 3442 973 3449 976
rect 3446 906 3449 973
rect 3442 903 3449 906
rect 3418 823 3437 826
rect 3394 796 3397 816
rect 3386 793 3397 796
rect 3402 803 3421 806
rect 3386 746 3389 793
rect 3386 743 3397 746
rect 3378 723 3389 726
rect 3322 693 3325 703
rect 3378 633 3381 723
rect 3394 716 3397 743
rect 3386 713 3397 716
rect 3402 713 3405 803
rect 3410 713 3413 736
rect 3410 693 3413 706
rect 3378 606 3381 626
rect 3386 623 3413 626
rect 3418 623 3421 726
rect 3434 713 3437 823
rect 3442 813 3445 903
rect 3450 676 3453 696
rect 3442 673 3453 676
rect 3386 613 3389 623
rect 3394 613 3413 616
rect 3314 573 3317 606
rect 3362 593 3365 606
rect 3378 603 3389 606
rect 3154 516 3157 526
rect 3162 523 3173 526
rect 3154 513 3181 516
rect 3146 493 3157 496
rect 3154 426 3157 493
rect 3218 436 3221 526
rect 3250 513 3253 536
rect 3266 513 3269 546
rect 3306 533 3309 546
rect 3274 503 3277 526
rect 3210 433 3221 436
rect 3154 423 3165 426
rect 3146 413 3157 416
rect 3162 403 3165 423
rect 3170 403 3173 416
rect 3178 396 3181 426
rect 3186 403 3189 416
rect 3210 403 3213 433
rect 3170 393 3181 396
rect 3218 346 3221 426
rect 3226 416 3229 436
rect 3266 433 3293 436
rect 3250 423 3261 426
rect 3266 416 3269 433
rect 3226 413 3237 416
rect 3242 413 3269 416
rect 3290 413 3293 433
rect 3138 333 3141 346
rect 3218 343 3229 346
rect 3218 323 3221 336
rect 3226 293 3229 343
rect 3234 333 3237 413
rect 3258 403 3269 406
rect 3314 403 3317 436
rect 3322 383 3325 556
rect 3346 533 3349 566
rect 3354 533 3381 536
rect 3330 506 3333 526
rect 3378 516 3381 533
rect 3370 513 3381 516
rect 3386 513 3389 603
rect 3394 593 3397 613
rect 3410 593 3413 606
rect 3418 586 3421 606
rect 3394 583 3421 586
rect 3330 503 3341 506
rect 3338 436 3341 503
rect 3370 446 3373 513
rect 3370 443 3381 446
rect 3330 433 3341 436
rect 3330 413 3333 433
rect 3378 413 3381 443
rect 3394 433 3397 583
rect 3442 566 3445 673
rect 3442 563 3453 566
rect 3418 513 3421 526
rect 3402 423 3437 426
rect 3338 403 3357 406
rect 3402 403 3405 423
rect 3418 406 3421 416
rect 3434 413 3437 423
rect 3442 406 3445 546
rect 3282 333 3285 346
rect 3098 213 3101 246
rect 3138 213 3141 226
rect 3090 133 3093 186
rect 3098 133 3101 206
rect 3082 116 3085 126
rect 3106 123 3109 156
rect 3082 113 3133 116
rect 3138 113 3141 136
rect 3162 93 3165 256
rect 3186 123 3189 206
rect 3194 203 3197 236
rect 3242 213 3245 326
rect 3250 306 3253 326
rect 3250 303 3261 306
rect 3258 226 3261 303
rect 3306 293 3309 326
rect 3330 313 3333 336
rect 3338 323 3341 403
rect 3346 323 3349 346
rect 3354 296 3357 396
rect 3410 393 3413 406
rect 3418 403 3445 406
rect 3362 323 3365 386
rect 3386 333 3389 356
rect 3394 333 3413 336
rect 3410 326 3413 333
rect 3370 323 3389 326
rect 3410 323 3421 326
rect 3386 313 3413 316
rect 3354 293 3373 296
rect 3250 223 3261 226
rect 3250 123 3253 223
rect 3314 213 3317 226
rect 3274 173 3277 206
rect 3290 166 3293 206
rect 3370 196 3373 293
rect 3354 193 3373 196
rect 3354 176 3357 193
rect 3418 186 3421 323
rect 3426 313 3429 326
rect 3442 213 3445 403
rect 3450 353 3453 563
rect 3418 183 3445 186
rect 3266 163 3293 166
rect 3346 173 3357 176
rect 3266 93 3269 163
rect 3290 103 3293 126
rect 3346 123 3349 173
rect 3362 93 3365 136
rect 3386 113 3389 126
rect 3442 123 3445 183
rect 3462 37 3482 3403
rect 3486 13 3506 3427
<< metal3 >>
rect 1897 3432 2118 3437
rect 1593 3422 1854 3427
rect 1593 3417 1598 3422
rect 1297 3412 1598 3417
rect 1849 3417 1854 3422
rect 1897 3417 1902 3432
rect 2113 3417 2118 3432
rect 1849 3412 1902 3417
rect 1921 3412 2094 3417
rect 2113 3412 2142 3417
rect 2345 3412 2454 3417
rect 1921 3407 1926 3412
rect 1633 3402 1710 3407
rect 1745 3402 1926 3407
rect 2089 3407 2094 3412
rect 2345 3407 2350 3412
rect 2089 3402 2350 3407
rect 2449 3407 2454 3412
rect 2521 3412 2662 3417
rect 2449 3402 2478 3407
rect 1633 3397 1638 3402
rect 1609 3392 1638 3397
rect 1705 3397 1710 3402
rect 1961 3397 2070 3402
rect 2521 3397 2526 3412
rect 2657 3397 2662 3412
rect 2705 3412 2806 3417
rect 2705 3397 2710 3412
rect 1705 3392 1734 3397
rect 1937 3392 1966 3397
rect 2065 3392 2094 3397
rect 2361 3392 2526 3397
rect 2561 3392 2638 3397
rect 2657 3392 2710 3397
rect 2801 3397 2806 3412
rect 2961 3402 3102 3407
rect 2961 3397 2966 3402
rect 2801 3392 2830 3397
rect 2937 3392 2966 3397
rect 3097 3397 3102 3402
rect 3097 3392 3198 3397
rect 3217 3392 3294 3397
rect 1753 3387 1918 3392
rect 2561 3387 2566 3392
rect 1441 3382 1758 3387
rect 1913 3382 2110 3387
rect 2537 3382 2566 3387
rect 2633 3387 2638 3392
rect 2985 3387 3078 3392
rect 3217 3387 3222 3392
rect 2633 3382 2990 3387
rect 3073 3382 3222 3387
rect 3289 3387 3294 3392
rect 3289 3382 3334 3387
rect 2321 3377 2518 3382
rect 401 3372 678 3377
rect 1617 3372 2006 3377
rect 2025 3372 2054 3377
rect 2121 3372 2326 3377
rect 2513 3372 3206 3377
rect 401 3347 406 3372
rect 673 3357 678 3372
rect 1393 3367 1598 3372
rect 2049 3367 2126 3372
rect 729 3362 854 3367
rect 1265 3362 1350 3367
rect 1369 3362 1398 3367
rect 1593 3362 1638 3367
rect 1721 3362 1854 3367
rect 1929 3362 2014 3367
rect 2337 3362 3078 3367
rect 3217 3362 3278 3367
rect 1265 3357 1270 3362
rect 673 3352 702 3357
rect 841 3352 910 3357
rect 1241 3352 1270 3357
rect 1345 3357 1350 3362
rect 3073 3357 3222 3362
rect 1345 3352 1390 3357
rect 1449 3352 1958 3357
rect 2033 3352 2238 3357
rect 2257 3352 2438 3357
rect 2465 3352 3054 3357
rect 2033 3347 2038 3352
rect 281 3342 406 3347
rect 425 3342 478 3347
rect 561 3342 670 3347
rect 793 3342 1022 3347
rect 1281 3342 1478 3347
rect 1553 3342 1846 3347
rect 1857 3342 2038 3347
rect 2233 3347 2238 3352
rect 2233 3342 2294 3347
rect 1185 3337 1286 3342
rect 2057 3337 2214 3342
rect 2289 3337 2422 3342
rect 2465 3337 2470 3352
rect 2489 3342 2774 3347
rect 2857 3342 3118 3347
rect 3137 3342 3214 3347
rect 2769 3337 2862 3342
rect 3137 3337 3142 3342
rect 129 3332 222 3337
rect 1065 3332 1142 3337
rect 1185 3327 1190 3337
rect 1305 3332 2062 3337
rect 2209 3332 2278 3337
rect 2417 3332 2470 3337
rect 2537 3332 2558 3337
rect 2657 3332 2750 3337
rect 2881 3332 2982 3337
rect 3081 3332 3142 3337
rect 3209 3337 3214 3342
rect 3209 3332 3238 3337
rect 2537 3327 2542 3332
rect 905 3322 934 3327
rect 929 3317 934 3322
rect 993 3322 1054 3327
rect 993 3317 998 3322
rect 465 3312 886 3317
rect 929 3312 998 3317
rect 1049 3317 1054 3322
rect 1113 3322 1190 3327
rect 1217 3322 2542 3327
rect 2657 3322 2662 3332
rect 2881 3327 2886 3332
rect 2737 3322 2886 3327
rect 3065 3322 3222 3327
rect 1113 3317 1118 3322
rect 1217 3317 1222 3322
rect 2905 3317 3046 3322
rect 1049 3312 1118 3317
rect 1137 3312 1222 3317
rect 1241 3312 2430 3317
rect 2537 3312 2910 3317
rect 3041 3312 3358 3317
rect 265 3302 510 3307
rect 505 3297 510 3302
rect 649 3302 678 3307
rect 1185 3302 1214 3307
rect 1449 3302 1758 3307
rect 1985 3302 2182 3307
rect 2241 3302 2350 3307
rect 2417 3302 3374 3307
rect 649 3297 654 3302
rect 361 3292 390 3297
rect 505 3292 654 3297
rect 689 3292 814 3297
rect 1017 3292 1102 3297
rect 385 3277 390 3292
rect 689 3277 694 3292
rect 1209 3287 1214 3302
rect 1345 3297 1454 3302
rect 1777 3297 1878 3302
rect 1345 3287 1350 3297
rect 1473 3292 1510 3297
rect 1553 3292 1630 3297
rect 1721 3292 1782 3297
rect 1873 3292 2022 3297
rect 2129 3292 2166 3297
rect 2193 3292 2486 3297
rect 2633 3292 2918 3297
rect 2937 3292 2974 3297
rect 3081 3292 3366 3297
rect 2161 3287 2166 3292
rect 2505 3287 2614 3292
rect 2969 3287 3086 3292
rect 785 3282 838 3287
rect 1209 3282 1350 3287
rect 1369 3282 1398 3287
rect 1481 3282 1574 3287
rect 1641 3282 2118 3287
rect 2161 3282 2358 3287
rect 2393 3282 2510 3287
rect 2609 3282 2646 3287
rect 2817 3282 2950 3287
rect 3105 3282 3206 3287
rect 3217 3282 3294 3287
rect 2665 3277 2758 3282
rect 3201 3277 3206 3282
rect 385 3272 694 3277
rect 1705 3272 2670 3277
rect 2753 3272 2806 3277
rect 2897 3272 3174 3277
rect 3201 3272 3262 3277
rect 2801 3267 2902 3272
rect 1497 3262 1582 3267
rect 1601 3262 1742 3267
rect 1769 3262 1974 3267
rect 2081 3262 2198 3267
rect 2313 3262 2526 3267
rect 2673 3262 2742 3267
rect 2921 3262 3390 3267
rect 1497 3257 1502 3262
rect 1337 3252 1502 3257
rect 1577 3257 1582 3262
rect 2545 3257 2654 3262
rect 1577 3252 2550 3257
rect 2649 3252 2758 3257
rect 2825 3252 3286 3257
rect 985 3242 1070 3247
rect 1513 3242 1790 3247
rect 2137 3242 2982 3247
rect 985 3237 990 3242
rect 585 3232 990 3237
rect 1065 3237 1070 3242
rect 1849 3237 2118 3242
rect 2977 3237 2982 3242
rect 3049 3242 3078 3247
rect 3201 3242 3230 3247
rect 3049 3237 3054 3242
rect 1065 3232 1222 3237
rect 1361 3232 1638 3237
rect 1825 3232 1854 3237
rect 2113 3232 2918 3237
rect 2977 3232 3054 3237
rect 3209 3232 3294 3237
rect 3313 3232 3374 3237
rect 1721 3227 1806 3232
rect 3313 3227 3318 3232
rect 849 3222 878 3227
rect 1241 3222 1342 3227
rect 1505 3222 1726 3227
rect 1801 3222 2654 3227
rect 2705 3222 2750 3227
rect 2849 3222 2934 3227
rect 3185 3222 3246 3227
rect 3265 3222 3318 3227
rect 3353 3222 3398 3227
rect 1241 3217 1246 3222
rect 841 3212 894 3217
rect 953 3212 1102 3217
rect 1193 3212 1246 3217
rect 1337 3217 1342 3222
rect 2745 3217 2854 3222
rect 3265 3217 3270 3222
rect 1337 3212 1494 3217
rect 1737 3212 2398 3217
rect 2409 3212 2590 3217
rect 2625 3212 2726 3217
rect 2953 3212 3038 3217
rect 3097 3212 3270 3217
rect 1489 3207 1742 3212
rect 2953 3207 2958 3212
rect 377 3202 446 3207
rect 777 3202 974 3207
rect 1761 3202 2046 3207
rect 2057 3202 2182 3207
rect 2385 3202 2574 3207
rect 2673 3202 2822 3207
rect 2841 3202 2878 3207
rect 2905 3202 2958 3207
rect 3033 3207 3038 3212
rect 3033 3202 3062 3207
rect 3137 3202 3254 3207
rect 3265 3202 3406 3207
rect 377 3197 382 3202
rect 89 3192 342 3197
rect 353 3192 382 3197
rect 441 3197 446 3202
rect 2201 3197 2366 3202
rect 441 3192 470 3197
rect 897 3192 1046 3197
rect 1201 3192 1358 3197
rect 1393 3192 1454 3197
rect 1505 3192 1630 3197
rect 1649 3192 1742 3197
rect 1769 3192 1806 3197
rect 1817 3192 2206 3197
rect 2361 3192 2798 3197
rect 2969 3192 3150 3197
rect 337 3177 342 3192
rect 1649 3187 1654 3192
rect 481 3182 526 3187
rect 801 3182 902 3187
rect 913 3182 934 3187
rect 1001 3182 1110 3187
rect 1305 3182 1382 3187
rect 1425 3182 1654 3187
rect 1737 3187 1742 3192
rect 2793 3187 2974 3192
rect 1737 3182 2414 3187
rect 2457 3182 2662 3187
rect 3289 3182 3366 3187
rect 481 3177 486 3182
rect 913 3177 918 3182
rect 2681 3177 2774 3182
rect 337 3172 486 3177
rect 833 3172 918 3177
rect 937 3172 1190 3177
rect 1225 3172 1590 3177
rect 1665 3172 1942 3177
rect 2057 3172 2686 3177
rect 2769 3172 2934 3177
rect 2953 3172 3102 3177
rect 3121 3172 3278 3177
rect 3361 3172 3390 3177
rect 1185 3167 1190 3172
rect 1585 3167 1670 3172
rect 1937 3167 2062 3172
rect 2953 3167 2958 3172
rect 265 3162 318 3167
rect 729 3162 1174 3167
rect 1185 3162 1238 3167
rect 1401 3162 1566 3167
rect 1761 3162 1918 3167
rect 2081 3162 2502 3167
rect 2513 3162 2958 3167
rect 3097 3167 3102 3172
rect 3273 3167 3366 3172
rect 3097 3162 3142 3167
rect 1281 3157 1382 3162
rect 2497 3157 2502 3162
rect 569 3152 622 3157
rect 745 3152 798 3157
rect 809 3152 910 3157
rect 921 3152 998 3157
rect 1033 3152 1126 3157
rect 1201 3152 1286 3157
rect 1377 3152 1430 3157
rect 1441 3152 1550 3157
rect 1681 3152 1814 3157
rect 1937 3152 2038 3157
rect 2057 3152 2414 3157
rect 2497 3152 2982 3157
rect 2993 3152 3094 3157
rect 3217 3152 3246 3157
rect 3257 3152 3294 3157
rect 1937 3147 1942 3152
rect 193 3142 598 3147
rect 793 3142 894 3147
rect 929 3142 1078 3147
rect 1297 3142 1366 3147
rect 1473 3142 1502 3147
rect 1817 3142 1942 3147
rect 2033 3147 2038 3152
rect 2033 3142 2702 3147
rect 2761 3142 2942 3147
rect 3353 3142 3422 3147
rect 1473 3137 1478 3142
rect 3001 3137 3334 3142
rect 225 3132 270 3137
rect 1097 3132 1478 3137
rect 1569 3132 1798 3137
rect 1953 3132 2366 3137
rect 2401 3132 3006 3137
rect 3329 3132 3438 3137
rect 913 3127 998 3132
rect 1097 3127 1102 3132
rect 1569 3127 1574 3132
rect 1793 3127 1934 3132
rect 217 3122 342 3127
rect 337 3117 342 3122
rect 505 3122 534 3127
rect 889 3122 918 3127
rect 993 3122 1102 3127
rect 1449 3122 1574 3127
rect 1929 3122 2510 3127
rect 2529 3122 2598 3127
rect 2641 3122 2950 3127
rect 3017 3122 3366 3127
rect 505 3117 510 3122
rect 1209 3117 1366 3122
rect 1681 3117 1774 3122
rect 137 3112 174 3117
rect 257 3112 318 3117
rect 337 3112 510 3117
rect 769 3112 982 3117
rect 1073 3112 1214 3117
rect 1361 3112 1686 3117
rect 1769 3112 2246 3117
rect 2257 3112 2838 3117
rect 2921 3112 3342 3117
rect 2241 3107 2246 3112
rect 545 3102 638 3107
rect 913 3102 1214 3107
rect 1249 3102 1350 3107
rect 1449 3102 1502 3107
rect 1553 3102 2078 3107
rect 2241 3102 2566 3107
rect 2585 3102 2686 3107
rect 2737 3102 3030 3107
rect 3105 3102 3238 3107
rect 3265 3102 3358 3107
rect 1345 3097 1454 3102
rect 1297 3092 1326 3097
rect 1473 3087 1478 3102
rect 2097 3097 2222 3102
rect 1513 3092 2102 3097
rect 2217 3092 2542 3097
rect 2601 3092 2854 3097
rect 2953 3092 3142 3097
rect 3313 3092 3398 3097
rect 665 3082 1038 3087
rect 1121 3082 1454 3087
rect 1473 3082 1542 3087
rect 1649 3082 1790 3087
rect 1913 3082 2014 3087
rect 2049 3082 2158 3087
rect 2169 3082 2262 3087
rect 2297 3082 3110 3087
rect 3129 3082 3246 3087
rect 3105 3077 3110 3082
rect 305 3072 398 3077
rect 1113 3072 1142 3077
rect 1137 3067 1142 3072
rect 1481 3072 2550 3077
rect 2577 3072 2670 3077
rect 2681 3072 2926 3077
rect 3105 3072 3310 3077
rect 1481 3067 1486 3072
rect 2577 3067 2582 3072
rect 2921 3067 3094 3072
rect 785 3062 838 3067
rect 1137 3062 1486 3067
rect 1561 3062 1694 3067
rect 1721 3062 1766 3067
rect 1937 3062 2054 3067
rect 2161 3062 2350 3067
rect 2385 3062 2582 3067
rect 2609 3062 2902 3067
rect 3089 3062 3206 3067
rect 785 3057 790 3062
rect 1761 3057 1942 3062
rect 2049 3057 2166 3062
rect 585 3052 790 3057
rect 801 3052 830 3057
rect 881 3052 1062 3057
rect 1521 3052 1646 3057
rect 1665 3052 1742 3057
rect 265 3042 350 3047
rect 497 3042 814 3047
rect 265 3037 270 3042
rect 217 3032 270 3037
rect 345 3037 350 3042
rect 881 3037 886 3052
rect 345 3032 470 3037
rect 665 3032 750 3037
rect 833 3032 886 3037
rect 1057 3037 1062 3052
rect 1665 3047 1670 3052
rect 1737 3047 1742 3052
rect 1961 3052 2030 3057
rect 2185 3052 3326 3057
rect 1961 3047 1966 3052
rect 1505 3042 1534 3047
rect 1577 3042 1670 3047
rect 1713 3037 1718 3047
rect 1737 3042 1966 3047
rect 2097 3042 2430 3047
rect 2521 3042 2630 3047
rect 2649 3042 2678 3047
rect 2769 3042 2870 3047
rect 2913 3042 2942 3047
rect 3121 3042 3198 3047
rect 3217 3042 3238 3047
rect 2673 3037 2678 3042
rect 2937 3037 3126 3042
rect 1057 3032 1142 3037
rect 1201 3032 1310 3037
rect 1433 3032 1574 3037
rect 1689 3032 1718 3037
rect 1985 3032 2654 3037
rect 2673 3032 2886 3037
rect 489 3027 646 3032
rect 745 3027 838 3032
rect 1569 3027 1694 3032
rect 281 3022 334 3027
rect 441 3022 494 3027
rect 641 3022 710 3027
rect 873 3022 974 3027
rect 1025 3022 1046 3027
rect 1441 3022 1550 3027
rect 1785 3022 1830 3027
rect 1929 3022 1974 3027
rect 2081 3022 2254 3027
rect 2281 3022 2974 3027
rect 3001 3022 3046 3027
rect 3073 3022 3166 3027
rect 3265 3022 3286 3027
rect 3385 3022 3414 3027
rect 1025 3017 1030 3022
rect 1969 3017 1974 3022
rect 3073 3017 3078 3022
rect 129 3012 166 3017
rect 489 3012 846 3017
rect 1001 3012 1030 3017
rect 1041 3012 1150 3017
rect 1225 3012 1270 3017
rect 1497 3012 1734 3017
rect 1849 3012 1950 3017
rect 1969 3012 2326 3017
rect 2449 3012 2662 3017
rect 2745 3012 2814 3017
rect 2873 3012 3078 3017
rect 3097 3012 3310 3017
rect 3417 3012 3454 3017
rect 161 3007 166 3012
rect 841 3007 1006 3012
rect 161 3002 214 3007
rect 481 3002 678 3007
rect 1193 3002 1366 3007
rect 1385 3002 1478 3007
rect 1513 3002 1590 3007
rect 1689 3002 1942 3007
rect 2097 3002 2222 3007
rect 2313 3002 2398 3007
rect 2441 3002 2942 3007
rect 2961 3002 3022 3007
rect 3073 3002 3126 3007
rect 481 2997 486 3002
rect 1385 2997 1390 3002
rect 433 2992 486 2997
rect 497 2992 734 2997
rect 745 2992 894 2997
rect 937 2992 1070 2997
rect 1137 2992 1278 2997
rect 1345 2992 1390 2997
rect 1473 2997 1478 3002
rect 1985 2997 2078 3002
rect 1473 2992 1678 2997
rect 1953 2992 1990 2997
rect 2073 2992 3174 2997
rect 1673 2987 1958 2992
rect 457 2982 606 2987
rect 1049 2982 1302 2987
rect 1329 2982 1638 2987
rect 2001 2982 2502 2987
rect 2513 2982 2918 2987
rect 2977 2982 3102 2987
rect 3161 2982 3206 2987
rect 1297 2977 1302 2982
rect 2913 2977 2918 2982
rect 401 2972 614 2977
rect 625 2972 846 2977
rect 1089 2972 1206 2977
rect 1297 2972 1326 2977
rect 1353 2972 1390 2977
rect 1505 2972 1550 2977
rect 1585 2972 2174 2977
rect 2185 2972 2894 2977
rect 2913 2972 3270 2977
rect 3337 2972 3366 2977
rect 1297 2967 1302 2972
rect 377 2962 702 2967
rect 945 2962 998 2967
rect 1049 2962 1182 2967
rect 1297 2962 1414 2967
rect 1513 2962 1574 2967
rect 2153 2962 2310 2967
rect 2329 2962 2454 2967
rect 2473 2962 2526 2967
rect 2537 2962 3238 2967
rect 3321 2962 3374 2967
rect 1593 2957 1902 2962
rect 1953 2957 2134 2962
rect 129 2952 238 2957
rect 273 2952 318 2957
rect 465 2952 590 2957
rect 745 2952 902 2957
rect 1017 2952 1126 2957
rect 1273 2952 1406 2957
rect 1465 2952 1598 2957
rect 1897 2952 1958 2957
rect 2129 2952 2670 2957
rect 2769 2952 2974 2957
rect 2993 2952 3118 2957
rect 3169 2952 3246 2957
rect 3313 2952 3406 2957
rect 1121 2947 1126 2952
rect 2665 2947 2774 2952
rect 2993 2947 2998 2952
rect 441 2942 502 2947
rect 529 2942 598 2947
rect 617 2942 702 2947
rect 849 2942 918 2947
rect 993 2942 1070 2947
rect 1121 2942 1238 2947
rect 1257 2942 1886 2947
rect 1969 2942 2102 2947
rect 2121 2942 2222 2947
rect 2249 2942 2646 2947
rect 2793 2942 2998 2947
rect 3033 2942 3094 2947
rect 3185 2942 3254 2947
rect 3297 2942 3334 2947
rect 617 2937 622 2942
rect 217 2932 246 2937
rect 417 2932 550 2937
rect 569 2932 622 2937
rect 697 2937 702 2942
rect 1881 2937 1974 2942
rect 697 2932 726 2937
rect 737 2932 886 2937
rect 1105 2932 1206 2937
rect 1385 2932 1710 2937
rect 1833 2932 1862 2937
rect 1993 2932 3174 2937
rect 1201 2927 1390 2932
rect 1705 2927 1838 2932
rect 3185 2927 3190 2942
rect 3201 2932 3230 2937
rect 0 2922 430 2927
rect 521 2922 550 2927
rect 641 2922 710 2927
rect 729 2922 838 2927
rect 945 2922 1022 2927
rect 1105 2922 1182 2927
rect 1409 2922 1686 2927
rect 1913 2922 2062 2927
rect 2137 2922 2454 2927
rect 2529 2922 2622 2927
rect 2705 2922 2798 2927
rect 2849 2922 3190 2927
rect 3225 2927 3230 2932
rect 3297 2932 3326 2937
rect 3297 2927 3302 2932
rect 3225 2922 3302 2927
rect 545 2917 646 2922
rect 377 2907 454 2912
rect 705 2907 710 2922
rect 945 2917 950 2922
rect 921 2912 950 2917
rect 1017 2917 1022 2922
rect 1017 2912 1478 2917
rect 1537 2912 1766 2917
rect 1817 2912 2814 2917
rect 2849 2912 2870 2917
rect 2881 2912 2966 2917
rect 3065 2912 3198 2917
rect 3353 2912 3374 2917
rect 2881 2907 2886 2912
rect 233 2902 382 2907
rect 449 2902 478 2907
rect 521 2902 550 2907
rect 545 2897 550 2902
rect 609 2902 694 2907
rect 705 2902 1054 2907
rect 1481 2902 2054 2907
rect 2113 2902 2166 2907
rect 2177 2902 2726 2907
rect 2865 2902 2886 2907
rect 2945 2902 3078 2907
rect 3105 2902 3126 2907
rect 3209 2902 3238 2907
rect 609 2897 614 2902
rect 1169 2897 1294 2902
rect 2745 2897 2846 2902
rect 265 2892 294 2897
rect 289 2887 294 2892
rect 393 2892 422 2897
rect 545 2892 614 2897
rect 977 2892 1006 2897
rect 393 2887 398 2892
rect 289 2882 398 2887
rect 1001 2887 1006 2892
rect 1065 2892 1102 2897
rect 1145 2892 1174 2897
rect 1289 2892 1318 2897
rect 1521 2892 1622 2897
rect 1801 2892 2750 2897
rect 2841 2892 3198 2897
rect 3273 2892 3342 2897
rect 1065 2887 1070 2892
rect 1617 2887 1806 2892
rect 3193 2887 3278 2892
rect 1001 2882 1070 2887
rect 1177 2882 1598 2887
rect 1825 2882 1854 2887
rect 1905 2882 2086 2887
rect 2097 2882 2262 2887
rect 2345 2882 3094 2887
rect 633 2872 726 2877
rect 745 2872 766 2877
rect 929 2872 966 2877
rect 1169 2872 1270 2877
rect 1281 2872 1318 2877
rect 1537 2872 1934 2877
rect 2033 2872 2150 2877
rect 2353 2872 3302 2877
rect 633 2867 638 2872
rect 505 2862 638 2867
rect 721 2867 726 2872
rect 961 2867 966 2872
rect 1337 2867 1510 2872
rect 721 2862 862 2867
rect 961 2862 1342 2867
rect 1505 2862 1534 2867
rect 1793 2862 1822 2867
rect 1993 2862 2254 2867
rect 2377 2862 2982 2867
rect 3001 2862 3046 2867
rect 2977 2857 2982 2862
rect 401 2852 446 2857
rect 649 2852 822 2857
rect 1233 2852 1590 2857
rect 1689 2852 2590 2857
rect 2681 2852 2934 2857
rect 2977 2852 3278 2857
rect 3305 2852 3350 2857
rect 273 2842 366 2847
rect 401 2842 462 2847
rect 705 2842 982 2847
rect 1241 2842 1862 2847
rect 2025 2842 2070 2847
rect 2113 2842 2374 2847
rect 2401 2842 2542 2847
rect 2609 2842 2718 2847
rect 2753 2842 2774 2847
rect 2793 2842 3086 2847
rect 273 2837 278 2842
rect 249 2832 278 2837
rect 361 2837 366 2842
rect 1881 2837 2006 2842
rect 361 2832 462 2837
rect 529 2832 710 2837
rect 769 2832 806 2837
rect 913 2832 950 2837
rect 1209 2832 1246 2837
rect 1265 2832 1286 2837
rect 1353 2832 1542 2837
rect 1625 2832 1886 2837
rect 2001 2832 3334 2837
rect 3385 2832 3430 2837
rect 305 2822 350 2827
rect 497 2822 670 2827
rect 681 2822 790 2827
rect 1265 2817 1270 2832
rect 1457 2822 1494 2827
rect 1513 2822 2038 2827
rect 2049 2822 2166 2827
rect 2185 2822 2390 2827
rect 2409 2822 2526 2827
rect 2561 2822 2606 2827
rect 2689 2822 2734 2827
rect 2769 2822 2838 2827
rect 2889 2822 2942 2827
rect 2977 2822 3150 2827
rect 3265 2822 3294 2827
rect 2033 2817 2038 2822
rect 3145 2817 3270 2822
rect 3313 2817 3318 2827
rect 3337 2822 3406 2827
rect 153 2812 262 2817
rect 617 2812 838 2817
rect 1073 2812 1270 2817
rect 1569 2812 2014 2817
rect 2033 2812 2278 2817
rect 2289 2812 3006 2817
rect 3313 2812 3334 2817
rect 3385 2812 3414 2817
rect 457 2807 598 2812
rect 3057 2807 3126 2812
rect 129 2802 158 2807
rect 153 2797 158 2802
rect 217 2802 246 2807
rect 433 2802 462 2807
rect 593 2802 926 2807
rect 1233 2802 1270 2807
rect 1665 2802 1750 2807
rect 1801 2802 3062 2807
rect 3121 2802 3302 2807
rect 3313 2802 3358 2807
rect 217 2797 222 2802
rect 1553 2797 1646 2802
rect 153 2792 222 2797
rect 457 2792 582 2797
rect 689 2792 870 2797
rect 1105 2792 1342 2797
rect 1393 2792 1502 2797
rect 1529 2792 1558 2797
rect 1641 2792 2190 2797
rect 2297 2792 2486 2797
rect 2497 2792 2942 2797
rect 3073 2792 3110 2797
rect 3233 2792 3366 2797
rect 521 2782 590 2787
rect 633 2782 758 2787
rect 1065 2782 1110 2787
rect 1553 2782 1686 2787
rect 1857 2782 2422 2787
rect 2433 2782 2462 2787
rect 2489 2782 2654 2787
rect 2681 2782 2774 2787
rect 2809 2782 2862 2787
rect 2929 2782 2958 2787
rect 2969 2782 3014 2787
rect 3089 2782 3214 2787
rect 3329 2782 3406 2787
rect 1105 2777 1110 2782
rect 1265 2777 1558 2782
rect 1769 2777 1838 2782
rect 241 2772 390 2777
rect 561 2772 750 2777
rect 825 2772 934 2777
rect 1105 2772 1270 2777
rect 1577 2772 1774 2777
rect 1833 2772 2950 2777
rect 3057 2772 3118 2777
rect 3145 2772 3238 2777
rect 3345 2772 3406 2777
rect 241 2767 246 2772
rect 0 2762 246 2767
rect 385 2767 390 2772
rect 385 2762 886 2767
rect 1289 2762 1702 2767
rect 1697 2757 1702 2762
rect 1785 2762 2102 2767
rect 2177 2762 3358 2767
rect 3377 2762 3438 2767
rect 1785 2757 1790 2762
rect 497 2752 774 2757
rect 825 2752 894 2757
rect 1017 2752 1046 2757
rect 1065 2752 1086 2757
rect 1345 2752 1678 2757
rect 1697 2752 1790 2757
rect 1881 2752 2030 2757
rect 2121 2752 2462 2757
rect 2553 2752 2974 2757
rect 3105 2752 3198 2757
rect 3257 2752 3414 2757
rect 3425 2752 3446 2757
rect 161 2742 190 2747
rect 185 2737 190 2742
rect 257 2742 286 2747
rect 321 2742 374 2747
rect 481 2742 574 2747
rect 809 2742 838 2747
rect 1001 2742 1094 2747
rect 1185 2742 1270 2747
rect 1361 2742 1390 2747
rect 1617 2742 1646 2747
rect 1809 2742 2110 2747
rect 2233 2742 3270 2747
rect 3393 2742 3422 2747
rect 257 2737 262 2742
rect 569 2737 574 2742
rect 697 2737 814 2742
rect 1185 2737 1190 2742
rect 1385 2737 1622 2742
rect 2105 2737 2238 2742
rect 3393 2737 3398 2742
rect 185 2732 262 2737
rect 345 2732 550 2737
rect 569 2732 702 2737
rect 889 2732 1190 2737
rect 1729 2732 1950 2737
rect 1977 2732 2054 2737
rect 2257 2727 2262 2737
rect 2281 2732 2342 2737
rect 2449 2732 2566 2737
rect 2601 2732 2686 2737
rect 2801 2732 2822 2737
rect 2929 2732 2966 2737
rect 3049 2732 3078 2737
rect 3089 2732 3134 2737
rect 3161 2732 3198 2737
rect 3369 2732 3398 2737
rect 2801 2727 2806 2732
rect 2961 2727 2966 2732
rect 3089 2727 3094 2732
rect 281 2722 302 2727
rect 721 2722 766 2727
rect 873 2722 942 2727
rect 1433 2722 1550 2727
rect 1577 2722 1694 2727
rect 1713 2722 2262 2727
rect 2273 2722 2654 2727
rect 2689 2722 2726 2727
rect 2761 2722 2806 2727
rect 2841 2722 2942 2727
rect 2961 2722 2982 2727
rect 3001 2722 3094 2727
rect 3145 2722 3182 2727
rect 3337 2722 3382 2727
rect 1577 2717 1582 2722
rect 505 2712 550 2717
rect 1273 2712 1390 2717
rect 1553 2712 1582 2717
rect 1689 2717 1694 2722
rect 1689 2712 1782 2717
rect 1857 2712 1910 2717
rect 1993 2712 2078 2717
rect 2209 2712 2494 2717
rect 2649 2712 2654 2722
rect 3441 2717 3446 2752
rect 2825 2712 3070 2717
rect 3193 2712 3310 2717
rect 3385 2712 3446 2717
rect 1857 2707 1862 2712
rect 2673 2707 2774 2712
rect 3065 2707 3198 2712
rect 473 2702 526 2707
rect 753 2702 838 2707
rect 889 2702 934 2707
rect 1089 2702 1862 2707
rect 1881 2702 1918 2707
rect 1937 2702 2142 2707
rect 2593 2702 2678 2707
rect 2769 2702 2798 2707
rect 2809 2702 2854 2707
rect 2913 2702 2942 2707
rect 2977 2702 3046 2707
rect 3249 2702 3366 2707
rect 929 2697 934 2702
rect 2161 2697 2486 2702
rect 2593 2697 2598 2702
rect 3041 2697 3046 2702
rect 809 2692 846 2697
rect 929 2692 1046 2697
rect 1297 2692 1358 2697
rect 1689 2692 2166 2697
rect 2481 2692 2598 2697
rect 2609 2692 2990 2697
rect 3041 2692 3334 2697
rect 329 2682 454 2687
rect 329 2677 334 2682
rect 305 2672 334 2677
rect 449 2677 454 2682
rect 593 2682 734 2687
rect 1385 2682 1606 2687
rect 1945 2682 2294 2687
rect 2305 2682 2534 2687
rect 2561 2682 2694 2687
rect 2809 2682 3086 2687
rect 3153 2682 3182 2687
rect 593 2677 598 2682
rect 449 2672 598 2677
rect 729 2677 734 2682
rect 1641 2677 1830 2682
rect 3177 2677 3182 2682
rect 3321 2682 3414 2687
rect 3321 2677 3326 2682
rect 729 2672 798 2677
rect 1049 2672 1406 2677
rect 1617 2672 1646 2677
rect 1825 2672 1854 2677
rect 1985 2672 2894 2677
rect 2913 2672 3134 2677
rect 3177 2672 3326 2677
rect 1401 2667 1406 2672
rect 1513 2667 1622 2672
rect 2913 2667 2918 2672
rect 609 2662 702 2667
rect 1401 2662 1518 2667
rect 1657 2662 1742 2667
rect 1753 2662 1862 2667
rect 1881 2662 2278 2667
rect 2289 2662 2358 2667
rect 2465 2662 2606 2667
rect 2641 2662 2758 2667
rect 2793 2662 2918 2667
rect 2929 2662 3054 2667
rect 3073 2657 3214 2662
rect 297 2652 502 2657
rect 705 2652 886 2657
rect 921 2652 950 2657
rect 1057 2652 1182 2657
rect 1201 2652 1238 2657
rect 1561 2652 1630 2657
rect 1649 2652 2382 2657
rect 2433 2652 2478 2657
rect 2489 2652 2958 2657
rect 3049 2652 3078 2657
rect 3209 2652 3398 2657
rect 1057 2647 1062 2652
rect 529 2642 598 2647
rect 617 2642 662 2647
rect 913 2642 958 2647
rect 1033 2642 1062 2647
rect 1177 2647 1182 2652
rect 1561 2647 1566 2652
rect 1177 2642 1254 2647
rect 1273 2642 1382 2647
rect 1537 2642 1566 2647
rect 1625 2647 1630 2652
rect 1625 2642 2630 2647
rect 2873 2642 3070 2647
rect 3081 2642 3198 2647
rect 1273 2637 1278 2642
rect 297 2632 446 2637
rect 561 2632 782 2637
rect 833 2632 854 2637
rect 929 2632 1094 2637
rect 1129 2632 1278 2637
rect 1377 2637 1382 2642
rect 2721 2637 2806 2642
rect 1377 2632 1606 2637
rect 1721 2632 1782 2637
rect 1833 2632 1926 2637
rect 1961 2632 2022 2637
rect 2097 2632 2294 2637
rect 2345 2632 2726 2637
rect 2801 2632 2966 2637
rect 3185 2632 3238 2637
rect 3305 2632 3398 2637
rect 129 2622 198 2627
rect 217 2622 238 2627
rect 473 2622 550 2627
rect 633 2622 814 2627
rect 129 2617 134 2622
rect 0 2612 134 2617
rect 193 2617 198 2622
rect 545 2617 638 2622
rect 929 2617 934 2632
rect 1601 2627 1726 2632
rect 1777 2627 1782 2632
rect 2961 2627 3190 2632
rect 193 2612 510 2617
rect 657 2612 734 2617
rect 833 2612 934 2617
rect 961 2617 966 2627
rect 1169 2622 1366 2627
rect 1465 2622 1494 2627
rect 1777 2622 2078 2627
rect 2129 2622 2230 2627
rect 2337 2622 2390 2627
rect 2473 2622 2622 2627
rect 2737 2622 2790 2627
rect 3209 2622 3350 2627
rect 3401 2622 3430 2627
rect 1489 2617 1582 2622
rect 2809 2617 2942 2622
rect 961 2612 1054 2617
rect 1121 2612 1174 2617
rect 1185 2612 1326 2617
rect 1577 2612 1774 2617
rect 1865 2612 2814 2617
rect 2937 2612 3158 2617
rect 3353 2612 3446 2617
rect 833 2607 838 2612
rect 1169 2607 1174 2612
rect 1769 2607 1870 2612
rect 201 2602 246 2607
rect 457 2602 710 2607
rect 753 2602 838 2607
rect 857 2602 998 2607
rect 1169 2602 1558 2607
rect 1889 2602 2462 2607
rect 2577 2602 2694 2607
rect 2785 2602 2854 2607
rect 2873 2602 2926 2607
rect 3097 2602 3310 2607
rect 3385 2602 3414 2607
rect 145 2592 174 2597
rect 169 2587 174 2592
rect 241 2592 302 2597
rect 361 2592 414 2597
rect 425 2592 486 2597
rect 529 2592 558 2597
rect 641 2592 766 2597
rect 817 2592 854 2597
rect 865 2592 1134 2597
rect 1241 2592 1334 2597
rect 1489 2592 1542 2597
rect 1617 2592 1726 2597
rect 1825 2592 2254 2597
rect 2361 2592 3086 2597
rect 3345 2592 3374 2597
rect 241 2587 246 2592
rect 849 2587 854 2592
rect 1353 2587 1470 2592
rect 1617 2587 1622 2592
rect 169 2582 246 2587
rect 417 2582 470 2587
rect 625 2582 662 2587
rect 689 2582 774 2587
rect 849 2582 894 2587
rect 1049 2582 1134 2587
rect 1153 2582 1358 2587
rect 1465 2582 1622 2587
rect 1721 2587 1726 2592
rect 2249 2587 2366 2592
rect 3081 2587 3350 2592
rect 1721 2582 2022 2587
rect 2073 2582 2182 2587
rect 2193 2582 2230 2587
rect 2385 2582 2478 2587
rect 2545 2582 2718 2587
rect 2785 2582 2822 2587
rect 2849 2582 2910 2587
rect 2985 2582 3030 2587
rect 265 2572 326 2577
rect 457 2572 526 2577
rect 777 2572 798 2577
rect 985 2572 1094 2577
rect 577 2567 718 2572
rect 513 2562 582 2567
rect 713 2562 742 2567
rect 801 2562 838 2567
rect 1065 2562 1126 2567
rect 897 2557 1046 2562
rect 0 2552 278 2557
rect 273 2547 278 2552
rect 337 2552 902 2557
rect 1041 2552 1070 2557
rect 1081 2552 1110 2557
rect 337 2547 342 2552
rect 1081 2547 1086 2552
rect 1153 2547 1158 2582
rect 1169 2572 1382 2577
rect 1417 2572 1550 2577
rect 1633 2572 1662 2577
rect 1881 2572 2230 2577
rect 2281 2572 2406 2577
rect 2457 2572 3046 2577
rect 3081 2572 3174 2577
rect 3193 2572 3214 2577
rect 3233 2572 3358 2577
rect 1657 2567 1662 2572
rect 1793 2567 1886 2572
rect 3081 2567 3086 2572
rect 1241 2562 1278 2567
rect 1337 2562 1430 2567
rect 1657 2562 1798 2567
rect 1905 2562 2150 2567
rect 2185 2562 2222 2567
rect 2617 2562 2782 2567
rect 2857 2562 2990 2567
rect 3017 2562 3086 2567
rect 3169 2567 3174 2572
rect 3233 2567 3238 2572
rect 3169 2562 3238 2567
rect 3353 2567 3358 2572
rect 3353 2562 3382 2567
rect 2433 2557 2558 2562
rect 1369 2552 1518 2557
rect 1873 2552 2294 2557
rect 2305 2552 2366 2557
rect 2409 2552 2438 2557
rect 2553 2552 2582 2557
rect 2593 2552 2798 2557
rect 2857 2552 2894 2557
rect 2945 2552 2998 2557
rect 3097 2552 3334 2557
rect 3345 2552 3446 2557
rect 273 2542 342 2547
rect 417 2542 790 2547
rect 809 2542 862 2547
rect 945 2542 1046 2547
rect 1065 2542 1086 2547
rect 1089 2542 1158 2547
rect 1169 2542 1622 2547
rect 1817 2542 2174 2547
rect 2353 2542 2614 2547
rect 2721 2542 2774 2547
rect 2785 2542 2814 2547
rect 2889 2542 2998 2547
rect 857 2537 862 2542
rect 209 2532 254 2537
rect 505 2532 606 2537
rect 601 2527 606 2532
rect 665 2532 758 2537
rect 857 2532 990 2537
rect 665 2527 670 2532
rect 1089 2527 1094 2542
rect 1169 2537 1174 2542
rect 2193 2537 2334 2542
rect 2625 2537 2726 2542
rect 2785 2537 2790 2542
rect 3009 2537 3014 2547
rect 3121 2542 3158 2547
rect 3217 2542 3294 2547
rect 1137 2532 1174 2537
rect 1185 2532 1278 2537
rect 1809 2532 1854 2537
rect 1921 2532 2198 2537
rect 2329 2532 2518 2537
rect 2577 2532 2630 2537
rect 2745 2532 2790 2537
rect 2809 2532 3150 2537
rect 3313 2532 3390 2537
rect 1369 2527 1454 2532
rect 3177 2527 3318 2532
rect 3385 2527 3390 2532
rect 225 2522 246 2527
rect 537 2522 582 2527
rect 601 2522 670 2527
rect 1041 2522 1094 2527
rect 1113 2522 1374 2527
rect 1449 2522 1638 2527
rect 1817 2522 2038 2527
rect 2161 2522 2246 2527
rect 2305 2522 2574 2527
rect 2681 2522 2710 2527
rect 2769 2522 2854 2527
rect 2929 2522 3182 2527
rect 3385 2522 3414 2527
rect 225 2517 230 2522
rect 857 2517 958 2522
rect 137 2512 230 2517
rect 297 2512 358 2517
rect 833 2512 862 2517
rect 953 2512 982 2517
rect 1153 2512 1302 2517
rect 1297 2507 1302 2512
rect 1385 2512 1438 2517
rect 1745 2512 1806 2517
rect 2009 2512 2854 2517
rect 2993 2512 3070 2517
rect 3193 2512 3342 2517
rect 3385 2512 3430 2517
rect 1385 2507 1390 2512
rect 1801 2507 2014 2512
rect 2849 2507 2854 2512
rect 241 2502 286 2507
rect 281 2497 286 2502
rect 369 2502 414 2507
rect 889 2502 942 2507
rect 1233 2502 1278 2507
rect 1297 2502 1390 2507
rect 1625 2502 1726 2507
rect 2033 2502 2118 2507
rect 2137 2502 2214 2507
rect 2321 2502 2382 2507
rect 2577 2502 2606 2507
rect 2745 2502 2838 2507
rect 2849 2502 3038 2507
rect 3417 2502 3454 2507
rect 369 2497 374 2502
rect 2401 2497 2558 2502
rect 2625 2497 2726 2502
rect 0 2492 126 2497
rect 281 2492 374 2497
rect 393 2492 870 2497
rect 121 2487 126 2492
rect 121 2482 230 2487
rect 225 2477 230 2482
rect 393 2477 398 2492
rect 865 2487 870 2492
rect 993 2492 1126 2497
rect 1409 2492 1462 2497
rect 1481 2492 1606 2497
rect 993 2487 998 2492
rect 1481 2487 1486 2492
rect 865 2482 998 2487
rect 1321 2482 1390 2487
rect 1425 2482 1486 2487
rect 1601 2487 1606 2492
rect 1833 2492 2014 2497
rect 2241 2492 2406 2497
rect 2553 2492 2630 2497
rect 2721 2492 3022 2497
rect 3177 2492 3230 2497
rect 1833 2487 1838 2492
rect 2009 2487 2222 2492
rect 1601 2482 1646 2487
rect 1809 2482 1838 2487
rect 2217 2482 2718 2487
rect 2793 2482 3102 2487
rect 1321 2477 1326 2482
rect 225 2472 398 2477
rect 1217 2472 1326 2477
rect 1385 2477 1390 2482
rect 1385 2472 1502 2477
rect 1681 2472 1766 2477
rect 1833 2472 2686 2477
rect 2737 2472 2790 2477
rect 2809 2472 2838 2477
rect 2849 2472 2958 2477
rect 3129 2472 3270 2477
rect 1681 2467 1686 2472
rect 1145 2462 1686 2467
rect 1761 2467 1766 2472
rect 1761 2462 1790 2467
rect 2097 2462 2318 2467
rect 2377 2462 2742 2467
rect 2753 2462 3142 2467
rect 1969 2457 2078 2462
rect 2737 2457 2742 2462
rect 3161 2457 3294 2462
rect 545 2452 590 2457
rect 761 2452 846 2457
rect 1105 2452 1150 2457
rect 1193 2452 1462 2457
rect 1633 2452 1830 2457
rect 1945 2452 1974 2457
rect 2073 2452 2486 2457
rect 2513 2452 2694 2457
rect 2737 2452 2862 2457
rect 3097 2452 3166 2457
rect 3289 2452 3318 2457
rect 545 2447 550 2452
rect 481 2442 550 2447
rect 577 2442 606 2447
rect 633 2442 678 2447
rect 737 2442 782 2447
rect 793 2442 822 2447
rect 905 2442 966 2447
rect 1017 2442 1110 2447
rect 1233 2442 1342 2447
rect 1489 2442 1710 2447
rect 1993 2442 2430 2447
rect 2521 2442 2574 2447
rect 2697 2442 2950 2447
rect 3073 2442 3270 2447
rect 3337 2442 3406 2447
rect 1833 2437 1974 2442
rect 3337 2437 3342 2442
rect 385 2432 798 2437
rect 865 2432 1030 2437
rect 1089 2432 1118 2437
rect 1169 2432 1390 2437
rect 1401 2432 1574 2437
rect 1737 2432 1838 2437
rect 1969 2432 2934 2437
rect 2945 2432 3006 2437
rect 3025 2432 3342 2437
rect 3401 2437 3406 2442
rect 3401 2432 3438 2437
rect 1601 2427 1702 2432
rect 393 2422 430 2427
rect 505 2422 542 2427
rect 601 2422 902 2427
rect 897 2417 902 2422
rect 993 2417 998 2427
rect 1153 2422 1198 2427
rect 1289 2422 1502 2427
rect 1585 2422 1606 2427
rect 1697 2422 1726 2427
rect 1849 2422 2006 2427
rect 2057 2422 2118 2427
rect 2169 2422 2830 2427
rect 2913 2422 3022 2427
rect 3145 2422 3262 2427
rect 1193 2417 1294 2422
rect 1497 2417 1590 2422
rect 0 2412 6 2417
rect 489 2412 742 2417
rect 897 2412 982 2417
rect 993 2412 1094 2417
rect 1121 2412 1174 2417
rect 1313 2412 1422 2417
rect 1441 2412 1478 2417
rect 1609 2412 1662 2417
rect 1697 2412 2150 2417
rect 2281 2412 2614 2417
rect 2689 2412 2950 2417
rect 2977 2412 3390 2417
rect 1 2387 6 2412
rect 977 2407 982 2412
rect 1441 2407 1446 2412
rect 2145 2407 2286 2412
rect 433 2402 558 2407
rect 665 2402 774 2407
rect 977 2402 1110 2407
rect 1177 2402 1230 2407
rect 1305 2402 1446 2407
rect 1457 2402 1526 2407
rect 1985 2402 2126 2407
rect 2305 2402 2390 2407
rect 2409 2402 2542 2407
rect 2569 2402 2766 2407
rect 2785 2402 2806 2407
rect 2905 2402 3086 2407
rect 3185 2402 3358 2407
rect 3369 2402 3430 2407
rect 553 2397 670 2402
rect 1545 2397 1910 2402
rect 241 2392 286 2397
rect 457 2392 534 2397
rect 689 2392 790 2397
rect 841 2392 966 2397
rect 961 2387 966 2392
rect 1025 2392 1054 2397
rect 1065 2392 1094 2397
rect 1113 2392 1142 2397
rect 1241 2392 1550 2397
rect 1905 2392 2198 2397
rect 2225 2392 2278 2397
rect 2289 2392 3182 2397
rect 3193 2392 3366 2397
rect 1025 2387 1030 2392
rect 1137 2387 1246 2392
rect 2225 2387 2230 2392
rect 1 2382 230 2387
rect 321 2382 606 2387
rect 633 2382 702 2387
rect 961 2382 1030 2387
rect 1337 2382 1718 2387
rect 1769 2382 1870 2387
rect 1985 2382 2230 2387
rect 2257 2382 2686 2387
rect 2753 2382 2790 2387
rect 2873 2382 2918 2387
rect 2929 2382 3030 2387
rect 3073 2382 3318 2387
rect 225 2377 326 2382
rect 1889 2377 1990 2382
rect 537 2372 718 2377
rect 1049 2372 1422 2377
rect 1513 2372 1542 2377
rect 1657 2372 1894 2377
rect 2297 2372 2750 2377
rect 2793 2372 3014 2377
rect 3201 2372 3334 2377
rect 417 2367 518 2372
rect 1417 2367 1518 2372
rect 2009 2367 2278 2372
rect 185 2362 326 2367
rect 393 2362 422 2367
rect 513 2362 662 2367
rect 1353 2362 1398 2367
rect 1745 2362 1814 2367
rect 1185 2357 1334 2362
rect 1809 2357 1814 2362
rect 1905 2362 2014 2367
rect 2273 2362 2902 2367
rect 3033 2362 3158 2367
rect 3177 2362 3286 2367
rect 3345 2362 3406 2367
rect 1905 2357 1910 2362
rect 3033 2357 3038 2362
rect 257 2352 334 2357
rect 361 2352 510 2357
rect 521 2352 654 2357
rect 753 2352 782 2357
rect 849 2352 902 2357
rect 993 2352 1078 2357
rect 1161 2352 1190 2357
rect 1329 2352 1366 2357
rect 1473 2352 1614 2357
rect 1625 2352 1758 2357
rect 1809 2352 1910 2357
rect 2025 2352 2254 2357
rect 2297 2352 2478 2357
rect 2569 2352 2598 2357
rect 2609 2352 2918 2357
rect 3001 2352 3038 2357
rect 3153 2357 3158 2362
rect 3281 2357 3350 2362
rect 3153 2352 3174 2357
rect 1473 2347 1478 2352
rect 2473 2347 2574 2352
rect 3169 2347 3174 2352
rect 3233 2352 3262 2357
rect 3233 2347 3238 2352
rect 0 2342 70 2347
rect 89 2342 270 2347
rect 313 2342 422 2347
rect 457 2342 518 2347
rect 625 2342 654 2347
rect 745 2342 782 2347
rect 833 2342 886 2347
rect 969 2342 1070 2347
rect 1137 2342 1270 2347
rect 1289 2342 1326 2347
rect 1353 2342 1382 2347
rect 1433 2342 1478 2347
rect 1489 2342 1510 2347
rect 1545 2342 1790 2347
rect 1929 2342 2294 2347
rect 2369 2342 2454 2347
rect 2593 2342 2694 2347
rect 2737 2342 2870 2347
rect 2881 2342 2934 2347
rect 3001 2342 3150 2347
rect 3169 2342 3238 2347
rect 3313 2342 3342 2347
rect 65 2337 70 2342
rect 1265 2337 1270 2342
rect 2369 2337 2374 2342
rect 2689 2337 2694 2342
rect 65 2332 94 2337
rect 201 2332 270 2337
rect 385 2332 430 2337
rect 561 2332 814 2337
rect 1265 2332 1654 2337
rect 1897 2332 2294 2337
rect 2313 2332 2374 2337
rect 2473 2332 2574 2337
rect 2617 2332 2662 2337
rect 2689 2332 2790 2337
rect 89 2327 206 2332
rect 265 2327 374 2332
rect 881 2327 1006 2332
rect 1177 2327 1246 2332
rect 1745 2327 1878 2332
rect 2289 2327 2294 2332
rect 2393 2327 2478 2332
rect 2569 2327 2574 2332
rect 2865 2327 2870 2342
rect 2905 2332 3078 2337
rect 225 2322 246 2327
rect 369 2322 534 2327
rect 673 2322 782 2327
rect 817 2322 838 2327
rect 857 2322 886 2327
rect 1001 2322 1030 2327
rect 1065 2322 1182 2327
rect 1241 2322 1750 2327
rect 1873 2322 2102 2327
rect 2289 2322 2398 2327
rect 2569 2322 2814 2327
rect 2865 2322 3086 2327
rect 3169 2322 3294 2327
rect 225 2317 230 2322
rect 529 2317 662 2322
rect 0 2312 78 2317
rect 137 2312 230 2317
rect 329 2312 486 2317
rect 657 2312 806 2317
rect 865 2312 1006 2317
rect 1025 2312 1030 2322
rect 2121 2317 2270 2322
rect 3169 2317 3174 2322
rect 1193 2312 1486 2317
rect 1601 2312 1646 2317
rect 1761 2312 1998 2317
rect 2057 2312 2126 2317
rect 2265 2312 3030 2317
rect 3073 2312 3174 2317
rect 3289 2317 3294 2322
rect 3289 2312 3334 2317
rect 3385 2312 3422 2317
rect 801 2307 806 2312
rect 249 2302 598 2307
rect 657 2302 686 2307
rect 761 2302 790 2307
rect 801 2302 1118 2307
rect 1145 2302 1190 2307
rect 1233 2302 1526 2307
rect 1625 2302 1670 2307
rect 1857 2302 2134 2307
rect 2153 2302 2318 2307
rect 2385 2302 2534 2307
rect 2545 2302 2638 2307
rect 2673 2302 3038 2307
rect 3065 2302 3174 2307
rect 2129 2297 2134 2302
rect 3193 2297 3294 2302
rect 0 2292 30 2297
rect 25 2287 30 2292
rect 177 2292 526 2297
rect 865 2292 926 2297
rect 985 2292 1022 2297
rect 1225 2292 1510 2297
rect 1921 2292 1990 2297
rect 2129 2292 2214 2297
rect 2273 2292 2542 2297
rect 2769 2292 3198 2297
rect 3289 2292 3342 2297
rect 177 2287 182 2292
rect 25 2282 182 2287
rect 201 2282 398 2287
rect 449 2282 478 2287
rect 761 2282 806 2287
rect 905 2282 934 2287
rect 1193 2282 1246 2287
rect 1369 2282 1574 2287
rect 1593 2282 1838 2287
rect 2209 2282 2598 2287
rect 2681 2282 3070 2287
rect 3105 2282 3254 2287
rect 3289 2282 3414 2287
rect 1593 2277 1598 2282
rect 1833 2277 2006 2282
rect 281 2272 310 2277
rect 393 2272 446 2277
rect 1145 2272 1286 2277
rect 1361 2272 1406 2277
rect 1473 2272 1598 2277
rect 2001 2272 2726 2277
rect 2745 2272 2782 2277
rect 2857 2272 3038 2277
rect 3081 2272 3174 2277
rect 305 2267 398 2272
rect 2721 2267 2726 2272
rect 417 2262 502 2267
rect 521 2262 630 2267
rect 1313 2262 1462 2267
rect 1609 2262 1990 2267
rect 2297 2262 2438 2267
rect 2449 2262 2534 2267
rect 2721 2262 2910 2267
rect 2929 2262 3006 2267
rect 3129 2262 3230 2267
rect 521 2257 526 2262
rect 73 2252 526 2257
rect 625 2257 630 2262
rect 1177 2257 1318 2262
rect 1457 2257 1614 2262
rect 2009 2257 2214 2262
rect 2433 2257 2438 2262
rect 2529 2257 2534 2262
rect 625 2252 1046 2257
rect 1153 2252 1182 2257
rect 1329 2252 1438 2257
rect 1769 2252 2014 2257
rect 2209 2252 2406 2257
rect 2433 2252 2502 2257
rect 2529 2252 2790 2257
rect 2913 2252 3222 2257
rect 1153 2247 1158 2252
rect 1329 2247 1334 2252
rect 409 2242 574 2247
rect 601 2242 630 2247
rect 777 2242 886 2247
rect 1073 2242 1158 2247
rect 1177 2242 1334 2247
rect 1345 2242 1566 2247
rect 1585 2242 1694 2247
rect 1713 2242 2014 2247
rect 2049 2242 2094 2247
rect 2121 2242 2198 2247
rect 2297 2242 2678 2247
rect 2865 2242 3166 2247
rect 1585 2237 1590 2242
rect 177 2232 222 2237
rect 249 2232 286 2237
rect 281 2227 286 2232
rect 409 2232 462 2237
rect 473 2232 622 2237
rect 641 2232 742 2237
rect 809 2232 950 2237
rect 1121 2232 1174 2237
rect 1185 2232 1310 2237
rect 1457 2232 1590 2237
rect 1689 2237 1694 2242
rect 1689 2232 1750 2237
rect 1841 2232 2158 2237
rect 2185 2232 2230 2237
rect 2417 2232 2566 2237
rect 2625 2232 2742 2237
rect 2761 2232 3014 2237
rect 3257 2232 3318 2237
rect 409 2227 414 2232
rect 1329 2227 1438 2232
rect 1745 2227 1846 2232
rect 2329 2227 2398 2232
rect 281 2222 414 2227
rect 433 2222 750 2227
rect 1073 2222 1334 2227
rect 1433 2222 1726 2227
rect 1865 2222 2334 2227
rect 2393 2222 2462 2227
rect 2529 2222 2678 2227
rect 2873 2222 3062 2227
rect 3393 2222 3430 2227
rect 2737 2217 2838 2222
rect 505 2212 550 2217
rect 577 2212 638 2217
rect 689 2212 846 2217
rect 1009 2212 1094 2217
rect 1113 2212 1654 2217
rect 1769 2212 2038 2217
rect 2217 2212 2254 2217
rect 2345 2212 2390 2217
rect 2505 2212 2550 2217
rect 2681 2212 2742 2217
rect 2833 2212 2974 2217
rect 3081 2212 3238 2217
rect 545 2207 550 2212
rect 1089 2207 1094 2212
rect 2057 2207 2198 2212
rect 2569 2207 2662 2212
rect 3081 2207 3086 2212
rect 217 2202 262 2207
rect 473 2202 526 2207
rect 545 2202 654 2207
rect 1089 2202 1118 2207
rect 1217 2202 1806 2207
rect 1841 2202 2062 2207
rect 2193 2202 2574 2207
rect 2657 2202 2918 2207
rect 2985 2202 3086 2207
rect 3233 2207 3238 2212
rect 3233 2202 3302 2207
rect 3361 2202 3414 2207
rect 1113 2197 1222 2202
rect 1841 2197 1846 2202
rect 2913 2197 2990 2202
rect 3105 2197 3214 2202
rect 3425 2197 3430 2222
rect 113 2192 254 2197
rect 297 2192 350 2197
rect 441 2192 486 2197
rect 561 2192 806 2197
rect 913 2192 1014 2197
rect 1073 2192 1094 2197
rect 1241 2192 1494 2197
rect 1561 2192 1670 2197
rect 1785 2192 1846 2197
rect 1865 2192 1942 2197
rect 1985 2192 2574 2197
rect 2617 2192 2894 2197
rect 3041 2192 3110 2197
rect 3209 2192 3294 2197
rect 3385 2192 3430 2197
rect 449 2182 750 2187
rect 1049 2182 1462 2187
rect 1865 2182 2390 2187
rect 2401 2182 3094 2187
rect 3113 2182 3230 2187
rect 3281 2182 3318 2187
rect 3089 2177 3094 2182
rect 569 2172 598 2177
rect 609 2172 678 2177
rect 793 2172 902 2177
rect 985 2172 1054 2177
rect 1201 2172 1262 2177
rect 1433 2172 1486 2177
rect 1505 2172 1606 2177
rect 1833 2172 2358 2177
rect 2417 2172 2790 2177
rect 2897 2172 2950 2177
rect 3089 2172 3142 2177
rect 1281 2167 1414 2172
rect 1505 2167 1510 2172
rect 129 2162 374 2167
rect 729 2162 982 2167
rect 1065 2162 1286 2167
rect 1409 2162 1510 2167
rect 1601 2167 1606 2172
rect 3177 2167 3246 2172
rect 3305 2167 3374 2172
rect 1601 2162 1630 2167
rect 1649 2162 1726 2167
rect 1945 2162 2030 2167
rect 2129 2162 2318 2167
rect 2337 2162 3182 2167
rect 3241 2162 3310 2167
rect 3369 2162 3398 2167
rect 129 2157 134 2162
rect 0 2152 134 2157
rect 369 2157 374 2162
rect 977 2157 1070 2162
rect 1649 2157 1654 2162
rect 369 2152 838 2157
rect 1209 2152 1654 2157
rect 1721 2157 1726 2162
rect 1721 2152 2510 2157
rect 2553 2152 2646 2157
rect 2705 2152 2966 2157
rect 1209 2147 1214 2152
rect 313 2142 358 2147
rect 457 2142 598 2147
rect 145 2132 254 2137
rect 489 2132 710 2137
rect 721 2127 726 2147
rect 737 2142 822 2147
rect 937 2142 1030 2147
rect 1105 2142 1214 2147
rect 1233 2142 1262 2147
rect 1353 2142 1518 2147
rect 1841 2142 1870 2147
rect 2153 2142 2262 2147
rect 2273 2142 2358 2147
rect 2377 2142 2838 2147
rect 2881 2142 3134 2147
rect 569 2122 726 2127
rect 817 2127 822 2142
rect 841 2127 998 2132
rect 817 2122 846 2127
rect 993 2122 1022 2127
rect 433 2112 558 2117
rect 257 2102 462 2107
rect 473 2102 518 2107
rect 553 2097 558 2112
rect 697 2112 758 2117
rect 841 2112 974 2117
rect 697 2097 702 2112
rect 1105 2107 1110 2142
rect 1257 2137 1358 2142
rect 1537 2137 1606 2142
rect 1865 2137 2158 2142
rect 3153 2137 3158 2162
rect 3177 2152 3230 2157
rect 3321 2152 3422 2157
rect 3241 2142 3310 2147
rect 3385 2142 3414 2147
rect 3305 2137 3390 2142
rect 1497 2132 1542 2137
rect 1601 2132 1710 2137
rect 2177 2132 2518 2137
rect 2569 2132 2902 2137
rect 3153 2132 3230 2137
rect 2961 2127 3094 2132
rect 1177 2122 1382 2127
rect 1393 2122 1430 2127
rect 1545 2122 1590 2127
rect 1881 2122 2158 2127
rect 2177 2122 2422 2127
rect 2465 2122 2678 2127
rect 2713 2122 2966 2127
rect 3089 2122 3118 2127
rect 3345 2122 3374 2127
rect 1609 2117 1710 2122
rect 2177 2117 2182 2122
rect 2673 2117 2678 2122
rect 1121 2112 1614 2117
rect 1705 2112 1734 2117
rect 1945 2112 1990 2117
rect 2129 2112 2182 2117
rect 2193 2112 2342 2117
rect 2369 2112 2406 2117
rect 2425 2112 2630 2117
rect 2673 2112 3062 2117
rect 3129 2112 3286 2117
rect 2001 2107 2134 2112
rect 3057 2107 3134 2112
rect 801 2102 886 2107
rect 881 2097 886 2102
rect 977 2102 1006 2107
rect 1025 2102 1110 2107
rect 1137 2102 1270 2107
rect 1289 2102 1318 2107
rect 977 2097 982 2102
rect 1313 2097 1318 2102
rect 1433 2102 1542 2107
rect 1601 2102 1726 2107
rect 1857 2102 1926 2107
rect 1961 2102 2006 2107
rect 2153 2102 2382 2107
rect 2465 2102 2574 2107
rect 2601 2102 2686 2107
rect 2721 2102 2774 2107
rect 2849 2102 2918 2107
rect 2953 2102 3038 2107
rect 3241 2102 3262 2107
rect 1433 2097 1438 2102
rect 1857 2097 1862 2102
rect 401 2092 502 2097
rect 553 2092 702 2097
rect 721 2092 758 2097
rect 833 2092 862 2097
rect 881 2092 982 2097
rect 1081 2092 1110 2097
rect 1313 2092 1438 2097
rect 1833 2092 1862 2097
rect 1921 2097 1926 2102
rect 1921 2092 2710 2097
rect 2761 2092 2910 2097
rect 3057 2092 3150 2097
rect 3233 2092 3262 2097
rect 857 2077 862 2092
rect 1081 2077 1086 2092
rect 2929 2087 3062 2092
rect 3145 2087 3150 2092
rect 1105 2082 1134 2087
rect 857 2072 1086 2077
rect 1129 2077 1134 2082
rect 1249 2082 1286 2087
rect 1689 2082 1822 2087
rect 1937 2082 1966 2087
rect 2129 2082 2470 2087
rect 2481 2082 2726 2087
rect 2897 2082 2934 2087
rect 3145 2082 3174 2087
rect 1249 2077 1254 2082
rect 1817 2077 1942 2082
rect 2721 2077 2814 2082
rect 1129 2072 1254 2077
rect 1369 2072 1406 2077
rect 2169 2072 2358 2077
rect 2449 2072 2710 2077
rect 2809 2072 2838 2077
rect 2889 2072 3350 2077
rect 1449 2062 1670 2067
rect 1273 2052 1318 2057
rect 1393 2052 1414 2057
rect 1449 2047 1454 2062
rect 281 2042 366 2047
rect 1281 2042 1374 2047
rect 1425 2042 1454 2047
rect 1665 2047 1670 2062
rect 1841 2062 2110 2067
rect 2193 2062 2934 2067
rect 3273 2062 3454 2067
rect 1841 2057 1846 2062
rect 1817 2052 1846 2057
rect 2105 2057 2110 2062
rect 2929 2057 3014 2062
rect 3273 2057 3278 2062
rect 2105 2052 2390 2057
rect 2433 2052 2486 2057
rect 2537 2052 2590 2057
rect 2625 2052 2814 2057
rect 3009 2052 3278 2057
rect 1665 2042 1790 2047
rect 1841 2042 1918 2047
rect 1961 2042 2014 2047
rect 2137 2042 2190 2047
rect 2241 2042 2318 2047
rect 2593 2042 2686 2047
rect 2737 2042 2830 2047
rect 2849 2042 2990 2047
rect 281 2037 286 2042
rect 257 2032 286 2037
rect 361 2037 366 2042
rect 2337 2037 2574 2042
rect 2849 2037 2854 2042
rect 361 2032 462 2037
rect 625 2032 710 2037
rect 785 2032 814 2037
rect 1017 2032 1078 2037
rect 1169 2032 1758 2037
rect 1897 2032 1926 2037
rect 2025 2032 2342 2037
rect 2569 2032 2646 2037
rect 2657 2032 2854 2037
rect 2985 2037 2990 2042
rect 2985 2032 3182 2037
rect 3225 2032 3294 2037
rect 3313 2032 3398 2037
rect 1921 2027 2030 2032
rect 2641 2027 2646 2032
rect 3225 2027 3230 2032
rect 273 2022 350 2027
rect 497 2022 534 2027
rect 569 2022 598 2027
rect 817 2022 990 2027
rect 1025 2022 1086 2027
rect 1193 2022 1278 2027
rect 1313 2022 1366 2027
rect 1553 2022 1686 2027
rect 1385 2017 1534 2022
rect 1697 2017 1702 2027
rect 2057 2022 2190 2027
rect 2209 2022 2254 2027
rect 2329 2022 2550 2027
rect 2641 2022 2878 2027
rect 2889 2022 2974 2027
rect 3201 2022 3230 2027
rect 3289 2027 3294 2032
rect 3289 2022 3310 2027
rect 2209 2017 2214 2022
rect 3305 2017 3310 2022
rect 3393 2022 3422 2027
rect 3393 2017 3398 2022
rect 505 2012 542 2017
rect 649 2012 766 2017
rect 833 2007 838 2017
rect 1265 2012 1326 2017
rect 1345 2012 1390 2017
rect 1529 2012 1702 2017
rect 1777 2012 2030 2017
rect 2049 2012 2214 2017
rect 2321 2012 2542 2017
rect 2649 2012 2718 2017
rect 2793 2012 2886 2017
rect 3153 2012 3172 2017
rect 3241 2012 3278 2017
rect 3305 2012 3398 2017
rect 1345 2007 1350 2012
rect 1777 2007 1782 2012
rect 169 2002 238 2007
rect 433 2002 806 2007
rect 817 2002 838 2007
rect 953 2002 1046 2007
rect 1073 2002 1182 2007
rect 1241 2002 1286 2007
rect 1297 2002 1350 2007
rect 1409 2002 1782 2007
rect 2025 2007 2030 2012
rect 3167 2007 3172 2012
rect 2025 2002 2766 2007
rect 2777 2002 2854 2007
rect 2905 2002 3126 2007
rect 3167 2002 3182 2007
rect 169 1997 174 2002
rect 0 1992 134 1997
rect 145 1992 174 1997
rect 233 1997 238 2002
rect 2905 1997 2910 2002
rect 233 1992 262 1997
rect 449 1992 702 1997
rect 793 1992 838 1997
rect 985 1992 1022 1997
rect 1065 1992 1574 1997
rect 1657 1992 1726 1997
rect 1793 1992 2406 1997
rect 2449 1992 2806 1997
rect 2825 1992 2910 1997
rect 3121 1997 3126 2002
rect 3121 1992 3150 1997
rect 3297 1992 3342 1997
rect 129 1977 134 1992
rect 1569 1987 1662 1992
rect 1721 1987 1798 1992
rect 2801 1987 2806 1992
rect 273 1982 446 1987
rect 473 1982 630 1987
rect 713 1982 790 1987
rect 825 1982 870 1987
rect 1001 1982 1294 1987
rect 1313 1982 1446 1987
rect 1473 1982 1550 1987
rect 1681 1982 1702 1987
rect 1977 1982 2118 1987
rect 2145 1982 2430 1987
rect 2585 1982 2750 1987
rect 2801 1982 2902 1987
rect 2953 1982 2998 1987
rect 3041 1982 3350 1987
rect 273 1977 278 1982
rect 625 1977 718 1982
rect 1697 1977 1702 1982
rect 129 1972 278 1977
rect 465 1972 526 1977
rect 785 1972 814 1977
rect 881 1972 1118 1977
rect 1185 1972 1206 1977
rect 1281 1972 1638 1977
rect 1697 1972 1854 1977
rect 1905 1972 2182 1977
rect 2289 1972 2550 1977
rect 2857 1972 2918 1977
rect 2945 1972 2982 1977
rect 2993 1972 3198 1977
rect 809 1967 886 1972
rect 2177 1967 2294 1972
rect 2569 1967 2710 1972
rect 2745 1967 2838 1972
rect 2945 1967 2950 1972
rect 449 1962 486 1967
rect 585 1962 782 1967
rect 993 1962 1086 1967
rect 1417 1962 1454 1967
rect 1489 1962 1630 1967
rect 1785 1962 2158 1967
rect 2313 1962 2574 1967
rect 2705 1962 2750 1967
rect 2833 1962 2950 1967
rect 1241 1957 1398 1962
rect 1649 1957 1766 1962
rect 2969 1957 3070 1962
rect 401 1952 846 1957
rect 1009 1952 1062 1957
rect 1161 1952 1246 1957
rect 1393 1952 1654 1957
rect 1761 1952 1854 1957
rect 1993 1952 2054 1957
rect 2073 1952 2206 1957
rect 2217 1952 2310 1957
rect 2337 1952 2694 1957
rect 2761 1952 2910 1957
rect 2937 1952 2974 1957
rect 3065 1952 3094 1957
rect 3289 1952 3326 1957
rect 1993 1947 1998 1952
rect 161 1942 254 1947
rect 281 1942 342 1947
rect 425 1942 486 1947
rect 569 1942 750 1947
rect 961 1942 1086 1947
rect 1097 1942 1182 1947
rect 1257 1942 1318 1947
rect 1337 1942 1430 1947
rect 1457 1942 1558 1947
rect 1609 1942 1774 1947
rect 1873 1942 1998 1947
rect 2017 1942 2438 1947
rect 2609 1942 2830 1947
rect 2881 1942 3086 1947
rect 3113 1942 3206 1947
rect 161 1937 166 1942
rect 1313 1937 1318 1942
rect 1873 1937 1878 1942
rect 2473 1937 2590 1942
rect 3113 1937 3118 1942
rect 137 1932 166 1937
rect 217 1932 262 1937
rect 673 1932 790 1937
rect 873 1932 1190 1937
rect 1313 1932 1878 1937
rect 2041 1932 2070 1937
rect 2097 1932 2166 1937
rect 2225 1932 2326 1937
rect 2345 1932 2478 1937
rect 2585 1932 2774 1937
rect 2881 1932 3118 1937
rect 3201 1937 3206 1942
rect 3201 1932 3230 1937
rect 3393 1932 3414 1937
rect 321 1927 406 1932
rect 593 1927 678 1932
rect 2769 1927 2886 1932
rect 249 1922 326 1927
rect 401 1922 430 1927
rect 441 1922 598 1927
rect 865 1922 1214 1927
rect 1345 1922 1518 1927
rect 1577 1922 1646 1927
rect 1761 1922 1798 1927
rect 1897 1922 1998 1927
rect 2049 1922 2246 1927
rect 2281 1922 2390 1927
rect 2489 1922 2750 1927
rect 2905 1922 2934 1927
rect 3041 1922 3318 1927
rect 1817 1917 1902 1922
rect 1993 1917 1998 1922
rect 2385 1917 2494 1922
rect 2929 1917 3046 1922
rect 337 1912 422 1917
rect 569 1912 630 1917
rect 897 1912 1006 1917
rect 1089 1912 1334 1917
rect 1417 1912 1822 1917
rect 1993 1912 2358 1917
rect 2513 1912 2662 1917
rect 2705 1912 2806 1917
rect 3065 1912 3118 1917
rect 3193 1912 3414 1917
rect 1329 1907 1422 1912
rect 0 1902 238 1907
rect 233 1897 238 1902
rect 353 1902 1206 1907
rect 1441 1902 1790 1907
rect 1849 1902 2422 1907
rect 2433 1902 2686 1907
rect 2705 1902 2710 1912
rect 2737 1902 2774 1907
rect 2833 1902 2966 1907
rect 3057 1902 3094 1907
rect 3201 1902 3230 1907
rect 3321 1902 3422 1907
rect 353 1897 358 1902
rect 233 1892 358 1897
rect 425 1892 454 1897
rect 449 1887 454 1892
rect 593 1892 638 1897
rect 769 1892 798 1897
rect 593 1887 598 1892
rect 449 1882 598 1887
rect 793 1887 798 1892
rect 889 1892 950 1897
rect 1049 1892 1102 1897
rect 1337 1892 1374 1897
rect 1449 1892 1494 1897
rect 1697 1892 2822 1897
rect 2833 1892 3038 1897
rect 3161 1892 3430 1897
rect 889 1887 894 1892
rect 1513 1887 1670 1892
rect 2817 1887 2822 1892
rect 793 1882 894 1887
rect 913 1882 958 1887
rect 1193 1882 1518 1887
rect 1665 1882 1694 1887
rect 1689 1877 1694 1882
rect 1809 1882 2094 1887
rect 2313 1882 2518 1887
rect 2577 1882 2782 1887
rect 2817 1882 2910 1887
rect 1809 1877 1814 1882
rect 2153 1877 2294 1882
rect 2905 1877 2910 1882
rect 3049 1882 3150 1887
rect 3049 1877 3054 1882
rect 1369 1872 1670 1877
rect 1689 1872 1814 1877
rect 1993 1872 2086 1877
rect 2129 1872 2158 1877
rect 2289 1872 2886 1877
rect 2905 1872 3054 1877
rect 3145 1877 3150 1882
rect 3273 1882 3342 1887
rect 3273 1877 3278 1882
rect 3145 1872 3278 1877
rect 1857 1867 1974 1872
rect 1393 1862 1550 1867
rect 1833 1862 1862 1867
rect 1969 1862 2782 1867
rect 25 1852 182 1857
rect 201 1852 302 1857
rect 489 1852 518 1857
rect 1089 1852 1166 1857
rect 1241 1852 1350 1857
rect 1417 1852 1470 1857
rect 1521 1852 1574 1857
rect 1593 1852 1694 1857
rect 1745 1852 2030 1857
rect 2041 1852 2062 1857
rect 2137 1852 2174 1857
rect 2433 1852 2478 1857
rect 2697 1852 2734 1857
rect 2889 1852 3094 1857
rect 3113 1852 3318 1857
rect 25 1847 30 1852
rect 0 1842 30 1847
rect 177 1847 182 1852
rect 1593 1847 1598 1852
rect 177 1842 406 1847
rect 1169 1842 1294 1847
rect 1345 1842 1406 1847
rect 1505 1842 1598 1847
rect 1689 1847 1694 1852
rect 2193 1847 2358 1852
rect 2497 1847 2598 1852
rect 1689 1842 1718 1847
rect 1793 1842 2198 1847
rect 2353 1842 2502 1847
rect 2593 1842 2758 1847
rect 3113 1837 3118 1852
rect 73 1832 158 1837
rect 553 1832 646 1837
rect 689 1832 710 1837
rect 1089 1832 2342 1837
rect 2497 1832 2782 1837
rect 2817 1832 2990 1837
rect 3009 1832 3118 1837
rect 3313 1837 3318 1852
rect 3313 1832 3342 1837
rect 73 1827 78 1832
rect 153 1827 366 1832
rect 2817 1827 2822 1832
rect 0 1822 78 1827
rect 361 1822 430 1827
rect 489 1822 542 1827
rect 937 1822 1046 1827
rect 1065 1822 1150 1827
rect 1193 1822 1838 1827
rect 1985 1822 2822 1827
rect 3081 1822 3390 1827
rect 1857 1817 1966 1822
rect 89 1812 222 1817
rect 241 1812 350 1817
rect 433 1812 694 1817
rect 1217 1812 1286 1817
rect 1401 1812 1430 1817
rect 1537 1812 1862 1817
rect 1961 1812 2142 1817
rect 2353 1812 2406 1817
rect 2505 1812 2574 1817
rect 2649 1812 2686 1817
rect 2769 1812 2846 1817
rect 2857 1812 2918 1817
rect 2985 1812 3070 1817
rect 1425 1807 1542 1812
rect 2161 1807 2334 1812
rect 193 1802 526 1807
rect 193 1792 198 1802
rect 521 1797 526 1802
rect 649 1802 814 1807
rect 1001 1802 1086 1807
rect 1113 1802 1390 1807
rect 1737 1802 1902 1807
rect 1961 1802 2102 1807
rect 2121 1802 2166 1807
rect 2329 1802 2670 1807
rect 2769 1802 2774 1812
rect 2897 1802 3014 1807
rect 649 1797 654 1802
rect 1561 1797 1686 1802
rect 3265 1797 3270 1822
rect 3289 1812 3358 1817
rect 3329 1802 3406 1807
rect 257 1792 286 1797
rect 281 1787 286 1792
rect 345 1792 374 1797
rect 417 1792 462 1797
rect 521 1792 654 1797
rect 689 1792 734 1797
rect 905 1792 1078 1797
rect 1289 1792 1374 1797
rect 1409 1792 1454 1797
rect 1497 1792 1566 1797
rect 1681 1792 1750 1797
rect 1761 1792 1790 1797
rect 1881 1792 2718 1797
rect 2737 1792 2766 1797
rect 2833 1792 2934 1797
rect 2969 1792 3094 1797
rect 3265 1792 3350 1797
rect 345 1787 350 1792
rect 1073 1787 1254 1792
rect 145 1782 222 1787
rect 281 1782 350 1787
rect 409 1782 430 1787
rect 465 1782 502 1787
rect 673 1782 814 1787
rect 1249 1782 1446 1787
rect 1577 1782 1726 1787
rect 1745 1777 1750 1792
rect 1785 1787 1886 1792
rect 1905 1782 2478 1787
rect 2489 1782 2526 1787
rect 2561 1782 2758 1787
rect 2777 1782 2886 1787
rect 3049 1782 3134 1787
rect 3321 1782 3390 1787
rect 2881 1777 3054 1782
rect 401 1772 454 1777
rect 569 1772 622 1777
rect 649 1772 710 1777
rect 1017 1772 1126 1777
rect 1185 1772 1614 1777
rect 1745 1772 2206 1777
rect 2305 1772 2438 1777
rect 2481 1772 2862 1777
rect 3073 1772 3190 1777
rect 313 1762 790 1767
rect 1105 1762 1214 1767
rect 1265 1762 1318 1767
rect 1369 1762 1566 1767
rect 1697 1762 1766 1767
rect 1945 1762 1998 1767
rect 2081 1762 2118 1767
rect 2185 1762 2286 1767
rect 2417 1762 2470 1767
rect 2481 1762 2574 1767
rect 2617 1762 2870 1767
rect 2913 1762 2950 1767
rect 3209 1762 3294 1767
rect 1825 1757 1926 1762
rect 2305 1757 2398 1762
rect 3209 1757 3214 1762
rect 609 1752 702 1757
rect 1113 1752 1134 1757
rect 1201 1752 1406 1757
rect 1425 1752 1494 1757
rect 1585 1752 1678 1757
rect 1801 1752 1830 1757
rect 1921 1752 2310 1757
rect 2393 1752 3214 1757
rect 3289 1757 3294 1762
rect 3289 1752 3318 1757
rect 3337 1752 3414 1757
rect 361 1747 494 1752
rect 1585 1747 1590 1752
rect 1673 1747 1782 1752
rect 3337 1747 3342 1752
rect 145 1742 254 1747
rect 337 1742 366 1747
rect 489 1742 646 1747
rect 873 1742 902 1747
rect 1121 1742 1590 1747
rect 1777 1742 1822 1747
rect 1865 1742 2198 1747
rect 2249 1742 2342 1747
rect 2353 1742 2422 1747
rect 2433 1742 2470 1747
rect 2481 1742 2542 1747
rect 2633 1742 2678 1747
rect 2705 1742 2742 1747
rect 2761 1742 2806 1747
rect 2833 1742 2862 1747
rect 2953 1742 3078 1747
rect 3097 1742 3342 1747
rect 3409 1747 3414 1752
rect 3409 1742 3438 1747
rect 2737 1737 2742 1742
rect 2833 1737 2838 1742
rect 2857 1737 2958 1742
rect 3073 1737 3078 1742
rect 353 1732 478 1737
rect 609 1732 670 1737
rect 1129 1732 1318 1737
rect 1329 1732 1382 1737
rect 1393 1732 1798 1737
rect 1985 1732 2558 1737
rect 2657 1732 2718 1737
rect 2737 1732 2758 1737
rect 2785 1732 2838 1737
rect 2977 1732 3054 1737
rect 3073 1732 3398 1737
rect 1793 1727 1990 1732
rect 313 1722 350 1727
rect 489 1722 630 1727
rect 873 1722 942 1727
rect 1049 1722 1414 1727
rect 1505 1722 1558 1727
rect 1609 1722 1774 1727
rect 2009 1722 2086 1727
rect 2145 1722 2966 1727
rect 345 1717 494 1722
rect 625 1717 694 1722
rect 2961 1717 2966 1722
rect 3257 1722 3414 1727
rect 3257 1717 3262 1722
rect 297 1712 326 1717
rect 545 1712 606 1717
rect 689 1712 758 1717
rect 817 1712 870 1717
rect 905 1712 1046 1717
rect 1081 1712 1166 1717
rect 1177 1712 1230 1717
rect 1313 1712 1398 1717
rect 1489 1712 1574 1717
rect 1721 1712 1782 1717
rect 1889 1712 1966 1717
rect 1985 1712 2030 1717
rect 2113 1712 2470 1717
rect 2481 1712 2526 1717
rect 2609 1712 2854 1717
rect 2961 1712 3262 1717
rect 3297 1712 3374 1717
rect 1393 1707 1398 1712
rect 1889 1707 1894 1712
rect 449 1702 518 1707
rect 641 1702 678 1707
rect 1001 1702 1030 1707
rect 1089 1702 1118 1707
rect 1113 1697 1118 1702
rect 1241 1702 1374 1707
rect 1393 1702 1430 1707
rect 1449 1702 1710 1707
rect 1865 1702 1894 1707
rect 1961 1707 1966 1712
rect 1961 1702 2486 1707
rect 2537 1702 2598 1707
rect 2697 1702 2734 1707
rect 2873 1702 2942 1707
rect 3281 1702 3318 1707
rect 1241 1697 1246 1702
rect 1425 1697 1430 1702
rect 2873 1697 2878 1702
rect 249 1692 350 1697
rect 881 1692 1054 1697
rect 1113 1692 1246 1697
rect 1329 1692 1398 1697
rect 1425 1692 1598 1697
rect 1689 1692 1758 1697
rect 1889 1692 1942 1697
rect 1969 1692 2014 1697
rect 2033 1692 2126 1697
rect 2153 1692 2262 1697
rect 2321 1692 2502 1697
rect 2537 1692 2878 1697
rect 2937 1697 2942 1702
rect 2937 1692 2966 1697
rect 2985 1692 3262 1697
rect 3289 1692 3414 1697
rect 1425 1687 1430 1692
rect 2033 1687 2038 1692
rect 2985 1687 2990 1692
rect 1009 1682 1062 1687
rect 1297 1682 1390 1687
rect 1401 1682 1430 1687
rect 1449 1682 1510 1687
rect 1929 1682 2038 1687
rect 2057 1682 2254 1687
rect 2345 1682 2758 1687
rect 2865 1682 2990 1687
rect 3257 1687 3262 1692
rect 3257 1682 3286 1687
rect 3377 1682 3438 1687
rect 2753 1677 2870 1682
rect 1121 1672 1174 1677
rect 1305 1672 1518 1677
rect 1009 1667 1102 1672
rect 457 1662 526 1667
rect 577 1662 654 1667
rect 689 1662 966 1667
rect 985 1662 1014 1667
rect 1097 1662 1142 1667
rect 689 1657 694 1662
rect 393 1652 694 1657
rect 961 1657 966 1662
rect 961 1652 1110 1657
rect 145 1642 374 1647
rect 409 1642 542 1647
rect 713 1642 830 1647
rect 865 1642 926 1647
rect 145 1637 150 1642
rect 0 1632 150 1637
rect 369 1637 374 1642
rect 713 1637 718 1642
rect 369 1632 422 1637
rect 609 1632 718 1637
rect 825 1637 830 1642
rect 825 1632 854 1637
rect 961 1632 1094 1637
rect 849 1627 966 1632
rect 1121 1627 1126 1662
rect 1169 1657 1174 1672
rect 1513 1667 1518 1672
rect 1609 1672 1678 1677
rect 1609 1667 1614 1672
rect 1225 1662 1494 1667
rect 1513 1662 1614 1667
rect 1673 1667 1678 1672
rect 1753 1672 2494 1677
rect 2569 1672 2646 1677
rect 2689 1672 2734 1677
rect 2889 1672 3182 1677
rect 1753 1667 1758 1672
rect 1673 1662 1758 1667
rect 1945 1662 2190 1667
rect 2209 1662 3382 1667
rect 1857 1657 1926 1662
rect 1169 1652 1422 1657
rect 1441 1652 1462 1657
rect 1777 1652 1862 1657
rect 1921 1652 2086 1657
rect 2377 1652 3094 1657
rect 2081 1647 2382 1652
rect 3089 1647 3094 1652
rect 3177 1652 3206 1657
rect 3177 1647 3182 1652
rect 1185 1642 1486 1647
rect 1873 1642 2062 1647
rect 2401 1642 2446 1647
rect 2473 1642 2646 1647
rect 2657 1642 2806 1647
rect 3089 1642 3182 1647
rect 2825 1637 3046 1642
rect 1169 1632 1246 1637
rect 1289 1632 1510 1637
rect 1529 1632 1606 1637
rect 1681 1632 1774 1637
rect 1873 1632 1950 1637
rect 1985 1632 2086 1637
rect 2121 1632 2254 1637
rect 2313 1632 2830 1637
rect 3041 1632 3070 1637
rect 3241 1632 3318 1637
rect 1529 1627 1534 1632
rect 281 1622 326 1627
rect 337 1622 494 1627
rect 505 1622 814 1627
rect 993 1622 1046 1627
rect 1057 1622 1126 1627
rect 1209 1622 1326 1627
rect 1425 1622 1454 1627
rect 1497 1622 1534 1627
rect 1601 1627 1606 1632
rect 1601 1622 1630 1627
rect 1737 1622 2454 1627
rect 2497 1622 3142 1627
rect 3297 1622 3358 1627
rect 337 1617 342 1622
rect 161 1612 342 1617
rect 425 1612 606 1617
rect 697 1612 742 1617
rect 913 1612 950 1617
rect 1057 1607 1062 1622
rect 2449 1617 2454 1622
rect 1097 1612 1198 1617
rect 1337 1612 1798 1617
rect 1849 1612 1894 1617
rect 1929 1612 1966 1617
rect 2009 1612 2190 1617
rect 2305 1612 2430 1617
rect 2449 1612 2598 1617
rect 2641 1612 2694 1617
rect 2713 1612 2798 1617
rect 2897 1612 3022 1617
rect 3097 1612 3150 1617
rect 3201 1612 3270 1617
rect 1193 1607 1342 1612
rect 121 1602 174 1607
rect 225 1602 326 1607
rect 521 1602 582 1607
rect 641 1602 694 1607
rect 721 1602 886 1607
rect 945 1602 1062 1607
rect 1105 1602 1174 1607
rect 1409 1602 1542 1607
rect 1825 1602 2126 1607
rect 2153 1602 2214 1607
rect 2225 1602 2510 1607
rect 2529 1602 2886 1607
rect 2929 1602 3078 1607
rect 3289 1602 3374 1607
rect 401 1597 502 1602
rect 89 1592 118 1597
rect 113 1587 118 1592
rect 177 1592 206 1597
rect 249 1592 358 1597
rect 377 1592 406 1597
rect 497 1592 742 1597
rect 833 1592 870 1597
rect 177 1587 182 1592
rect 0 1582 78 1587
rect 113 1582 182 1587
rect 369 1582 654 1587
rect 809 1582 830 1587
rect 73 1567 78 1582
rect 369 1567 374 1582
rect 489 1572 550 1577
rect 561 1572 590 1577
rect 617 1572 646 1577
rect 857 1572 918 1577
rect 945 1572 950 1602
rect 1825 1597 1830 1602
rect 2209 1597 2214 1602
rect 1041 1592 1126 1597
rect 1185 1592 1246 1597
rect 1305 1592 1414 1597
rect 1441 1592 1478 1597
rect 1593 1592 1702 1597
rect 1809 1592 1830 1597
rect 1865 1592 2030 1597
rect 2049 1592 2086 1597
rect 2121 1592 2198 1597
rect 2209 1592 2302 1597
rect 2321 1592 2414 1597
rect 2425 1592 2518 1597
rect 2545 1592 2918 1597
rect 3033 1592 3102 1597
rect 3121 1592 3198 1597
rect 3241 1592 3318 1597
rect 1041 1587 1046 1592
rect 969 1582 1046 1587
rect 1057 1582 1078 1587
rect 1137 1582 1206 1587
rect 1417 1582 1494 1587
rect 1569 1582 1766 1587
rect 1297 1577 1398 1582
rect 1809 1577 1814 1592
rect 3121 1587 3126 1592
rect 1825 1582 1870 1587
rect 2033 1582 2950 1587
rect 2961 1582 3038 1587
rect 3073 1582 3126 1587
rect 3193 1587 3198 1592
rect 3193 1582 3222 1587
rect 3233 1582 3374 1587
rect 1889 1577 2014 1582
rect 3233 1577 3238 1582
rect 993 1572 1302 1577
rect 1393 1572 1446 1577
rect 1457 1572 1614 1577
rect 1681 1572 1814 1577
rect 1841 1572 1894 1577
rect 2009 1572 2062 1577
rect 2129 1572 2278 1577
rect 2329 1572 2622 1577
rect 2657 1572 2726 1577
rect 2793 1572 3238 1577
rect 3257 1572 3318 1577
rect 913 1567 918 1572
rect 73 1562 374 1567
rect 433 1562 510 1567
rect 553 1562 726 1567
rect 801 1562 902 1567
rect 913 1562 942 1567
rect 1041 1562 1150 1567
rect 1313 1562 1670 1567
rect 1761 1562 2598 1567
rect 2721 1562 2854 1567
rect 2881 1562 2958 1567
rect 3041 1562 3262 1567
rect 1177 1557 1294 1562
rect 417 1552 1110 1557
rect 1153 1552 1182 1557
rect 1289 1552 1910 1557
rect 1929 1552 2014 1557
rect 2033 1552 2142 1557
rect 2193 1552 2310 1557
rect 2321 1552 2414 1557
rect 2433 1552 2558 1557
rect 2713 1552 3198 1557
rect 1153 1547 1158 1552
rect 2321 1547 2326 1552
rect 393 1542 678 1547
rect 785 1542 910 1547
rect 953 1542 982 1547
rect 1041 1542 1158 1547
rect 1177 1542 1630 1547
rect 1681 1542 2230 1547
rect 2249 1542 2286 1547
rect 2297 1542 2326 1547
rect 2369 1542 2470 1547
rect 2513 1542 2574 1547
rect 2689 1542 2766 1547
rect 2785 1542 2862 1547
rect 2969 1542 3150 1547
rect 3385 1542 3406 1547
rect 113 1532 166 1537
rect 289 1532 382 1537
rect 561 1532 838 1537
rect 377 1527 566 1532
rect 977 1527 982 1542
rect 1073 1532 1102 1537
rect 1193 1532 1766 1537
rect 1889 1532 2638 1537
rect 1097 1527 1198 1532
rect 585 1522 654 1527
rect 697 1522 750 1527
rect 809 1522 830 1527
rect 977 1522 1054 1527
rect 1329 1522 1406 1527
rect 1513 1522 1646 1527
rect 1657 1522 2406 1527
rect 2481 1522 2510 1527
rect 2553 1522 2590 1527
rect 2689 1522 2694 1542
rect 2705 1532 2758 1537
rect 3081 1532 3118 1537
rect 3217 1532 3286 1537
rect 3217 1527 3222 1532
rect 2737 1522 3222 1527
rect 3281 1527 3286 1532
rect 3313 1532 3422 1537
rect 3313 1527 3318 1532
rect 3281 1522 3318 1527
rect 3337 1522 3406 1527
rect 233 1517 310 1522
rect 1217 1517 1310 1522
rect 2609 1517 2694 1522
rect 0 1512 238 1517
rect 305 1512 406 1517
rect 441 1512 502 1517
rect 513 1512 614 1517
rect 753 1512 862 1517
rect 1025 1512 1062 1517
rect 1089 1512 1118 1517
rect 1113 1507 1118 1512
rect 1193 1512 1222 1517
rect 1305 1512 1630 1517
rect 1897 1512 2342 1517
rect 2441 1512 2494 1517
rect 2513 1512 2614 1517
rect 2993 1512 3110 1517
rect 1193 1507 1198 1512
rect 1625 1507 1734 1512
rect 1897 1507 1902 1512
rect 2713 1507 2806 1512
rect 249 1502 294 1507
rect 361 1502 462 1507
rect 569 1502 718 1507
rect 1113 1502 1198 1507
rect 1249 1502 1278 1507
rect 1289 1502 1606 1507
rect 1729 1502 1902 1507
rect 1921 1502 2094 1507
rect 2113 1502 2718 1507
rect 2801 1502 2862 1507
rect 2881 1502 2958 1507
rect 3081 1502 3150 1507
rect 3233 1502 3270 1507
rect 3377 1502 3414 1507
rect 2881 1497 2886 1502
rect 177 1492 398 1497
rect 1217 1492 1278 1497
rect 1321 1492 1398 1497
rect 1473 1492 1710 1497
rect 1969 1492 2382 1497
rect 2449 1492 2886 1497
rect 2953 1497 2958 1502
rect 2953 1492 2982 1497
rect 3273 1492 3350 1497
rect 1865 1487 1950 1492
rect 0 1482 166 1487
rect 161 1477 166 1482
rect 473 1482 558 1487
rect 473 1477 478 1482
rect 161 1472 478 1477
rect 553 1477 558 1482
rect 641 1482 1054 1487
rect 1337 1482 1870 1487
rect 1945 1482 2142 1487
rect 2177 1482 3286 1487
rect 641 1477 646 1482
rect 553 1472 646 1477
rect 1425 1472 1526 1477
rect 1561 1472 1702 1477
rect 1881 1472 1918 1477
rect 1929 1472 2038 1477
rect 2057 1472 2990 1477
rect 3297 1472 3366 1477
rect 1769 1467 1862 1472
rect 2985 1467 2990 1472
rect 3081 1467 3302 1472
rect 689 1462 830 1467
rect 689 1457 694 1462
rect 145 1452 214 1457
rect 665 1452 694 1457
rect 825 1457 830 1462
rect 1073 1462 1166 1467
rect 1185 1462 1230 1467
rect 1249 1462 1358 1467
rect 1377 1462 1446 1467
rect 1625 1462 1774 1467
rect 1857 1462 2462 1467
rect 2473 1462 2606 1467
rect 2673 1462 2702 1467
rect 2793 1462 2966 1467
rect 2985 1462 3086 1467
rect 1073 1457 1078 1462
rect 825 1452 878 1457
rect 1009 1452 1078 1457
rect 1161 1457 1166 1462
rect 1249 1457 1254 1462
rect 1161 1452 1254 1457
rect 1353 1457 1358 1462
rect 2697 1457 2798 1462
rect 1353 1452 1382 1457
rect 1457 1452 1614 1457
rect 1785 1452 1854 1457
rect 1865 1452 1966 1457
rect 1985 1452 2078 1457
rect 2129 1452 2214 1457
rect 2257 1452 2334 1457
rect 2353 1452 2390 1457
rect 2409 1452 2494 1457
rect 2505 1452 2630 1457
rect 3105 1452 3142 1457
rect 3161 1452 3254 1457
rect 1377 1447 1462 1452
rect 1609 1447 1702 1452
rect 1785 1447 1790 1452
rect 2129 1447 2134 1452
rect 2625 1447 2630 1452
rect 2817 1447 3014 1452
rect 377 1442 654 1447
rect 713 1442 742 1447
rect 769 1442 814 1447
rect 1025 1442 1342 1447
rect 1697 1442 1790 1447
rect 1817 1442 2134 1447
rect 2153 1442 2182 1447
rect 2193 1442 2238 1447
rect 2289 1442 2310 1447
rect 2321 1442 2526 1447
rect 2625 1442 2710 1447
rect 2729 1442 2822 1447
rect 3009 1442 3038 1447
rect 3057 1442 3190 1447
rect 3265 1442 3334 1447
rect 649 1437 718 1442
rect 833 1437 942 1442
rect 2705 1437 2710 1442
rect 3185 1437 3270 1442
rect 233 1432 406 1437
rect 417 1432 446 1437
rect 753 1432 838 1437
rect 937 1432 966 1437
rect 1073 1432 1118 1437
rect 1161 1432 1310 1437
rect 1409 1432 1678 1437
rect 1809 1432 2550 1437
rect 2705 1432 2750 1437
rect 2833 1432 2974 1437
rect 3097 1432 3166 1437
rect 401 1427 406 1432
rect 753 1427 758 1432
rect 401 1422 430 1427
rect 657 1422 782 1427
rect 793 1422 950 1427
rect 1081 1422 1398 1427
rect 1521 1422 1630 1427
rect 1393 1417 1526 1422
rect 1625 1417 1630 1422
rect 1689 1422 1766 1427
rect 1913 1422 1950 1427
rect 1969 1422 2006 1427
rect 2033 1422 2318 1427
rect 2361 1422 2406 1427
rect 2417 1422 2486 1427
rect 2609 1422 2798 1427
rect 2881 1422 3294 1427
rect 3361 1422 3438 1427
rect 1689 1417 1694 1422
rect 481 1412 566 1417
rect 697 1412 1046 1417
rect 1105 1412 1326 1417
rect 1545 1412 1606 1417
rect 1625 1412 1694 1417
rect 1809 1412 1894 1417
rect 1921 1412 2190 1417
rect 2241 1412 2342 1417
rect 2353 1412 2910 1417
rect 3033 1412 3214 1417
rect 3241 1412 3270 1417
rect 137 1402 214 1407
rect 729 1402 806 1407
rect 841 1402 886 1407
rect 1137 1402 1222 1407
rect 1257 1402 1502 1407
rect 137 1397 142 1402
rect 113 1392 142 1397
rect 209 1397 214 1402
rect 209 1392 238 1397
rect 281 1392 310 1397
rect 537 1392 574 1397
rect 769 1392 846 1397
rect 881 1392 886 1402
rect 1553 1397 1670 1402
rect 1809 1397 1814 1412
rect 1889 1407 1894 1412
rect 2905 1407 3038 1412
rect 1889 1402 2886 1407
rect 3057 1402 3158 1407
rect 3265 1397 3270 1412
rect 913 1392 1014 1397
rect 1089 1392 1134 1397
rect 1153 1392 1246 1397
rect 1337 1392 1374 1397
rect 1457 1392 1558 1397
rect 1665 1392 1814 1397
rect 1841 1392 1966 1397
rect 2057 1392 2118 1397
rect 2153 1392 2358 1397
rect 2385 1392 2478 1397
rect 2497 1392 2606 1397
rect 2673 1392 2822 1397
rect 2857 1392 3054 1397
rect 3049 1387 3054 1392
rect 3137 1392 3182 1397
rect 3233 1392 3270 1397
rect 3137 1387 3142 1392
rect 441 1382 494 1387
rect 585 1382 662 1387
rect 833 1382 950 1387
rect 961 1382 1134 1387
rect 1241 1382 1478 1387
rect 1569 1382 1654 1387
rect 1809 1382 2078 1387
rect 2089 1382 2118 1387
rect 2153 1382 2174 1387
rect 2185 1382 2662 1387
rect 2753 1382 2902 1387
rect 3049 1382 3142 1387
rect 3161 1382 3198 1387
rect 3241 1382 3366 1387
rect 1129 1377 1246 1382
rect 2657 1377 2758 1382
rect 121 1372 278 1377
rect 417 1372 678 1377
rect 1073 1372 1110 1377
rect 1265 1372 1334 1377
rect 1457 1372 1590 1377
rect 1793 1372 2446 1377
rect 2465 1372 2550 1377
rect 2921 1372 3030 1377
rect 1265 1367 1270 1372
rect 2921 1367 2926 1372
rect 393 1362 742 1367
rect 969 1362 1070 1367
rect 1113 1362 1270 1367
rect 1281 1362 1390 1367
rect 1473 1362 1630 1367
rect 1865 1362 1966 1367
rect 1985 1362 2126 1367
rect 2137 1362 2182 1367
rect 2201 1362 2662 1367
rect 2729 1362 2758 1367
rect 2817 1362 2926 1367
rect 3025 1367 3030 1372
rect 3089 1367 3254 1372
rect 3025 1362 3054 1367
rect 3065 1362 3094 1367
rect 3249 1362 3406 1367
rect 425 1352 518 1357
rect 585 1352 646 1357
rect 673 1352 758 1357
rect 937 1352 998 1357
rect 1009 1352 1102 1357
rect 1145 1352 1174 1357
rect 1241 1352 1534 1357
rect 1553 1352 1718 1357
rect 1801 1352 2494 1357
rect 2929 1352 3238 1357
rect 673 1347 678 1352
rect 2489 1347 2630 1352
rect 113 1342 238 1347
rect 273 1342 326 1347
rect 409 1342 582 1347
rect 625 1342 678 1347
rect 689 1342 710 1347
rect 849 1342 902 1347
rect 921 1342 950 1347
rect 961 1342 1094 1347
rect 1153 1342 1190 1347
rect 1225 1342 1246 1347
rect 1313 1342 1614 1347
rect 1809 1342 2142 1347
rect 2169 1342 2222 1347
rect 2249 1342 2358 1347
rect 2441 1342 2470 1347
rect 2625 1342 2814 1347
rect 2873 1342 2958 1347
rect 3145 1342 3374 1347
rect 3409 1342 3454 1347
rect 2353 1337 2358 1342
rect 2465 1337 2470 1342
rect 377 1332 478 1337
rect 521 1332 550 1337
rect 569 1332 622 1337
rect 633 1332 726 1337
rect 753 1332 838 1337
rect 545 1327 550 1332
rect 385 1322 438 1327
rect 545 1322 694 1327
rect 225 1312 422 1317
rect 513 1312 702 1317
rect 721 1307 726 1332
rect 833 1327 838 1332
rect 929 1332 1414 1337
rect 1521 1332 1670 1337
rect 1801 1332 1870 1337
rect 1897 1332 2030 1337
rect 2097 1332 2206 1337
rect 2353 1332 2446 1337
rect 2465 1332 2670 1337
rect 2985 1332 3302 1337
rect 929 1327 934 1332
rect 1665 1327 1670 1332
rect 2225 1327 2334 1332
rect 745 1322 798 1327
rect 833 1322 934 1327
rect 953 1322 1022 1327
rect 777 1312 814 1317
rect 449 1302 574 1307
rect 649 1302 726 1307
rect 769 1302 1006 1307
rect 1057 1302 1062 1327
rect 1177 1322 1214 1327
rect 1233 1322 1286 1327
rect 1417 1322 1646 1327
rect 1665 1322 1926 1327
rect 1945 1322 2230 1327
rect 2329 1322 2606 1327
rect 2697 1322 2758 1327
rect 2801 1322 2934 1327
rect 3153 1322 3190 1327
rect 1233 1317 1238 1322
rect 1169 1312 1238 1317
rect 1297 1312 1382 1317
rect 1489 1312 1686 1317
rect 1857 1312 2494 1317
rect 2529 1312 2590 1317
rect 2625 1312 2718 1317
rect 3017 1312 3294 1317
rect 3321 1312 3350 1317
rect 2529 1307 2534 1312
rect 2713 1307 2870 1312
rect 3017 1307 3022 1312
rect 1129 1302 1806 1307
rect 1865 1302 1894 1307
rect 1961 1302 2014 1307
rect 2097 1302 2326 1307
rect 2385 1302 2534 1307
rect 2553 1302 2694 1307
rect 2865 1302 3022 1307
rect 3217 1297 3350 1302
rect 617 1292 726 1297
rect 1065 1292 1702 1297
rect 1793 1292 2358 1297
rect 2457 1292 2542 1297
rect 2561 1292 2846 1297
rect 3041 1292 3166 1297
rect 3193 1292 3222 1297
rect 3345 1292 3414 1297
rect 417 1287 598 1292
rect 393 1282 422 1287
rect 593 1282 654 1287
rect 737 1282 846 1287
rect 881 1282 918 1287
rect 1137 1282 1310 1287
rect 1385 1282 1430 1287
rect 1529 1282 1646 1287
rect 1817 1282 1886 1287
rect 1897 1282 1966 1287
rect 1977 1282 2086 1287
rect 2097 1282 2198 1287
rect 2249 1282 2302 1287
rect 2313 1282 2598 1287
rect 2785 1282 2822 1287
rect 3169 1282 3334 1287
rect 649 1277 742 1282
rect 1665 1277 1798 1282
rect 2617 1277 2734 1282
rect 449 1272 534 1277
rect 553 1272 630 1277
rect 921 1272 1046 1277
rect 1129 1272 1294 1277
rect 1617 1272 1670 1277
rect 1793 1272 2454 1277
rect 2505 1272 2566 1277
rect 2585 1272 2622 1277
rect 2729 1272 3294 1277
rect 1041 1267 1046 1272
rect 1313 1267 1542 1272
rect 1617 1267 1622 1272
rect 409 1262 486 1267
rect 561 1262 894 1267
rect 1041 1262 1214 1267
rect 1257 1262 1318 1267
rect 1537 1262 1622 1267
rect 1665 1262 2206 1267
rect 2281 1262 2342 1267
rect 2409 1262 2718 1267
rect 2825 1262 2886 1267
rect 3097 1262 3190 1267
rect 889 1257 1030 1262
rect 2713 1257 2830 1262
rect 257 1252 462 1257
rect 545 1252 606 1257
rect 1025 1252 1070 1257
rect 1065 1247 1070 1252
rect 1145 1252 1526 1257
rect 1777 1252 2614 1257
rect 2665 1252 2694 1257
rect 1145 1247 1150 1252
rect 2689 1247 2694 1252
rect 2921 1252 3022 1257
rect 3041 1252 3094 1257
rect 2921 1247 2926 1252
rect 425 1242 470 1247
rect 481 1242 542 1247
rect 721 1242 774 1247
rect 785 1242 822 1247
rect 873 1242 934 1247
rect 1065 1242 1150 1247
rect 1177 1242 1214 1247
rect 1289 1242 1486 1247
rect 1625 1242 1758 1247
rect 1881 1242 2334 1247
rect 2345 1242 2542 1247
rect 2689 1242 2926 1247
rect 3017 1247 3022 1252
rect 3017 1242 3222 1247
rect 3241 1242 3326 1247
rect 561 1237 702 1242
rect 1625 1237 1630 1242
rect 329 1232 566 1237
rect 697 1232 750 1237
rect 905 1232 1030 1237
rect 1169 1232 1198 1237
rect 1353 1232 1406 1237
rect 1457 1232 1630 1237
rect 1753 1237 1758 1242
rect 3217 1237 3222 1242
rect 1753 1232 1838 1237
rect 1929 1232 1974 1237
rect 2009 1232 2038 1237
rect 2081 1232 2710 1237
rect 2769 1232 2846 1237
rect 2937 1232 3206 1237
rect 3217 1232 3262 1237
rect 1217 1227 1334 1232
rect 2081 1227 2086 1232
rect 2705 1227 2710 1232
rect 3257 1227 3262 1232
rect 3337 1232 3414 1237
rect 3337 1227 3342 1232
rect 305 1222 358 1227
rect 449 1222 478 1227
rect 577 1222 670 1227
rect 473 1217 582 1222
rect 665 1217 670 1222
rect 729 1222 758 1227
rect 801 1222 910 1227
rect 1145 1222 1222 1227
rect 1329 1222 1382 1227
rect 1577 1222 1926 1227
rect 1977 1222 2086 1227
rect 2153 1222 2350 1227
rect 2457 1222 2518 1227
rect 2529 1222 2582 1227
rect 2705 1222 2982 1227
rect 3257 1222 3342 1227
rect 729 1217 734 1222
rect 1401 1217 1526 1222
rect 2529 1217 2534 1222
rect 3057 1217 3158 1222
rect 601 1212 646 1217
rect 665 1212 734 1217
rect 1081 1212 1254 1217
rect 1273 1212 1406 1217
rect 1521 1212 2534 1217
rect 3033 1212 3062 1217
rect 3153 1212 3182 1217
rect 1249 1207 1254 1212
rect 2753 1207 2830 1212
rect 2889 1207 3014 1212
rect 217 1202 286 1207
rect 457 1202 502 1207
rect 569 1202 614 1207
rect 1153 1202 1230 1207
rect 1249 1202 1510 1207
rect 1601 1202 1902 1207
rect 1921 1202 2030 1207
rect 2105 1202 2134 1207
rect 2225 1202 2406 1207
rect 2657 1202 2678 1207
rect 2729 1202 2758 1207
rect 2825 1202 2894 1207
rect 3009 1202 3238 1207
rect 217 1197 222 1202
rect 145 1192 182 1197
rect 193 1192 222 1197
rect 281 1197 286 1202
rect 1505 1197 1606 1202
rect 2425 1197 2638 1202
rect 281 1192 806 1197
rect 825 1192 950 1197
rect 985 1192 1086 1197
rect 1153 1192 1182 1197
rect 1193 1192 1318 1197
rect 1401 1192 1486 1197
rect 1625 1192 1990 1197
rect 2009 1192 2430 1197
rect 2633 1192 2814 1197
rect 177 1187 182 1192
rect 801 1187 806 1192
rect 177 1182 262 1187
rect 433 1182 470 1187
rect 545 1182 582 1187
rect 601 1182 678 1187
rect 801 1182 822 1187
rect 97 1172 166 1177
rect 161 1167 166 1172
rect 273 1172 342 1177
rect 553 1172 662 1177
rect 801 1172 822 1177
rect 273 1167 278 1172
rect 161 1162 278 1167
rect 633 1162 750 1167
rect 777 1162 806 1167
rect 649 1152 782 1157
rect 97 1142 214 1147
rect 337 1142 462 1147
rect 481 1142 526 1147
rect 537 1142 622 1147
rect 641 1142 686 1147
rect 337 1137 342 1142
rect 313 1132 342 1137
rect 457 1137 462 1142
rect 457 1132 766 1137
rect 817 1127 822 1172
rect 849 1147 854 1192
rect 1985 1187 1990 1192
rect 2809 1187 2814 1192
rect 2905 1192 3286 1197
rect 3329 1192 3366 1197
rect 2905 1187 2910 1192
rect 945 1182 1582 1187
rect 1737 1182 1894 1187
rect 1985 1182 2118 1187
rect 2153 1182 2174 1187
rect 2193 1182 2790 1187
rect 2809 1182 2910 1187
rect 2985 1182 3070 1187
rect 3121 1182 3166 1187
rect 3217 1182 3286 1187
rect 873 1172 990 1177
rect 1001 1172 1046 1177
rect 1233 1172 1398 1177
rect 1433 1172 1630 1177
rect 1713 1172 1958 1177
rect 1985 1172 2086 1177
rect 2097 1172 2782 1177
rect 2929 1172 3086 1177
rect 1065 1167 1214 1172
rect 3281 1167 3350 1172
rect 881 1162 902 1167
rect 953 1162 1022 1167
rect 1041 1162 1070 1167
rect 1209 1162 1374 1167
rect 1449 1162 1518 1167
rect 1665 1162 1774 1167
rect 1897 1162 2054 1167
rect 2073 1162 2214 1167
rect 2321 1162 2422 1167
rect 2489 1162 3286 1167
rect 3345 1162 3374 1167
rect 1537 1157 1646 1162
rect 1049 1152 1094 1157
rect 1153 1152 1542 1157
rect 1641 1152 1798 1157
rect 2009 1152 2118 1157
rect 2129 1152 2270 1157
rect 2353 1152 2382 1157
rect 2417 1152 2638 1157
rect 2681 1152 2766 1157
rect 2961 1152 3014 1157
rect 3033 1152 3110 1157
rect 3297 1152 3422 1157
rect 1841 1147 1990 1152
rect 2849 1147 2942 1152
rect 833 1142 854 1147
rect 897 1142 1022 1147
rect 1081 1142 1174 1147
rect 1209 1142 1270 1147
rect 1425 1142 1678 1147
rect 1817 1142 1846 1147
rect 1985 1142 2094 1147
rect 2177 1142 2198 1147
rect 2233 1142 2854 1147
rect 2937 1142 3094 1147
rect 1169 1137 1174 1142
rect 1289 1137 1406 1142
rect 961 1132 1006 1137
rect 1169 1132 1294 1137
rect 1401 1132 1974 1137
rect 2073 1132 2574 1137
rect 2689 1132 2758 1137
rect 2865 1132 2942 1137
rect 3105 1132 3334 1137
rect 161 1122 294 1127
rect 393 1122 494 1127
rect 609 1122 654 1127
rect 769 1122 822 1127
rect 841 1122 942 1127
rect 961 1122 966 1132
rect 2753 1127 2870 1132
rect 2937 1127 3110 1132
rect 985 1122 1366 1127
rect 1377 1122 1662 1127
rect 1865 1122 1918 1127
rect 2001 1122 2134 1127
rect 2337 1122 2454 1127
rect 2673 1122 2734 1127
rect 2889 1122 2918 1127
rect 3313 1122 3390 1127
rect 161 1117 166 1122
rect 289 1117 374 1122
rect 841 1117 846 1122
rect 73 1112 166 1117
rect 369 1112 670 1117
rect 777 1112 846 1117
rect 937 1117 942 1122
rect 1361 1117 1366 1122
rect 2153 1117 2254 1122
rect 937 1112 1046 1117
rect 1137 1112 1310 1117
rect 1361 1112 2158 1117
rect 2249 1112 2278 1117
rect 2409 1112 2502 1117
rect 2625 1112 2726 1117
rect 2769 1112 2902 1117
rect 2929 1112 3046 1117
rect 3065 1112 3126 1117
rect 2297 1107 2390 1112
rect 177 1102 1086 1107
rect 1161 1102 1182 1107
rect 1193 1102 1222 1107
rect 1233 1102 1278 1107
rect 1377 1102 1470 1107
rect 1489 1102 1566 1107
rect 1601 1102 1654 1107
rect 1897 1102 2302 1107
rect 2385 1102 2614 1107
rect 2705 1102 2742 1107
rect 2801 1102 2838 1107
rect 2857 1102 3014 1107
rect 177 1097 182 1102
rect 1649 1097 1654 1102
rect 2833 1097 2838 1102
rect 0 1092 182 1097
rect 193 1092 758 1097
rect 937 1092 998 1097
rect 1049 1092 1094 1097
rect 1177 1092 1262 1097
rect 1273 1092 1422 1097
rect 1433 1092 1614 1097
rect 1649 1092 1774 1097
rect 1833 1092 1918 1097
rect 2009 1092 2086 1097
rect 2185 1092 2262 1097
rect 2289 1092 2422 1097
rect 2441 1092 2822 1097
rect 2833 1092 2918 1097
rect 3177 1092 3294 1097
rect 793 1087 918 1092
rect 2081 1087 2190 1092
rect 2817 1087 2822 1092
rect 377 1082 422 1087
rect 449 1082 630 1087
rect 689 1082 798 1087
rect 913 1082 942 1087
rect 1153 1082 1318 1087
rect 1337 1082 1454 1087
rect 1497 1082 1526 1087
rect 1561 1082 1590 1087
rect 1793 1082 1902 1087
rect 1945 1082 1982 1087
rect 2017 1082 2062 1087
rect 2209 1082 2270 1087
rect 2625 1082 2774 1087
rect 2817 1082 2942 1087
rect 121 1077 270 1082
rect 449 1077 454 1082
rect 625 1077 630 1082
rect 961 1077 1094 1082
rect 1609 1077 1774 1082
rect 2425 1077 2606 1082
rect 0 1072 126 1077
rect 265 1072 454 1077
rect 521 1072 614 1077
rect 625 1072 966 1077
rect 1089 1072 1118 1077
rect 1145 1072 1390 1077
rect 1441 1072 1614 1077
rect 1769 1072 1822 1077
rect 2001 1072 2182 1077
rect 2265 1072 2302 1077
rect 2401 1072 2430 1077
rect 2601 1072 2894 1077
rect 1441 1067 1446 1072
rect 1841 1067 1982 1072
rect 137 1062 254 1067
rect 649 1062 950 1067
rect 985 1062 1446 1067
rect 1513 1062 1742 1067
rect 1785 1062 1846 1067
rect 1977 1062 2790 1067
rect 2809 1062 2998 1067
rect 369 1057 614 1062
rect 193 1052 374 1057
rect 609 1052 638 1057
rect 745 1052 790 1057
rect 1009 1052 1110 1057
rect 1153 1052 1294 1057
rect 817 1047 910 1052
rect 0 1042 686 1047
rect 793 1042 822 1047
rect 905 1042 934 1047
rect 1153 1042 1158 1052
rect 1377 1047 1382 1057
rect 1441 1052 1534 1057
rect 1553 1052 1654 1057
rect 1753 1052 2462 1057
rect 2577 1052 2670 1057
rect 2713 1052 3038 1057
rect 1209 1042 1334 1047
rect 1377 1042 1422 1047
rect 1433 1042 1590 1047
rect 1753 1042 2062 1047
rect 2097 1042 2134 1047
rect 2145 1042 2430 1047
rect 2641 1042 2766 1047
rect 2793 1042 3214 1047
rect 1001 1037 1158 1042
rect 2449 1037 2622 1042
rect 193 1032 1006 1037
rect 1193 1032 1254 1037
rect 1353 1032 1662 1037
rect 1761 1032 2454 1037
rect 2617 1032 3014 1037
rect 3049 1032 3094 1037
rect 3193 1032 3374 1037
rect 193 1027 198 1032
rect 0 1022 198 1027
rect 241 1022 286 1027
rect 305 1022 366 1027
rect 441 1022 470 1027
rect 761 1022 782 1027
rect 793 1022 822 1027
rect 905 1022 934 1027
rect 1017 1022 1046 1027
rect 1073 1022 1838 1027
rect 1849 1022 2438 1027
rect 2497 1022 2702 1027
rect 2721 1022 2750 1027
rect 2777 1022 2854 1027
rect 2881 1022 3086 1027
rect 3185 1022 3214 1027
rect 817 1017 910 1022
rect 1041 1017 1046 1022
rect 2721 1017 2726 1022
rect 3209 1017 3214 1022
rect 3273 1022 3422 1027
rect 3273 1017 3278 1022
rect 161 1012 334 1017
rect 465 1012 550 1017
rect 569 1012 638 1017
rect 1041 1012 1062 1017
rect 1097 1012 1238 1017
rect 1313 1012 1734 1017
rect 1897 1012 2038 1017
rect 2089 1012 2166 1017
rect 2257 1012 2502 1017
rect 2513 1012 2726 1017
rect 2777 1012 3046 1017
rect 3209 1012 3278 1017
rect 3297 1012 3326 1017
rect 569 1007 574 1012
rect 0 1002 86 1007
rect 113 1002 150 1007
rect 225 1002 262 1007
rect 321 1002 366 1007
rect 385 1002 486 1007
rect 513 1002 574 1007
rect 633 1007 638 1012
rect 1057 1007 1062 1012
rect 1753 1007 1854 1012
rect 633 1002 662 1007
rect 769 1002 878 1007
rect 897 1002 982 1007
rect 1057 1002 1758 1007
rect 1849 1002 1886 1007
rect 1953 1002 2134 1007
rect 2193 1002 2302 1007
rect 81 987 86 1002
rect 1881 997 1958 1002
rect 2129 997 2134 1002
rect 2497 997 2502 1012
rect 2601 1002 2638 1007
rect 2649 1002 3150 1007
rect 3281 997 3350 1002
rect 97 992 174 997
rect 209 992 294 997
rect 337 992 382 997
rect 449 992 582 997
rect 593 992 678 997
rect 713 992 782 997
rect 889 992 934 997
rect 1121 992 1222 997
rect 1265 992 1302 997
rect 1313 992 1334 997
rect 1353 992 1414 997
rect 1433 992 1662 997
rect 1713 992 1838 997
rect 1977 992 2022 997
rect 2073 992 2118 997
rect 2129 992 2214 997
rect 2273 992 2318 997
rect 2337 992 2478 997
rect 2497 992 2598 997
rect 2641 992 2822 997
rect 2833 992 2902 997
rect 2929 992 2998 997
rect 3153 992 3286 997
rect 3345 992 3446 997
rect 953 987 1046 992
rect 0 982 70 987
rect 81 982 958 987
rect 1041 982 1070 987
rect 1121 982 1158 987
rect 1169 982 1390 987
rect 65 977 70 982
rect 1409 977 1414 992
rect 2337 987 2342 992
rect 1449 982 1606 987
rect 1649 982 1686 987
rect 1777 982 1814 987
rect 1873 982 2342 987
rect 2473 987 2478 992
rect 2473 982 2934 987
rect 2985 982 3054 987
rect 3121 982 3214 987
rect 3297 982 3334 987
rect 1681 977 1782 982
rect 1873 977 1878 982
rect 2361 977 2446 982
rect 65 972 1046 977
rect 1129 972 1382 977
rect 1409 972 1662 977
rect 1801 972 1878 977
rect 1889 972 2094 977
rect 2129 972 2190 977
rect 2289 972 2366 977
rect 2441 972 2518 977
rect 2561 972 2622 977
rect 2697 972 2750 977
rect 2873 972 2942 977
rect 3033 972 3238 977
rect 0 962 30 967
rect 273 962 774 967
rect 889 962 918 967
rect 1049 962 1718 967
rect 1777 962 2006 967
rect 2033 962 2254 967
rect 2281 962 2430 967
rect 25 957 278 962
rect 769 957 894 962
rect 2513 957 2518 972
rect 2601 962 3054 967
rect 3193 962 3222 967
rect 3337 962 3414 967
rect 3049 957 3198 962
rect 297 952 438 957
rect 449 952 558 957
rect 673 952 750 957
rect 1025 952 1230 957
rect 1337 952 1558 957
rect 1673 952 1870 957
rect 1929 952 2502 957
rect 2513 952 2862 957
rect 2905 952 3030 957
rect 1553 947 1678 952
rect 2497 947 2502 952
rect 0 942 78 947
rect 89 942 214 947
rect 305 942 374 947
rect 401 942 494 947
rect 529 942 590 947
rect 817 942 926 947
rect 1017 942 1062 947
rect 1081 942 1142 947
rect 1193 942 1334 947
rect 1417 942 1478 947
rect 1489 942 1526 947
rect 1697 942 1734 947
rect 1889 942 1958 947
rect 2001 942 2174 947
rect 2265 942 2390 947
rect 2401 942 2454 947
rect 2497 942 2590 947
rect 2665 942 3358 947
rect 529 937 534 942
rect 817 937 822 942
rect 353 932 534 937
rect 681 932 822 937
rect 921 937 926 942
rect 921 932 1046 937
rect 1057 932 1062 942
rect 2385 937 2390 942
rect 1313 932 1430 937
rect 1481 932 1574 937
rect 1593 932 1926 937
rect 2025 932 2134 937
rect 2177 932 2254 937
rect 2385 932 2550 937
rect 2713 932 2822 937
rect 2929 932 2982 937
rect 3017 932 3070 937
rect 1057 927 1294 932
rect 2249 927 2374 932
rect 2569 927 2654 932
rect 2929 927 2934 932
rect 0 922 30 927
rect 25 917 30 922
rect 209 922 678 927
rect 833 922 998 927
rect 1289 922 1526 927
rect 1577 922 1622 927
rect 1745 922 2198 927
rect 2369 922 2574 927
rect 2649 922 2742 927
rect 209 917 214 922
rect 673 917 678 922
rect 25 912 214 917
rect 345 912 374 917
rect 409 912 478 917
rect 673 912 710 917
rect 1105 912 1190 917
rect 1201 912 1286 917
rect 1297 912 1510 917
rect 1521 907 1526 922
rect 1537 912 1686 917
rect 1753 912 2094 917
rect 2297 912 2342 917
rect 2409 912 2454 917
rect 2561 912 2638 917
rect 2737 912 2742 922
rect 2849 922 2934 927
rect 2985 922 3046 927
rect 3089 922 3182 927
rect 3241 922 3358 927
rect 2849 917 2854 922
rect 3241 917 3246 922
rect 2785 912 2830 917
rect 2849 912 2878 917
rect 2897 912 2942 917
rect 2977 912 3014 917
rect 3217 912 3246 917
rect 3353 917 3358 922
rect 3353 912 3438 917
rect 377 902 838 907
rect 937 902 1022 907
rect 1113 902 1134 907
rect 1241 902 1510 907
rect 1521 902 1814 907
rect 1825 902 1886 907
rect 1929 902 2006 907
rect 2097 902 2150 907
rect 2721 902 3126 907
rect 3225 902 3366 907
rect 1505 897 1510 902
rect 2249 897 2486 902
rect 2721 897 2726 902
rect 233 892 334 897
rect 329 887 334 892
rect 417 892 446 897
rect 1009 892 1278 897
rect 1401 892 1438 897
rect 1505 892 1758 897
rect 1769 892 1806 897
rect 1833 892 2254 897
rect 2481 892 2726 897
rect 2737 892 3070 897
rect 3161 892 3190 897
rect 3241 892 3334 897
rect 417 887 422 892
rect 3065 887 3166 892
rect 3329 887 3334 892
rect 3401 892 3430 897
rect 3401 887 3406 892
rect 185 882 246 887
rect 329 882 422 887
rect 457 882 686 887
rect 1065 882 1214 887
rect 1345 882 1494 887
rect 1521 882 2526 887
rect 2625 882 3046 887
rect 3329 882 3406 887
rect 1209 877 1302 882
rect 2521 877 2630 882
rect 761 872 782 877
rect 921 872 950 877
rect 1113 872 1190 877
rect 1297 872 1822 877
rect 1849 872 2206 877
rect 2241 872 2502 877
rect 2649 872 3142 877
rect 3137 867 3142 872
rect 3281 872 3310 877
rect 3281 867 3286 872
rect 465 862 534 867
rect 553 862 718 867
rect 1089 862 1150 867
rect 1169 862 1262 867
rect 1385 862 1454 867
rect 1473 862 1542 867
rect 1585 862 1622 867
rect 1633 862 1662 867
rect 1777 862 1838 867
rect 1953 862 3038 867
rect 3137 862 3286 867
rect 553 857 558 862
rect 409 852 558 857
rect 713 857 718 862
rect 1473 857 1478 862
rect 713 852 790 857
rect 897 852 990 857
rect 1105 852 1398 857
rect 1417 852 1478 857
rect 1489 852 1710 857
rect 1857 852 2070 857
rect 2081 852 2246 857
rect 2305 852 2566 857
rect 2657 852 2734 857
rect 2793 852 2950 857
rect 577 847 694 852
rect 1489 847 1494 852
rect 313 842 398 847
rect 521 842 582 847
rect 689 842 774 847
rect 1065 842 1494 847
rect 1513 842 1742 847
rect 1825 842 2238 847
rect 2249 842 2550 847
rect 2633 842 2678 847
rect 2801 842 2902 847
rect 2961 842 3118 847
rect 153 832 278 837
rect 577 832 686 837
rect 153 827 158 832
rect 121 822 158 827
rect 273 827 278 832
rect 681 827 686 832
rect 769 832 1054 837
rect 1177 832 1294 837
rect 1337 832 1446 837
rect 1481 832 1534 837
rect 1545 832 1654 837
rect 1689 832 1766 837
rect 1833 832 1998 837
rect 2209 832 2342 837
rect 2385 832 2462 837
rect 2529 832 2790 837
rect 2865 832 2926 837
rect 3065 832 3222 837
rect 3289 832 3374 837
rect 769 827 774 832
rect 2017 827 2190 832
rect 2785 827 2790 832
rect 2945 827 3070 832
rect 273 822 302 827
rect 353 822 382 827
rect 513 822 574 827
rect 609 822 662 827
rect 681 822 774 827
rect 793 822 886 827
rect 1217 822 1374 827
rect 1425 822 1582 827
rect 1593 822 1638 827
rect 1745 822 2022 827
rect 2185 822 2454 827
rect 2465 822 2622 827
rect 2713 822 2742 827
rect 2785 822 2950 827
rect 3089 822 3166 827
rect 3201 822 3398 827
rect 2449 817 2454 822
rect 3089 817 3094 822
rect 169 812 414 817
rect 537 812 606 817
rect 1033 812 1862 817
rect 1881 812 2230 817
rect 2329 812 2422 817
rect 2449 812 2582 817
rect 2601 812 3094 817
rect 3105 812 3246 817
rect 2417 807 2422 812
rect 289 802 326 807
rect 665 802 726 807
rect 953 802 1030 807
rect 1233 802 1358 807
rect 1377 802 1798 807
rect 1817 802 1926 807
rect 1937 802 1998 807
rect 2201 802 2310 807
rect 2337 802 2374 807
rect 2417 802 2486 807
rect 2569 802 2734 807
rect 2753 802 2798 807
rect 2913 802 2974 807
rect 1377 797 1382 802
rect 305 792 438 797
rect 745 792 910 797
rect 969 792 1062 797
rect 1337 792 1382 797
rect 1393 792 1414 797
rect 1457 792 1566 797
rect 1601 792 1662 797
rect 1713 792 1766 797
rect 1793 787 1798 802
rect 2081 797 2182 802
rect 2753 797 2758 802
rect 1833 792 1862 797
rect 1945 792 1966 797
rect 2057 792 2086 797
rect 2177 792 2758 797
rect 2769 792 2846 797
rect 2937 792 3014 797
rect 3129 792 3230 797
rect 3281 792 3326 797
rect 249 782 406 787
rect 457 782 646 787
rect 697 782 838 787
rect 1369 782 1718 787
rect 1793 782 2158 787
rect 2217 782 3086 787
rect 3297 782 3318 787
rect 457 777 462 782
rect 281 772 462 777
rect 641 777 646 782
rect 641 772 702 777
rect 921 772 1094 777
rect 1113 772 1198 777
rect 1249 772 1366 777
rect 1385 772 1470 777
rect 1505 772 1638 777
rect 1649 772 1726 777
rect 1801 772 2502 777
rect 2641 772 3014 777
rect 3097 772 3278 777
rect 513 767 614 772
rect 729 767 798 772
rect 921 767 926 772
rect 313 762 342 767
rect 473 762 518 767
rect 609 762 638 767
rect 705 762 734 767
rect 793 762 926 767
rect 1089 767 1094 772
rect 1649 767 1654 772
rect 2497 767 2630 772
rect 3009 767 3102 772
rect 1089 762 1550 767
rect 1561 762 1654 767
rect 1833 762 1926 767
rect 2001 762 2086 767
rect 2121 762 2246 767
rect 2353 762 2438 767
rect 2625 762 2758 767
rect 337 757 478 762
rect 2785 757 2990 762
rect 529 752 614 757
rect 705 752 782 757
rect 937 752 1046 757
rect 1089 752 1118 757
rect 1129 752 1206 757
rect 1217 752 1246 757
rect 1265 752 1334 757
rect 1369 752 1430 757
rect 1449 752 1558 757
rect 1617 752 1646 757
rect 1681 752 1750 757
rect 1937 752 2790 757
rect 2985 752 3046 757
rect 1873 747 1942 752
rect 385 742 582 747
rect 729 742 1302 747
rect 1313 742 1342 747
rect 1353 742 1438 747
rect 1449 742 1702 747
rect 1873 737 1878 747
rect 2025 742 2718 747
rect 2713 737 2718 742
rect 2801 742 2990 747
rect 3113 742 3182 747
rect 3217 742 3350 747
rect 2801 737 2806 742
rect 3217 737 3222 742
rect 153 732 222 737
rect 481 732 678 737
rect 689 732 822 737
rect 1153 732 1174 737
rect 1321 732 1502 737
rect 1537 732 1630 737
rect 1657 732 1710 737
rect 1761 732 1790 737
rect 1825 732 1878 737
rect 1889 732 2022 737
rect 2065 732 2230 737
rect 2297 732 2366 737
rect 2417 732 2494 737
rect 2569 732 2614 737
rect 2625 732 2694 737
rect 2713 732 2806 737
rect 2825 732 3054 737
rect 3145 732 3222 737
rect 3345 737 3350 742
rect 3345 732 3414 737
rect 673 727 678 732
rect 1033 727 1134 732
rect 1193 727 1302 732
rect 2625 727 2630 732
rect 81 722 182 727
rect 337 722 462 727
rect 489 722 550 727
rect 577 722 606 727
rect 673 722 854 727
rect 873 722 1038 727
rect 1129 722 1198 727
rect 1297 722 2086 727
rect 2097 722 2150 727
rect 2177 722 2630 727
rect 2929 722 2950 727
rect 3233 722 3302 727
rect 337 717 342 722
rect 89 712 198 717
rect 209 712 254 717
rect 265 712 342 717
rect 457 717 462 722
rect 457 712 518 717
rect 513 707 518 712
rect 593 712 622 717
rect 769 712 798 717
rect 593 707 598 712
rect 353 702 454 707
rect 513 702 598 707
rect 793 697 798 712
rect 953 712 982 717
rect 1049 712 2198 717
rect 2217 712 2534 717
rect 2561 712 2598 717
rect 2769 712 2878 717
rect 2977 712 3046 717
rect 3089 712 3222 717
rect 3289 712 3342 717
rect 953 697 958 712
rect 2529 707 2534 712
rect 1041 702 1070 707
rect 1097 702 1398 707
rect 1489 702 1534 707
rect 1633 702 1718 707
rect 1841 702 1902 707
rect 1929 702 2142 707
rect 2321 702 2454 707
rect 2465 702 2518 707
rect 2529 702 2662 707
rect 2673 702 2822 707
rect 2833 702 2974 707
rect 2209 697 2302 702
rect 2465 697 2470 702
rect 2833 697 2838 702
rect 65 692 94 697
rect 89 687 94 692
rect 465 692 494 697
rect 793 692 958 697
rect 1121 692 1166 697
rect 1201 692 1246 697
rect 1265 692 1294 697
rect 1337 692 1518 697
rect 1529 692 1550 697
rect 1561 692 1622 697
rect 1729 692 2118 697
rect 2185 692 2214 697
rect 2297 692 2470 697
rect 2481 692 2838 697
rect 2969 697 2974 702
rect 3057 702 3086 707
rect 3161 702 3214 707
rect 3273 702 3318 707
rect 3057 697 3062 702
rect 2969 692 3062 697
rect 3201 692 3454 697
rect 89 682 342 687
rect 337 677 342 682
rect 465 677 470 692
rect 1265 687 1270 692
rect 1153 682 1190 687
rect 1217 682 1270 687
rect 1281 682 1446 687
rect 1497 682 1534 687
rect 1553 682 1814 687
rect 1833 682 1870 687
rect 1905 682 2886 687
rect 1553 677 1558 682
rect 337 672 470 677
rect 1057 672 1558 677
rect 1625 672 1838 677
rect 1945 672 2158 677
rect 2337 672 2406 677
rect 2417 672 2718 677
rect 2881 672 2950 677
rect 2177 667 2318 672
rect 777 662 966 667
rect 1129 662 1150 667
rect 1225 662 1582 667
rect 1593 662 1942 667
rect 1985 662 2182 667
rect 2313 662 2958 667
rect 777 647 782 662
rect 961 647 966 662
rect 1985 657 1990 662
rect 1321 652 1398 657
rect 1489 652 1678 657
rect 1713 652 1766 657
rect 1809 652 1870 657
rect 1921 652 1990 657
rect 2073 652 2310 657
rect 2321 652 2710 657
rect 2785 652 2838 657
rect 753 642 782 647
rect 833 642 942 647
rect 961 642 990 647
rect 1313 642 1862 647
rect 1873 642 1958 647
rect 1985 642 2182 647
rect 2353 642 2606 647
rect 2633 642 2686 647
rect 833 637 838 642
rect 689 632 838 637
rect 937 637 942 642
rect 1873 637 1878 642
rect 937 632 998 637
rect 1145 632 1174 637
rect 1249 632 1286 637
rect 1377 632 1606 637
rect 1617 632 1646 637
rect 1745 632 1878 637
rect 1969 632 2254 637
rect 2297 632 2350 637
rect 2361 632 2726 637
rect 2857 632 2998 637
rect 3137 632 3206 637
rect 1617 627 1622 632
rect 3137 627 3142 632
rect 217 622 342 627
rect 705 622 766 627
rect 849 622 926 627
rect 1033 622 1062 627
rect 1113 622 1622 627
rect 1801 622 1854 627
rect 1881 622 2046 627
rect 2169 622 2262 627
rect 2313 622 2414 627
rect 2425 622 2574 627
rect 2601 622 2694 627
rect 2721 622 2790 627
rect 2801 622 2918 627
rect 3113 622 3142 627
rect 3201 627 3206 632
rect 3377 627 3382 637
rect 3201 622 3230 627
rect 3265 622 3422 627
rect 217 617 222 622
rect 121 612 222 617
rect 337 617 342 622
rect 921 617 1038 622
rect 2721 617 2726 622
rect 2937 617 3094 622
rect 3265 617 3270 622
rect 337 612 366 617
rect 465 612 558 617
rect 745 612 862 617
rect 1121 612 1158 617
rect 1273 612 1566 617
rect 1593 612 1622 617
rect 1673 612 1766 617
rect 1817 612 1846 617
rect 1857 612 1910 617
rect 1953 612 2086 617
rect 2097 612 2190 617
rect 2273 612 2726 617
rect 2793 612 2942 617
rect 3089 612 3270 617
rect 465 607 470 612
rect 449 602 470 607
rect 553 607 558 612
rect 1857 607 1862 612
rect 2097 607 2102 612
rect 553 602 654 607
rect 737 602 766 607
rect 873 602 1278 607
rect 1369 602 1414 607
rect 1433 602 1862 607
rect 1897 602 1998 607
rect 2025 602 2102 607
rect 2201 602 3158 607
rect 449 597 454 602
rect 761 597 878 602
rect 233 592 454 597
rect 473 592 638 597
rect 953 592 1038 597
rect 1097 592 1238 597
rect 1297 592 1766 597
rect 1817 592 2214 597
rect 2257 592 2638 597
rect 2753 592 2934 597
rect 3017 592 3246 597
rect 3361 592 3398 597
rect 105 582 150 587
rect 353 582 382 587
rect 497 582 582 587
rect 649 582 726 587
rect 825 582 998 587
rect 1065 582 1142 587
rect 1249 582 1302 587
rect 1313 582 1334 587
rect 1345 582 1398 587
rect 1505 582 1558 587
rect 1633 582 1702 587
rect 377 577 502 582
rect 577 577 654 582
rect 1161 577 1254 582
rect 521 572 558 577
rect 553 567 558 572
rect 729 572 838 577
rect 945 572 1166 577
rect 1265 572 1422 577
rect 1457 572 1646 577
rect 729 567 734 572
rect 1761 567 1766 592
rect 1849 582 1958 587
rect 1969 582 2070 587
rect 2129 582 2390 587
rect 2401 582 2462 587
rect 2529 582 2630 587
rect 2665 582 2734 587
rect 3057 582 3126 587
rect 3209 582 3302 587
rect 2753 577 2862 582
rect 3409 577 3414 597
rect 1849 572 2006 577
rect 2049 572 2094 577
rect 2153 572 2238 577
rect 2249 572 2366 577
rect 2449 572 2486 577
rect 2569 572 2758 577
rect 2857 572 2886 577
rect 3025 572 3414 577
rect 2449 567 2454 572
rect 361 562 502 567
rect 553 562 734 567
rect 753 562 814 567
rect 849 562 878 567
rect 361 557 366 562
rect 113 552 222 557
rect 337 552 366 557
rect 497 557 502 562
rect 873 557 878 562
rect 937 562 1054 567
rect 1153 562 1206 567
rect 1249 562 1446 567
rect 1553 562 1654 567
rect 1761 562 1926 567
rect 1953 562 2454 567
rect 2473 562 2926 567
rect 3009 562 3350 567
rect 937 557 942 562
rect 497 552 534 557
rect 873 552 942 557
rect 1009 552 1062 557
rect 1081 552 1238 557
rect 1249 552 1430 557
rect 1489 552 1622 557
rect 1633 552 1926 557
rect 2009 552 2062 557
rect 2145 552 2342 557
rect 2353 552 2414 557
rect 2473 552 2686 557
rect 2745 552 2958 557
rect 3281 552 3390 557
rect 1633 547 1638 552
rect 3281 547 3286 552
rect 273 542 614 547
rect 689 542 822 547
rect 1001 542 1470 547
rect 1553 542 1638 547
rect 1809 542 2518 547
rect 2577 542 2854 547
rect 2865 542 2958 547
rect 3145 542 3286 547
rect 3305 542 3334 547
rect 1553 537 1558 542
rect 2513 537 2518 542
rect 2849 537 2854 542
rect 3329 537 3334 542
rect 3401 542 3446 547
rect 3401 537 3406 542
rect 305 532 422 537
rect 417 527 422 532
rect 529 532 574 537
rect 961 532 1046 537
rect 1089 532 1118 537
rect 1233 532 1558 537
rect 1577 532 1726 537
rect 1889 532 2078 537
rect 2121 532 2222 537
rect 2297 532 2494 537
rect 2513 532 2574 537
rect 2633 532 2734 537
rect 2761 532 2822 537
rect 2849 532 2878 537
rect 3329 532 3406 537
rect 529 527 534 532
rect 1113 527 1238 532
rect 2817 527 2822 532
rect 97 522 318 527
rect 417 522 534 527
rect 553 522 638 527
rect 985 522 1086 527
rect 1257 522 1438 527
rect 1521 522 1926 527
rect 2057 522 2150 527
rect 2233 522 2390 527
rect 2441 522 2478 527
rect 2585 522 2614 527
rect 2817 522 2886 527
rect 3097 522 3174 527
rect 1945 517 2038 522
rect 2145 517 2238 522
rect 1129 512 1254 517
rect 1297 512 1430 517
rect 1441 512 1694 517
rect 1809 512 1830 517
rect 1913 512 1950 517
rect 2033 512 2126 517
rect 2297 512 2598 517
rect 2713 512 2798 517
rect 2905 512 3022 517
rect 3249 512 3422 517
rect 489 502 542 507
rect 537 497 542 502
rect 649 502 1078 507
rect 1097 502 1262 507
rect 1321 502 1478 507
rect 1657 502 1878 507
rect 1889 502 1934 507
rect 1953 502 2038 507
rect 2113 502 2174 507
rect 2257 502 2646 507
rect 3217 502 3278 507
rect 649 497 654 502
rect 1497 497 1638 502
rect 1873 497 1878 502
rect 537 492 654 497
rect 1049 492 1502 497
rect 1633 492 1862 497
rect 1873 492 2030 497
rect 2049 492 2078 497
rect 2185 492 2278 497
rect 2353 492 2454 497
rect 2073 487 2190 492
rect 2473 487 2574 492
rect 1017 482 1310 487
rect 1409 482 1942 487
rect 2225 482 2334 487
rect 2409 482 2478 487
rect 2569 482 2598 487
rect 1025 472 1054 477
rect 1049 467 1054 472
rect 1145 472 1270 477
rect 1289 472 1582 477
rect 1713 472 1790 477
rect 1817 472 1934 477
rect 1953 472 2046 477
rect 2065 472 2206 477
rect 2265 472 2606 477
rect 1145 467 1150 472
rect 265 462 422 467
rect 1049 462 1150 467
rect 1177 462 1206 467
rect 265 447 270 462
rect 417 447 422 462
rect 465 452 558 457
rect 873 452 1030 457
rect 1169 452 1254 457
rect 465 447 470 452
rect 241 442 270 447
rect 289 442 390 447
rect 417 442 470 447
rect 577 442 646 447
rect 289 437 294 442
rect 209 432 294 437
rect 385 437 390 442
rect 577 437 582 442
rect 385 432 406 437
rect 537 432 582 437
rect 641 437 646 442
rect 1249 437 1254 452
rect 1265 447 1270 472
rect 1601 467 1694 472
rect 2065 467 2070 472
rect 1281 462 1606 467
rect 1689 462 1950 467
rect 1969 462 2070 467
rect 2201 467 2206 472
rect 2201 462 2310 467
rect 2369 462 2510 467
rect 2913 462 3006 467
rect 1281 452 1326 457
rect 1449 452 1678 457
rect 1697 447 1862 452
rect 1969 447 1974 462
rect 2089 457 2182 462
rect 2913 457 2918 462
rect 2041 452 2094 457
rect 2177 452 2270 457
rect 2281 452 2366 457
rect 2801 452 2918 457
rect 3001 457 3006 462
rect 3001 452 3030 457
rect 3049 452 3270 457
rect 2385 447 2462 452
rect 1265 442 1366 447
rect 1385 442 1470 447
rect 1481 442 1702 447
rect 1857 442 1886 447
rect 1905 442 1974 447
rect 1993 442 2390 447
rect 2457 442 2534 447
rect 2929 442 2966 447
rect 1361 437 1366 442
rect 1905 437 1910 442
rect 2961 437 2966 442
rect 3049 437 3054 452
rect 641 432 718 437
rect 1185 432 1238 437
rect 1249 432 1286 437
rect 1361 432 1910 437
rect 1929 432 2022 437
rect 2041 432 2166 437
rect 2241 432 2382 437
rect 2393 432 2446 437
rect 2513 432 2622 437
rect 2641 432 2782 437
rect 2961 432 2990 437
rect 3009 432 3054 437
rect 3265 437 3270 452
rect 3265 432 3318 437
rect 305 422 382 427
rect 297 412 374 417
rect 401 412 406 432
rect 2017 427 2022 432
rect 2393 427 2398 432
rect 2641 427 2646 432
rect 457 422 526 427
rect 673 422 702 427
rect 1177 422 1414 427
rect 1425 422 1510 427
rect 1529 422 1566 427
rect 1681 422 1726 427
rect 1737 422 1798 427
rect 1921 422 1942 427
rect 2017 422 2070 427
rect 2145 422 2286 427
rect 2321 422 2398 427
rect 2409 422 2502 427
rect 2569 422 2646 427
rect 2777 427 2782 432
rect 2777 422 2814 427
rect 2833 422 3102 427
rect 3177 422 3254 427
rect 521 417 590 422
rect 673 417 678 422
rect 2497 417 2574 422
rect 2665 417 2758 422
rect 2833 417 2838 422
rect 585 412 678 417
rect 1185 412 1230 417
rect 1345 412 1502 417
rect 1521 412 1622 417
rect 1649 412 2022 417
rect 2137 412 2278 417
rect 2289 412 2406 417
rect 2593 412 2670 417
rect 2753 412 2838 417
rect 2849 412 2926 417
rect 2993 412 3086 417
rect 3153 412 3174 417
rect 249 402 406 407
rect 497 402 566 407
rect 737 402 822 407
rect 1033 402 1126 407
rect 1145 402 1198 407
rect 1305 402 1646 407
rect 1745 402 1822 407
rect 1033 397 1038 402
rect 209 392 326 397
rect 505 392 606 397
rect 729 392 766 397
rect 929 392 1038 397
rect 1121 397 1126 402
rect 1641 397 1750 402
rect 1817 397 1822 402
rect 1929 402 2398 407
rect 2561 402 3062 407
rect 1929 397 1934 402
rect 3057 397 3062 402
rect 3161 402 3190 407
rect 3209 402 3262 407
rect 3161 397 3166 402
rect 3393 397 3398 437
rect 1121 392 1366 397
rect 1457 392 1622 397
rect 1769 392 1798 397
rect 1817 392 1934 397
rect 1953 392 2934 397
rect 2945 392 3038 397
rect 3057 392 3166 397
rect 3353 392 3414 397
rect 313 382 406 387
rect 1049 382 1574 387
rect 1593 382 1678 387
rect 1753 382 1790 387
rect 2009 382 2438 387
rect 2585 382 2790 387
rect 2929 382 2958 387
rect 3321 382 3366 387
rect 697 377 790 382
rect 1569 377 1574 382
rect 1881 377 1990 382
rect 2457 377 2566 382
rect 2785 377 2934 382
rect 113 372 262 377
rect 433 372 654 377
rect 673 372 702 377
rect 785 372 934 377
rect 1321 372 1558 377
rect 1569 372 1886 377
rect 1985 372 2462 377
rect 2561 372 2598 377
rect 2641 372 2766 377
rect 433 367 438 372
rect 409 362 438 367
rect 649 367 654 372
rect 1097 367 1302 372
rect 649 362 1102 367
rect 1297 362 1606 367
rect 1713 362 1830 367
rect 1897 362 2054 367
rect 2073 362 2262 367
rect 457 357 558 362
rect 2049 357 2054 362
rect 2369 357 2374 372
rect 2593 367 2598 372
rect 2393 362 2574 367
rect 2593 362 2622 367
rect 2705 362 2734 367
rect 2857 362 2942 367
rect 2617 357 2710 362
rect 2857 357 2862 362
rect 417 352 462 357
rect 553 352 830 357
rect 1113 352 1534 357
rect 1577 352 1766 357
rect 1777 352 1878 357
rect 1945 352 2014 357
rect 2049 352 2206 357
rect 2217 352 2358 357
rect 2369 352 2430 357
rect 2833 352 2862 357
rect 2937 357 2942 362
rect 3073 362 3158 367
rect 3073 357 3078 362
rect 2937 352 3078 357
rect 3153 357 3158 362
rect 3265 362 3366 367
rect 3265 357 3270 362
rect 3153 352 3270 357
rect 3361 357 3366 362
rect 3361 352 3454 357
rect 825 347 910 352
rect 1113 347 1118 352
rect 1777 347 1782 352
rect 345 342 422 347
rect 433 342 542 347
rect 657 342 678 347
rect 721 342 806 347
rect 905 342 1118 347
rect 1137 342 1206 347
rect 1329 342 1358 347
rect 1465 342 1694 347
rect 1713 342 1782 347
rect 1801 342 2070 347
rect 2169 342 2270 347
rect 2289 342 2414 347
rect 2441 342 2518 347
rect 2689 342 2782 347
rect 2865 342 2926 347
rect 3089 342 3142 347
rect 3281 342 3350 347
rect 657 337 662 342
rect 1353 337 1470 342
rect 1713 337 1718 342
rect 2289 337 2294 342
rect 465 332 662 337
rect 681 332 734 337
rect 865 332 886 337
rect 1489 332 1718 337
rect 1737 332 2294 337
rect 2305 332 2558 337
rect 1249 327 1334 332
rect 225 322 326 327
rect 569 322 694 327
rect 753 322 846 327
rect 225 317 230 322
rect 201 312 230 317
rect 321 317 326 322
rect 753 317 758 322
rect 321 312 350 317
rect 377 312 414 317
rect 553 312 758 317
rect 841 317 846 322
rect 905 322 974 327
rect 1145 322 1254 327
rect 1329 322 1670 327
rect 1689 322 1894 327
rect 2017 322 2214 327
rect 2233 322 2422 327
rect 2505 322 3038 327
rect 3217 322 3342 327
rect 3361 322 3430 327
rect 905 317 910 322
rect 841 312 910 317
rect 969 317 974 322
rect 1889 317 2022 322
rect 2209 317 2214 322
rect 2417 317 2510 322
rect 969 312 1014 317
rect 1105 312 1318 317
rect 217 302 278 307
rect 273 297 278 302
rect 401 302 430 307
rect 561 302 678 307
rect 769 302 878 307
rect 401 297 406 302
rect 273 292 406 297
rect 673 287 678 302
rect 1009 297 1014 312
rect 1313 307 1318 312
rect 1481 312 1870 317
rect 2209 312 2326 317
rect 2529 312 2622 317
rect 2897 312 2926 317
rect 3049 312 3206 317
rect 3305 312 3334 317
rect 1481 307 1486 312
rect 2041 307 2190 312
rect 2321 307 2326 312
rect 2921 307 3054 312
rect 3201 307 3310 312
rect 1033 302 1270 307
rect 1313 302 1486 307
rect 1505 302 1734 307
rect 1849 302 1894 307
rect 2017 302 2046 307
rect 2185 302 2310 307
rect 2321 302 2358 307
rect 2433 302 2750 307
rect 689 292 982 297
rect 1009 292 1158 297
rect 1241 292 1294 297
rect 1625 292 2566 297
rect 1153 287 1246 292
rect 2561 287 2566 292
rect 2705 292 2982 297
rect 3225 292 3310 297
rect 2705 287 2710 292
rect 673 282 902 287
rect 1265 282 1374 287
rect 1401 282 1606 287
rect 1777 282 2158 287
rect 2337 282 2542 287
rect 2561 282 2710 287
rect 1025 277 1134 282
rect 1401 277 1406 282
rect 1601 277 1758 282
rect 2153 277 2342 282
rect 521 272 686 277
rect 753 272 990 277
rect 1001 272 1030 277
rect 1129 272 1366 277
rect 1377 272 1406 277
rect 1753 272 1902 277
rect 2009 272 2134 277
rect 2361 272 2430 277
rect 2729 272 3054 277
rect 1361 267 1366 272
rect 2729 267 2734 272
rect 1041 262 1118 267
rect 1233 262 1318 267
rect 1361 262 2246 267
rect 2273 262 2582 267
rect 2705 262 2734 267
rect 3049 267 3054 272
rect 3049 262 3078 267
rect 1113 257 1238 262
rect 2241 257 2246 262
rect 2841 257 2990 262
rect 969 252 1030 257
rect 1257 252 1310 257
rect 1401 252 1718 257
rect 1817 252 2230 257
rect 2241 252 2846 257
rect 2985 252 3014 257
rect 3049 252 3166 257
rect 1025 247 1094 252
rect 1257 247 1262 252
rect 1305 247 1406 252
rect 1713 247 1822 252
rect 401 242 470 247
rect 713 242 878 247
rect 1089 242 1262 247
rect 1425 242 1454 247
rect 1617 242 1694 247
rect 1449 237 1622 242
rect 1689 237 1694 242
rect 1841 242 2022 247
rect 2049 242 2150 247
rect 2161 242 2198 247
rect 2297 242 2382 247
rect 2433 242 2902 247
rect 2937 242 3102 247
rect 1841 237 1846 242
rect 2193 237 2302 242
rect 2433 237 2438 242
rect 369 232 406 237
rect 665 232 766 237
rect 977 232 1070 237
rect 1289 232 1374 237
rect 1641 232 1670 237
rect 1689 232 1846 237
rect 1865 232 2174 237
rect 2321 232 2438 237
rect 2449 232 2478 237
rect 2585 232 3198 237
rect 977 227 982 232
rect 305 222 422 227
rect 569 222 726 227
rect 897 222 982 227
rect 1001 222 1246 227
rect 1377 222 1558 227
rect 913 217 918 222
rect 1665 217 1670 232
rect 1865 217 1870 232
rect 2473 227 2590 232
rect 1889 222 2254 227
rect 2609 222 2686 227
rect 2833 222 2862 227
rect 2897 222 2998 227
rect 3017 222 3318 227
rect 2833 217 2838 222
rect 393 212 566 217
rect 561 207 566 212
rect 633 212 662 217
rect 697 212 766 217
rect 873 212 918 217
rect 1537 212 1614 217
rect 1665 212 1870 217
rect 1953 212 2838 217
rect 2849 212 2950 217
rect 3025 212 3142 217
rect 633 207 638 212
rect 561 202 638 207
rect 1273 202 1302 207
rect 1385 202 1446 207
rect 1513 202 1550 207
rect 1889 202 1966 207
rect 2041 202 2166 207
rect 3041 202 3094 207
rect 2225 197 2366 202
rect 2881 197 2990 202
rect 449 192 478 197
rect 473 187 478 192
rect 777 192 894 197
rect 1393 192 1462 197
rect 1977 192 2118 197
rect 2201 192 2230 197
rect 2361 192 2502 197
rect 2513 192 2750 197
rect 2857 192 2886 197
rect 2985 192 3046 197
rect 777 187 782 192
rect 2497 187 2502 192
rect 161 182 246 187
rect 161 177 166 182
rect 137 172 166 177
rect 241 177 246 182
rect 289 182 374 187
rect 409 182 438 187
rect 473 182 782 187
rect 1905 182 2038 187
rect 2217 182 2350 187
rect 2497 182 2526 187
rect 2721 182 3094 187
rect 289 177 294 182
rect 241 172 294 177
rect 369 177 374 182
rect 369 172 398 177
rect 1353 172 1894 177
rect 1985 172 2230 177
rect 2697 172 2742 177
rect 3273 172 3350 177
rect 1889 167 1974 172
rect 809 162 982 167
rect 1969 162 2278 167
rect 2297 162 2446 167
rect 2465 162 2758 167
rect 361 157 454 162
rect 809 157 814 162
rect 177 152 366 157
rect 449 152 478 157
rect 585 152 814 157
rect 977 157 982 162
rect 2297 157 2302 162
rect 977 152 1110 157
rect 1241 152 1350 157
rect 1841 152 2046 157
rect 2169 152 2302 157
rect 2441 157 2446 162
rect 2753 157 2758 162
rect 2905 162 3102 167
rect 2905 157 2910 162
rect 2441 152 2510 157
rect 2753 152 2910 157
rect 2929 152 3110 157
rect 2505 147 2510 152
rect 217 142 246 147
rect 241 137 246 142
rect 377 142 422 147
rect 465 142 630 147
rect 377 137 382 142
rect 241 132 382 137
rect 401 132 486 137
rect 481 127 486 132
rect 577 132 606 137
rect 577 127 582 132
rect 481 122 582 127
rect 625 127 630 142
rect 825 142 878 147
rect 825 127 830 142
rect 873 137 878 142
rect 937 142 966 147
rect 1217 142 1262 147
rect 1417 142 1518 147
rect 1721 142 1814 147
rect 1865 142 2486 147
rect 2505 142 2726 147
rect 2929 142 2958 147
rect 937 137 942 142
rect 1721 137 1726 142
rect 873 132 942 137
rect 1633 132 1726 137
rect 1809 127 1814 142
rect 2953 137 2958 142
rect 3041 142 3070 147
rect 3041 137 3046 142
rect 1833 132 1894 137
rect 2953 132 3046 137
rect 3161 132 3310 137
rect 1913 127 2094 132
rect 2201 127 2478 132
rect 625 122 830 127
rect 1257 122 1294 127
rect 1777 122 1798 127
rect 1809 122 1918 127
rect 2089 122 2206 127
rect 2473 122 2646 127
rect 2657 122 2726 127
rect 3161 117 3166 132
rect 3305 117 3310 132
rect 201 112 462 117
rect 1009 112 1230 117
rect 1265 112 1310 117
rect 1385 112 1422 117
rect 1689 112 2078 117
rect 2217 112 2462 117
rect 2617 112 2646 117
rect 2745 112 2774 117
rect 2809 112 2926 117
rect 2945 112 3046 117
rect 3137 112 3166 117
rect 3185 112 3270 117
rect 3305 112 3390 117
rect 2073 107 2222 112
rect 2489 107 2582 112
rect 2641 107 2750 112
rect 2809 107 2814 112
rect 1361 102 1414 107
rect 1721 102 1750 107
rect 1745 97 1750 102
rect 1825 102 1974 107
rect 2009 102 2054 107
rect 2241 102 2398 107
rect 2473 102 2494 107
rect 2577 102 2606 107
rect 2785 102 2814 107
rect 2921 107 2926 112
rect 3185 107 3190 112
rect 2921 102 2982 107
rect 1825 97 1830 102
rect 2393 97 2478 102
rect 2601 97 2606 102
rect 2977 97 2982 102
rect 3057 102 3190 107
rect 3265 107 3270 112
rect 3265 102 3294 107
rect 3057 97 3062 102
rect 441 92 934 97
rect 1377 92 1494 97
rect 1569 92 1710 97
rect 1745 92 1830 97
rect 1945 92 2086 97
rect 2113 92 2230 97
rect 2505 92 2542 97
rect 2601 92 2806 97
rect 2977 92 3062 97
rect 3137 92 3366 97
rect 2225 87 2374 92
rect 2801 87 2806 92
rect 1393 82 1438 87
rect 1857 82 2134 87
rect 2369 82 2446 87
rect 2801 82 2958 87
rect 2953 77 2958 82
rect 3137 77 3142 92
rect 889 72 1366 77
rect 1361 67 1366 72
rect 1505 72 1558 77
rect 1505 67 1510 72
rect 1361 62 1510 67
rect 1553 67 1558 72
rect 1721 72 2358 77
rect 1721 67 1726 72
rect 2353 67 2358 72
rect 2457 72 2782 77
rect 2953 72 3142 77
rect 2457 67 2462 72
rect 1553 62 1726 67
rect 1873 62 1966 67
rect 2001 62 2030 67
rect 2025 57 2030 62
rect 2113 62 2142 67
rect 2353 62 2462 67
rect 2113 57 2118 62
rect 1745 52 1774 57
rect 2025 52 2118 57
rect 2793 52 2934 57
rect 1769 47 1774 52
rect 2793 47 2798 52
rect 1769 42 1862 47
rect 1857 37 1862 42
rect 2153 42 2798 47
rect 2153 37 2158 42
rect 1857 32 2158 37
rect 377 22 1038 27
use AND2X2  AND2X2_0
timestamp 1713453518
transform 1 0 2136 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1713453518
transform 1 0 1552 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1713453518
transform 1 0 3408 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1713453518
transform 1 0 3072 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1713453518
transform 1 0 3128 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1713453518
transform 1 0 3072 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1713453518
transform 1 0 3112 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1713453518
transform 1 0 3296 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1713453518
transform 1 0 3256 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1713453518
transform 1 0 3392 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1713453518
transform 1 0 3336 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1713453518
transform 1 0 1608 0 1 170
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1713453518
transform 1 0 1232 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1713453518
transform 1 0 1120 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1713453518
transform 1 0 1464 0 -1 370
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1713453518
transform 1 0 3328 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1713453518
transform 1 0 1528 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1713453518
transform 1 0 1936 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1713453518
transform 1 0 2128 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1713453518
transform 1 0 1880 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_20
timestamp 1713453518
transform 1 0 3384 0 -1 3170
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1713453518
transform 1 0 2264 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1713453518
transform 1 0 3040 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_23
timestamp 1713453518
transform 1 0 2792 0 -1 2770
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1713453518
transform 1 0 2440 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_25
timestamp 1713453518
transform 1 0 1296 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_26
timestamp 1713453518
transform 1 0 3072 0 -1 2970
box -8 -3 40 105
use AND2X2  AND2X2_27
timestamp 1713453518
transform 1 0 2984 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_28
timestamp 1713453518
transform 1 0 1816 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_29
timestamp 1713453518
transform 1 0 1744 0 1 2370
box -8 -3 40 105
use AND2X2  AND2X2_30
timestamp 1713453518
transform 1 0 3000 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_31
timestamp 1713453518
transform 1 0 1760 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_32
timestamp 1713453518
transform 1 0 2600 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_33
timestamp 1713453518
transform 1 0 1440 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_34
timestamp 1713453518
transform 1 0 2368 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_35
timestamp 1713453518
transform 1 0 584 0 -1 2770
box -8 -3 40 105
use AND2X2  AND2X2_36
timestamp 1713453518
transform 1 0 528 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_37
timestamp 1713453518
transform 1 0 344 0 -1 1170
box -8 -3 40 105
use AND2X2  AND2X2_38
timestamp 1713453518
transform 1 0 432 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_39
timestamp 1713453518
transform 1 0 632 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_40
timestamp 1713453518
transform 1 0 664 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_41
timestamp 1713453518
transform 1 0 408 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_42
timestamp 1713453518
transform 1 0 776 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_43
timestamp 1713453518
transform 1 0 520 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_44
timestamp 1713453518
transform 1 0 712 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_45
timestamp 1713453518
transform 1 0 1056 0 -1 170
box -8 -3 40 105
use AND2X2  AND2X2_46
timestamp 1713453518
transform 1 0 1056 0 1 170
box -8 -3 40 105
use AND2X2  AND2X2_47
timestamp 1713453518
transform 1 0 2392 0 -1 370
box -8 -3 40 105
use AND2X2  AND2X2_48
timestamp 1713453518
transform 1 0 2216 0 -1 370
box -8 -3 40 105
use AND2X2  AND2X2_49
timestamp 1713453518
transform 1 0 3032 0 1 170
box -8 -3 40 105
use AND2X2  AND2X2_50
timestamp 1713453518
transform 1 0 2960 0 -1 370
box -8 -3 40 105
use AND2X2  AND2X2_51
timestamp 1713453518
transform 1 0 2592 0 -1 370
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1713453518
transform 1 0 2512 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1713453518
transform 1 0 2904 0 1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1713453518
transform 1 0 2504 0 1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1713453518
transform 1 0 1920 0 -1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1713453518
transform 1 0 2192 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1713453518
transform 1 0 2976 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1713453518
transform 1 0 3256 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1713453518
transform 1 0 3024 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1713453518
transform 1 0 3352 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1713453518
transform 1 0 2160 0 1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1713453518
transform 1 0 3136 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1713453518
transform 1 0 2840 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1713453518
transform 1 0 2384 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1713453518
transform 1 0 1368 0 -1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1713453518
transform 1 0 2840 0 -1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1713453518
transform 1 0 1360 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1713453518
transform 1 0 3096 0 -1 3170
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1713453518
transform 1 0 3280 0 -1 3370
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1713453518
transform 1 0 3128 0 -1 3370
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1713453518
transform 1 0 3184 0 -1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1713453518
transform 1 0 3184 0 1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1713453518
transform 1 0 1288 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1713453518
transform 1 0 3200 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1713453518
transform 1 0 1240 0 -1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1713453518
transform 1 0 2816 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1713453518
transform 1 0 1504 0 1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1713453518
transform 1 0 2760 0 1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_27
timestamp 1713453518
transform 1 0 1232 0 1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_28
timestamp 1713453518
transform 1 0 2936 0 -1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_29
timestamp 1713453518
transform 1 0 3192 0 1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_30
timestamp 1713453518
transform 1 0 3184 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_31
timestamp 1713453518
transform 1 0 3136 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_32
timestamp 1713453518
transform 1 0 3064 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_33
timestamp 1713453518
transform 1 0 1520 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_34
timestamp 1713453518
transform 1 0 3192 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_35
timestamp 1713453518
transform 1 0 1496 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_36
timestamp 1713453518
transform 1 0 2992 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_37
timestamp 1713453518
transform 1 0 1464 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_38
timestamp 1713453518
transform 1 0 2712 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_39
timestamp 1713453518
transform 1 0 1184 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_40
timestamp 1713453518
transform 1 0 2720 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_41
timestamp 1713453518
transform 1 0 1160 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_42
timestamp 1713453518
transform 1 0 3272 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_43
timestamp 1713453518
transform 1 0 1136 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_44
timestamp 1713453518
transform 1 0 3264 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_45
timestamp 1713453518
transform 1 0 1152 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_46
timestamp 1713453518
transform 1 0 3064 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_47
timestamp 1713453518
transform 1 0 2672 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_48
timestamp 1713453518
transform 1 0 1488 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_49
timestamp 1713453518
transform 1 0 2648 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_50
timestamp 1713453518
transform 1 0 1544 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_51
timestamp 1713453518
transform 1 0 2704 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_52
timestamp 1713453518
transform 1 0 1528 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_53
timestamp 1713453518
transform 1 0 2976 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_54
timestamp 1713453518
transform 1 0 3024 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_55
timestamp 1713453518
transform 1 0 1368 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_56
timestamp 1713453518
transform 1 0 1760 0 -1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_57
timestamp 1713453518
transform 1 0 1400 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_58
timestamp 1713453518
transform 1 0 1880 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_59
timestamp 1713453518
transform 1 0 1288 0 -1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_60
timestamp 1713453518
transform 1 0 1808 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_61
timestamp 1713453518
transform 1 0 1488 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_62
timestamp 1713453518
transform 1 0 1968 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_63
timestamp 1713453518
transform 1 0 408 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_64
timestamp 1713453518
transform 1 0 328 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_65
timestamp 1713453518
transform 1 0 416 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_66
timestamp 1713453518
transform 1 0 560 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_67
timestamp 1713453518
transform 1 0 592 0 1 1770
box -7 -3 39 105
use AOI21X1  AOI21X1_68
timestamp 1713453518
transform 1 0 568 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_69
timestamp 1713453518
transform 1 0 536 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_70
timestamp 1713453518
transform 1 0 440 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_71
timestamp 1713453518
transform 1 0 424 0 -1 370
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1713453518
transform 1 0 2232 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1713453518
transform 1 0 3008 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1713453518
transform 1 0 2312 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1713453518
transform 1 0 2680 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1713453518
transform 1 0 2648 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1713453518
transform 1 0 2688 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1713453518
transform 1 0 2552 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1713453518
transform 1 0 2616 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1713453518
transform 1 0 2952 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1713453518
transform 1 0 2768 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1713453518
transform 1 0 2784 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1713453518
transform 1 0 2208 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1713453518
transform 1 0 2504 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1713453518
transform 1 0 2648 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1713453518
transform 1 0 2512 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1713453518
transform 1 0 2536 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1713453518
transform 1 0 2232 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1713453518
transform 1 0 2272 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1713453518
transform 1 0 2320 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1713453518
transform 1 0 2408 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1713453518
transform 1 0 2240 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1713453518
transform 1 0 2008 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1713453518
transform 1 0 2320 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1713453518
transform 1 0 2328 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1713453518
transform 1 0 2344 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1713453518
transform 1 0 2056 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1713453518
transform 1 0 1712 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1713453518
transform 1 0 2032 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1713453518
transform 1 0 1864 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1713453518
transform 1 0 2104 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1713453518
transform 1 0 1424 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1713453518
transform 1 0 2920 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1713453518
transform 1 0 2296 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1713453518
transform 1 0 2200 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1713453518
transform 1 0 2296 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1713453518
transform 1 0 2136 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1713453518
transform 1 0 2144 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1713453518
transform 1 0 2160 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1713453518
transform 1 0 2176 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1713453518
transform 1 0 1896 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1713453518
transform 1 0 1936 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1713453518
transform 1 0 1856 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1713453518
transform 1 0 3032 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1713453518
transform 1 0 3312 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1713453518
transform 1 0 3144 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1713453518
transform 1 0 2864 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1713453518
transform 1 0 2992 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1713453518
transform 1 0 2848 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1713453518
transform 1 0 3056 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1713453518
transform 1 0 3296 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1713453518
transform 1 0 3336 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1713453518
transform 1 0 3352 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1713453518
transform 1 0 3232 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1713453518
transform 1 0 2896 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1713453518
transform 1 0 3096 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_55
timestamp 1713453518
transform 1 0 2864 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1713453518
transform 1 0 2744 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_57
timestamp 1713453518
transform 1 0 2488 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_58
timestamp 1713453518
transform 1 0 2536 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_59
timestamp 1713453518
transform 1 0 2560 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_60
timestamp 1713453518
transform 1 0 2832 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_61
timestamp 1713453518
transform 1 0 2888 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_62
timestamp 1713453518
transform 1 0 2904 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_63
timestamp 1713453518
transform 1 0 3360 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_64
timestamp 1713453518
transform 1 0 3360 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_65
timestamp 1713453518
transform 1 0 3296 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_66
timestamp 1713453518
transform 1 0 2040 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_67
timestamp 1713453518
transform 1 0 3360 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_68
timestamp 1713453518
transform 1 0 2864 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_69
timestamp 1713453518
transform 1 0 2808 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_70
timestamp 1713453518
transform 1 0 2960 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_71
timestamp 1713453518
transform 1 0 2968 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1713453518
transform 1 0 2528 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_73
timestamp 1713453518
transform 1 0 2600 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_74
timestamp 1713453518
transform 1 0 2560 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_75
timestamp 1713453518
transform 1 0 2848 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_76
timestamp 1713453518
transform 1 0 2832 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_77
timestamp 1713453518
transform 1 0 2624 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_78
timestamp 1713453518
transform 1 0 2496 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_79
timestamp 1713453518
transform 1 0 2392 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_80
timestamp 1713453518
transform 1 0 2408 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_81
timestamp 1713453518
transform 1 0 2392 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_82
timestamp 1713453518
transform 1 0 1608 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_83
timestamp 1713453518
transform 1 0 1504 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_84
timestamp 1713453518
transform 1 0 1712 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_85
timestamp 1713453518
transform 1 0 2232 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_86
timestamp 1713453518
transform 1 0 1904 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_87
timestamp 1713453518
transform 1 0 2808 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_88
timestamp 1713453518
transform 1 0 2616 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_89
timestamp 1713453518
transform 1 0 2080 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_90
timestamp 1713453518
transform 1 0 3232 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_91
timestamp 1713453518
transform 1 0 2728 0 -1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_92
timestamp 1713453518
transform 1 0 2368 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_93
timestamp 1713453518
transform 1 0 3296 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_94
timestamp 1713453518
transform 1 0 2712 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_95
timestamp 1713453518
transform 1 0 2296 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_96
timestamp 1713453518
transform 1 0 3368 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_97
timestamp 1713453518
transform 1 0 2608 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_98
timestamp 1713453518
transform 1 0 2120 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_99
timestamp 1713453518
transform 1 0 3304 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_100
timestamp 1713453518
transform 1 0 1272 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_101
timestamp 1713453518
transform 1 0 2424 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_102
timestamp 1713453518
transform 1 0 1976 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_103
timestamp 1713453518
transform 1 0 3344 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_104
timestamp 1713453518
transform 1 0 2440 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_105
timestamp 1713453518
transform 1 0 1904 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_106
timestamp 1713453518
transform 1 0 3400 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_107
timestamp 1713453518
transform 1 0 2344 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_108
timestamp 1713453518
transform 1 0 1984 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_109
timestamp 1713453518
transform 1 0 2968 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_110
timestamp 1713453518
transform 1 0 2296 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_111
timestamp 1713453518
transform 1 0 2072 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_112
timestamp 1713453518
transform 1 0 2992 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_113
timestamp 1713453518
transform 1 0 1184 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_114
timestamp 1713453518
transform 1 0 2296 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_115
timestamp 1713453518
transform 1 0 2128 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_116
timestamp 1713453518
transform 1 0 3128 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_117
timestamp 1713453518
transform 1 0 2440 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_118
timestamp 1713453518
transform 1 0 1920 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_119
timestamp 1713453518
transform 1 0 3392 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_120
timestamp 1713453518
transform 1 0 2552 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_121
timestamp 1713453518
transform 1 0 2352 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_122
timestamp 1713453518
transform 1 0 3392 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_123
timestamp 1713453518
transform 1 0 2504 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_124
timestamp 1713453518
transform 1 0 2128 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_125
timestamp 1713453518
transform 1 0 3392 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_126
timestamp 1713453518
transform 1 0 1240 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_127
timestamp 1713453518
transform 1 0 2496 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_128
timestamp 1713453518
transform 1 0 2024 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_129
timestamp 1713453518
transform 1 0 3328 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_130
timestamp 1713453518
transform 1 0 2480 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_131
timestamp 1713453518
transform 1 0 2136 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_132
timestamp 1713453518
transform 1 0 3336 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_133
timestamp 1713453518
transform 1 0 2416 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_134
timestamp 1713453518
transform 1 0 2104 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_135
timestamp 1713453518
transform 1 0 3240 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_136
timestamp 1713453518
transform 1 0 2360 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_137
timestamp 1713453518
transform 1 0 1992 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_138
timestamp 1713453518
transform 1 0 2944 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_139
timestamp 1713453518
transform 1 0 1152 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_140
timestamp 1713453518
transform 1 0 2296 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_141
timestamp 1713453518
transform 1 0 1896 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_142
timestamp 1713453518
transform 1 0 2920 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_143
timestamp 1713453518
transform 1 0 2304 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_144
timestamp 1713453518
transform 1 0 1984 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_145
timestamp 1713453518
transform 1 0 3248 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_146
timestamp 1713453518
transform 1 0 2328 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_147
timestamp 1713453518
transform 1 0 2088 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_148
timestamp 1713453518
transform 1 0 3048 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_149
timestamp 1713453518
transform 1 0 2312 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_150
timestamp 1713453518
transform 1 0 1808 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_151
timestamp 1713453518
transform 1 0 2936 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_152
timestamp 1713453518
transform 1 0 1280 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_153
timestamp 1713453518
transform 1 0 1288 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_154
timestamp 1713453518
transform 1 0 2280 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_155
timestamp 1713453518
transform 1 0 2064 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_156
timestamp 1713453518
transform 1 0 2800 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_157
timestamp 1713453518
transform 1 0 2320 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_158
timestamp 1713453518
transform 1 0 2128 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_159
timestamp 1713453518
transform 1 0 2800 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_160
timestamp 1713453518
transform 1 0 2344 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_161
timestamp 1713453518
transform 1 0 2112 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_162
timestamp 1713453518
transform 1 0 2912 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_163
timestamp 1713453518
transform 1 0 2160 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_164
timestamp 1713453518
transform 1 0 2896 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_165
timestamp 1713453518
transform 1 0 1384 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_166
timestamp 1713453518
transform 1 0 1936 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_167
timestamp 1713453518
transform 1 0 1928 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_168
timestamp 1713453518
transform 1 0 1864 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_169
timestamp 1713453518
transform 1 0 1664 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_170
timestamp 1713453518
transform 1 0 1608 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_171
timestamp 1713453518
transform 1 0 3008 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_172
timestamp 1713453518
transform 1 0 2880 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_173
timestamp 1713453518
transform 1 0 2696 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_174
timestamp 1713453518
transform 1 0 2592 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_175
timestamp 1713453518
transform 1 0 3064 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_176
timestamp 1713453518
transform 1 0 2008 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_177
timestamp 1713453518
transform 1 0 304 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_178
timestamp 1713453518
transform 1 0 344 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_179
timestamp 1713453518
transform 1 0 408 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_180
timestamp 1713453518
transform 1 0 584 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_181
timestamp 1713453518
transform 1 0 440 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_182
timestamp 1713453518
transform 1 0 536 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_183
timestamp 1713453518
transform 1 0 400 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_184
timestamp 1713453518
transform 1 0 528 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_185
timestamp 1713453518
transform 1 0 384 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_186
timestamp 1713453518
transform 1 0 624 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_187
timestamp 1713453518
transform 1 0 400 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_188
timestamp 1713453518
transform 1 0 608 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_189
timestamp 1713453518
transform 1 0 368 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_190
timestamp 1713453518
transform 1 0 672 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_191
timestamp 1713453518
transform 1 0 328 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_192
timestamp 1713453518
transform 1 0 648 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_193
timestamp 1713453518
transform 1 0 416 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_194
timestamp 1713453518
transform 1 0 696 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_195
timestamp 1713453518
transform 1 0 440 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_196
timestamp 1713453518
transform 1 0 560 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_197
timestamp 1713453518
transform 1 0 440 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_198
timestamp 1713453518
transform 1 0 648 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_199
timestamp 1713453518
transform 1 0 440 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_200
timestamp 1713453518
transform 1 0 712 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_201
timestamp 1713453518
transform 1 0 480 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_202
timestamp 1713453518
transform 1 0 752 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_203
timestamp 1713453518
transform 1 0 576 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_204
timestamp 1713453518
transform 1 0 608 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_205
timestamp 1713453518
transform 1 0 392 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_206
timestamp 1713453518
transform 1 0 664 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_207
timestamp 1713453518
transform 1 0 424 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_208
timestamp 1713453518
transform 1 0 768 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_209
timestamp 1713453518
transform 1 0 480 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_210
timestamp 1713453518
transform 1 0 752 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_211
timestamp 1713453518
transform 1 0 440 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_212
timestamp 1713453518
transform 1 0 648 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_213
timestamp 1713453518
transform 1 0 640 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_214
timestamp 1713453518
transform 1 0 736 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_215
timestamp 1713453518
transform 1 0 640 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_216
timestamp 1713453518
transform 1 0 736 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_217
timestamp 1713453518
transform 1 0 520 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_218
timestamp 1713453518
transform 1 0 672 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_219
timestamp 1713453518
transform 1 0 400 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_220
timestamp 1713453518
transform 1 0 496 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_221
timestamp 1713453518
transform 1 0 520 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_222
timestamp 1713453518
transform 1 0 672 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_223
timestamp 1713453518
transform 1 0 448 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_224
timestamp 1713453518
transform 1 0 624 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_225
timestamp 1713453518
transform 1 0 456 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_226
timestamp 1713453518
transform 1 0 552 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_227
timestamp 1713453518
transform 1 0 584 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_228
timestamp 1713453518
transform 1 0 384 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_229
timestamp 1713453518
transform 1 0 400 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_230
timestamp 1713453518
transform 1 0 440 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_231
timestamp 1713453518
transform 1 0 384 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_232
timestamp 1713453518
transform 1 0 728 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_233
timestamp 1713453518
transform 1 0 664 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_234
timestamp 1713453518
transform 1 0 752 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_235
timestamp 1713453518
transform 1 0 736 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_236
timestamp 1713453518
transform 1 0 760 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_237
timestamp 1713453518
transform 1 0 696 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_238
timestamp 1713453518
transform 1 0 720 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_239
timestamp 1713453518
transform 1 0 752 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_240
timestamp 1713453518
transform 1 0 768 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_241
timestamp 1713453518
transform 1 0 704 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_242
timestamp 1713453518
transform 1 0 752 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_243
timestamp 1713453518
transform 1 0 832 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_244
timestamp 1713453518
transform 1 0 808 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_245
timestamp 1713453518
transform 1 0 808 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_246
timestamp 1713453518
transform 1 0 904 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_247
timestamp 1713453518
transform 1 0 968 0 1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_248
timestamp 1713453518
transform 1 0 896 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_249
timestamp 1713453518
transform 1 0 920 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_250
timestamp 1713453518
transform 1 0 848 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_251
timestamp 1713453518
transform 1 0 824 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_252
timestamp 1713453518
transform 1 0 792 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_253
timestamp 1713453518
transform 1 0 824 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_254
timestamp 1713453518
transform 1 0 856 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_255
timestamp 1713453518
transform 1 0 824 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_256
timestamp 1713453518
transform 1 0 768 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_257
timestamp 1713453518
transform 1 0 800 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_258
timestamp 1713453518
transform 1 0 784 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_259
timestamp 1713453518
transform 1 0 840 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_260
timestamp 1713453518
transform 1 0 888 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_261
timestamp 1713453518
transform 1 0 864 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_262
timestamp 1713453518
transform 1 0 920 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_263
timestamp 1713453518
transform 1 0 760 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_264
timestamp 1713453518
transform 1 0 848 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_265
timestamp 1713453518
transform 1 0 768 0 -1 970
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1713453518
transform 1 0 696 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1713453518
transform 1 0 712 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1713453518
transform 1 0 1688 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1713453518
transform 1 0 72 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1713453518
transform 1 0 96 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1713453518
transform 1 0 376 0 -1 170
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1713453518
transform 1 0 1584 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1713453518
transform 1 0 1480 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1713453518
transform 1 0 1480 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1713453518
transform 1 0 1544 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1713453518
transform 1 0 1096 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1713453518
transform 1 0 384 0 -1 370
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1713453518
transform 1 0 320 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1713453518
transform 1 0 1056 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1713453518
transform 1 0 1264 0 -1 370
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1713453518
transform 1 0 776 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1713453518
transform 1 0 832 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1713453518
transform 1 0 752 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1713453518
transform 1 0 856 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1713453518
transform 1 0 824 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1713453518
transform 1 0 840 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_21
timestamp 1713453518
transform 1 0 816 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_22
timestamp 1713453518
transform 1 0 3144 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_23
timestamp 1713453518
transform 1 0 720 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1713453518
transform 1 0 728 0 1 1170
box -5 -3 28 105
use BUFX2  BUFX2_25
timestamp 1713453518
transform 1 0 704 0 1 1170
box -5 -3 28 105
use BUFX2  BUFX2_26
timestamp 1713453518
transform 1 0 800 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_27
timestamp 1713453518
transform 1 0 896 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_28
timestamp 1713453518
transform 1 0 808 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_29
timestamp 1713453518
transform 1 0 2392 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_30
timestamp 1713453518
transform 1 0 2192 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_31
timestamp 1713453518
transform 1 0 608 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_32
timestamp 1713453518
transform 1 0 472 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_33
timestamp 1713453518
transform 1 0 2536 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_34
timestamp 1713453518
transform 1 0 2176 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_35
timestamp 1713453518
transform 1 0 2568 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_36
timestamp 1713453518
transform 1 0 2152 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_37
timestamp 1713453518
transform 1 0 2216 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_38
timestamp 1713453518
transform 1 0 3104 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_39
timestamp 1713453518
transform 1 0 1344 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_40
timestamp 1713453518
transform 1 0 1040 0 1 770
box -5 -3 28 105
use BUFX2  BUFX2_41
timestamp 1713453518
transform 1 0 1032 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_42
timestamp 1713453518
transform 1 0 2216 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_43
timestamp 1713453518
transform 1 0 2976 0 1 570
box -5 -3 28 105
use BUFX2  BUFX2_44
timestamp 1713453518
transform 1 0 1872 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_45
timestamp 1713453518
transform 1 0 1840 0 -1 2170
box -5 -3 28 105
use BUFX2  BUFX2_46
timestamp 1713453518
transform 1 0 464 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_47
timestamp 1713453518
transform 1 0 480 0 -1 2170
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1713453518
transform 1 0 2344 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1713453518
transform 1 0 2232 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1713453518
transform 1 0 1680 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1713453518
transform 1 0 1792 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1713453518
transform 1 0 3152 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1713453518
transform 1 0 3280 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1713453518
transform 1 0 3256 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1713453518
transform 1 0 3040 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1713453518
transform 1 0 3352 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1713453518
transform 1 0 1704 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1713453518
transform 1 0 1568 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1713453518
transform 1 0 1576 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1713453518
transform 1 0 1320 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1713453518
transform 1 0 1048 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1713453518
transform 1 0 2480 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1713453518
transform 1 0 2112 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1713453518
transform 1 0 3000 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1713453518
transform 1 0 2920 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1713453518
transform 1 0 2632 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1713453518
transform 1 0 2672 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1713453518
transform 1 0 2808 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1713453518
transform 1 0 792 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1713453518
transform 1 0 736 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1713453518
transform 1 0 784 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1713453518
transform 1 0 880 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1713453518
transform 1 0 912 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1713453518
transform 1 0 1008 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1713453518
transform 1 0 984 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1713453518
transform 1 0 936 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1713453518
transform 1 0 944 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1713453518
transform 1 0 904 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1713453518
transform 1 0 888 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1713453518
transform 1 0 936 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1713453518
transform 1 0 912 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1713453518
transform 1 0 856 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1713453518
transform 1 0 880 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1713453518
transform 1 0 896 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1713453518
transform 1 0 904 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1713453518
transform 1 0 944 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1713453518
transform 1 0 944 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1713453518
transform 1 0 896 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1713453518
transform 1 0 856 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1713453518
transform 1 0 936 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1713453518
transform 1 0 816 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1713453518
transform 1 0 912 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1713453518
transform 1 0 840 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1713453518
transform 1 0 888 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1713453518
transform 1 0 896 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1713453518
transform 1 0 840 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1713453518
transform 1 0 904 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1713453518
transform 1 0 936 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1713453518
transform 1 0 896 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1713453518
transform 1 0 736 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1713453518
transform 1 0 792 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1713453518
transform 1 0 480 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1713453518
transform 1 0 80 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1713453518
transform 1 0 80 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1713453518
transform 1 0 72 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1713453518
transform 1 0 168 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1713453518
transform 1 0 296 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1713453518
transform 1 0 504 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1713453518
transform 1 0 512 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1713453518
transform 1 0 80 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1713453518
transform 1 0 104 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1713453518
transform 1 0 88 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1713453518
transform 1 0 80 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1713453518
transform 1 0 80 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1713453518
transform 1 0 256 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1713453518
transform 1 0 80 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1713453518
transform 1 0 88 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1713453518
transform 1 0 88 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1713453518
transform 1 0 80 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1713453518
transform 1 0 88 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1713453518
transform 1 0 192 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1713453518
transform 1 0 208 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1713453518
transform 1 0 80 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1713453518
transform 1 0 80 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1713453518
transform 1 0 88 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1713453518
transform 1 0 80 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1713453518
transform 1 0 200 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1713453518
transform 1 0 96 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1713453518
transform 1 0 88 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1713453518
transform 1 0 80 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1713453518
transform 1 0 304 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1713453518
transform 1 0 152 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1713453518
transform 1 0 624 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1713453518
transform 1 0 304 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1713453518
transform 1 0 680 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1713453518
transform 1 0 280 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1713453518
transform 1 0 296 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1713453518
transform 1 0 272 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1713453518
transform 1 0 384 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1713453518
transform 1 0 368 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1713453518
transform 1 0 688 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1713453518
transform 1 0 688 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1713453518
transform 1 0 312 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1713453518
transform 1 0 360 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1713453518
transform 1 0 368 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1713453518
transform 1 0 312 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1713453518
transform 1 0 248 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1713453518
transform 1 0 472 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1713453518
transform 1 0 312 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1713453518
transform 1 0 312 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1713453518
transform 1 0 320 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1713453518
transform 1 0 304 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1713453518
transform 1 0 776 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1713453518
transform 1 0 720 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1713453518
transform 1 0 776 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1713453518
transform 1 0 256 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1713453518
transform 1 0 280 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1713453518
transform 1 0 320 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1713453518
transform 1 0 296 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1713453518
transform 1 0 200 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1713453518
transform 1 0 160 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1713453518
transform 1 0 264 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1713453518
transform 1 0 88 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1713453518
transform 1 0 600 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1713453518
transform 1 0 408 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1713453518
transform 1 0 776 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1713453518
transform 1 0 400 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1713453518
transform 1 0 1104 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1713453518
transform 1 0 944 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1713453518
transform 1 0 952 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1713453518
transform 1 0 1096 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1713453518
transform 1 0 624 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1713453518
transform 1 0 512 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1713453518
transform 1 0 576 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1713453518
transform 1 0 840 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_128
timestamp 1713453518
transform 1 0 736 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1713453518
transform 1 0 456 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_130
timestamp 1713453518
transform 1 0 256 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_131
timestamp 1713453518
transform 1 0 88 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_132
timestamp 1713453518
transform 1 0 128 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_133
timestamp 1713453518
transform 1 0 208 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1713453518
transform 1 0 80 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_135
timestamp 1713453518
transform 1 0 248 0 1 170
box -8 -3 104 105
use FILL  FILL_0
timestamp 1713453518
transform 1 0 3440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_1
timestamp 1713453518
transform 1 0 3432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2
timestamp 1713453518
transform 1 0 3424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3
timestamp 1713453518
transform 1 0 3416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_4
timestamp 1713453518
transform 1 0 3408 0 -1 3370
box -8 -3 16 105
use FILL  FILL_5
timestamp 1713453518
transform 1 0 3400 0 -1 3370
box -8 -3 16 105
use FILL  FILL_6
timestamp 1713453518
transform 1 0 3392 0 -1 3370
box -8 -3 16 105
use FILL  FILL_7
timestamp 1713453518
transform 1 0 3312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_8
timestamp 1713453518
transform 1 0 3272 0 -1 3370
box -8 -3 16 105
use FILL  FILL_9
timestamp 1713453518
transform 1 0 3264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_10
timestamp 1713453518
transform 1 0 3256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_11
timestamp 1713453518
transform 1 0 3168 0 -1 3370
box -8 -3 16 105
use FILL  FILL_12
timestamp 1713453518
transform 1 0 3160 0 -1 3370
box -8 -3 16 105
use FILL  FILL_13
timestamp 1713453518
transform 1 0 3088 0 -1 3370
box -8 -3 16 105
use FILL  FILL_14
timestamp 1713453518
transform 1 0 3080 0 -1 3370
box -8 -3 16 105
use FILL  FILL_15
timestamp 1713453518
transform 1 0 3024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_16
timestamp 1713453518
transform 1 0 3016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_17
timestamp 1713453518
transform 1 0 3008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_18
timestamp 1713453518
transform 1 0 2984 0 -1 3370
box -8 -3 16 105
use FILL  FILL_19
timestamp 1713453518
transform 1 0 2944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_20
timestamp 1713453518
transform 1 0 2936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_21
timestamp 1713453518
transform 1 0 2896 0 -1 3370
box -8 -3 16 105
use FILL  FILL_22
timestamp 1713453518
transform 1 0 2888 0 -1 3370
box -8 -3 16 105
use FILL  FILL_23
timestamp 1713453518
transform 1 0 2840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_24
timestamp 1713453518
transform 1 0 2832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_25
timestamp 1713453518
transform 1 0 2824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_26
timestamp 1713453518
transform 1 0 2792 0 -1 3370
box -8 -3 16 105
use FILL  FILL_27
timestamp 1713453518
transform 1 0 2784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_28
timestamp 1713453518
transform 1 0 2776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_29
timestamp 1713453518
transform 1 0 2768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_30
timestamp 1713453518
transform 1 0 2720 0 -1 3370
box -8 -3 16 105
use FILL  FILL_31
timestamp 1713453518
transform 1 0 2712 0 -1 3370
box -8 -3 16 105
use FILL  FILL_32
timestamp 1713453518
transform 1 0 2704 0 -1 3370
box -8 -3 16 105
use FILL  FILL_33
timestamp 1713453518
transform 1 0 2696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_34
timestamp 1713453518
transform 1 0 2688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_35
timestamp 1713453518
transform 1 0 2640 0 -1 3370
box -8 -3 16 105
use FILL  FILL_36
timestamp 1713453518
transform 1 0 2632 0 -1 3370
box -8 -3 16 105
use FILL  FILL_37
timestamp 1713453518
transform 1 0 2624 0 -1 3370
box -8 -3 16 105
use FILL  FILL_38
timestamp 1713453518
transform 1 0 2616 0 -1 3370
box -8 -3 16 105
use FILL  FILL_39
timestamp 1713453518
transform 1 0 2608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_40
timestamp 1713453518
transform 1 0 2576 0 -1 3370
box -8 -3 16 105
use FILL  FILL_41
timestamp 1713453518
transform 1 0 2568 0 -1 3370
box -8 -3 16 105
use FILL  FILL_42
timestamp 1713453518
transform 1 0 2528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_43
timestamp 1713453518
transform 1 0 2520 0 -1 3370
box -8 -3 16 105
use FILL  FILL_44
timestamp 1713453518
transform 1 0 2512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_45
timestamp 1713453518
transform 1 0 2504 0 -1 3370
box -8 -3 16 105
use FILL  FILL_46
timestamp 1713453518
transform 1 0 2496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_47
timestamp 1713453518
transform 1 0 2488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_48
timestamp 1713453518
transform 1 0 2456 0 -1 3370
box -8 -3 16 105
use FILL  FILL_49
timestamp 1713453518
transform 1 0 2448 0 -1 3370
box -8 -3 16 105
use FILL  FILL_50
timestamp 1713453518
transform 1 0 2440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_51
timestamp 1713453518
transform 1 0 2408 0 -1 3370
box -8 -3 16 105
use FILL  FILL_52
timestamp 1713453518
transform 1 0 2400 0 -1 3370
box -8 -3 16 105
use FILL  FILL_53
timestamp 1713453518
transform 1 0 2392 0 -1 3370
box -8 -3 16 105
use FILL  FILL_54
timestamp 1713453518
transform 1 0 2384 0 -1 3370
box -8 -3 16 105
use FILL  FILL_55
timestamp 1713453518
transform 1 0 2376 0 -1 3370
box -8 -3 16 105
use FILL  FILL_56
timestamp 1713453518
transform 1 0 2368 0 -1 3370
box -8 -3 16 105
use FILL  FILL_57
timestamp 1713453518
transform 1 0 2320 0 -1 3370
box -8 -3 16 105
use FILL  FILL_58
timestamp 1713453518
transform 1 0 2312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_59
timestamp 1713453518
transform 1 0 2304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_60
timestamp 1713453518
transform 1 0 2296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_61
timestamp 1713453518
transform 1 0 2288 0 -1 3370
box -8 -3 16 105
use FILL  FILL_62
timestamp 1713453518
transform 1 0 2280 0 -1 3370
box -8 -3 16 105
use FILL  FILL_63
timestamp 1713453518
transform 1 0 2248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_64
timestamp 1713453518
transform 1 0 2240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_65
timestamp 1713453518
transform 1 0 2232 0 -1 3370
box -8 -3 16 105
use FILL  FILL_66
timestamp 1713453518
transform 1 0 2224 0 -1 3370
box -8 -3 16 105
use FILL  FILL_67
timestamp 1713453518
transform 1 0 2192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_68
timestamp 1713453518
transform 1 0 2184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_69
timestamp 1713453518
transform 1 0 2176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_70
timestamp 1713453518
transform 1 0 2168 0 -1 3370
box -8 -3 16 105
use FILL  FILL_71
timestamp 1713453518
transform 1 0 2144 0 -1 3370
box -8 -3 16 105
use FILL  FILL_72
timestamp 1713453518
transform 1 0 2136 0 -1 3370
box -8 -3 16 105
use FILL  FILL_73
timestamp 1713453518
transform 1 0 2128 0 -1 3370
box -8 -3 16 105
use FILL  FILL_74
timestamp 1713453518
transform 1 0 2120 0 -1 3370
box -8 -3 16 105
use FILL  FILL_75
timestamp 1713453518
transform 1 0 2072 0 -1 3370
box -8 -3 16 105
use FILL  FILL_76
timestamp 1713453518
transform 1 0 2064 0 -1 3370
box -8 -3 16 105
use FILL  FILL_77
timestamp 1713453518
transform 1 0 2056 0 -1 3370
box -8 -3 16 105
use FILL  FILL_78
timestamp 1713453518
transform 1 0 2048 0 -1 3370
box -8 -3 16 105
use FILL  FILL_79
timestamp 1713453518
transform 1 0 2040 0 -1 3370
box -8 -3 16 105
use FILL  FILL_80
timestamp 1713453518
transform 1 0 2032 0 -1 3370
box -8 -3 16 105
use FILL  FILL_81
timestamp 1713453518
transform 1 0 2024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_82
timestamp 1713453518
transform 1 0 2016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_83
timestamp 1713453518
transform 1 0 1976 0 -1 3370
box -8 -3 16 105
use FILL  FILL_84
timestamp 1713453518
transform 1 0 1968 0 -1 3370
box -8 -3 16 105
use FILL  FILL_85
timestamp 1713453518
transform 1 0 1960 0 -1 3370
box -8 -3 16 105
use FILL  FILL_86
timestamp 1713453518
transform 1 0 1920 0 -1 3370
box -8 -3 16 105
use FILL  FILL_87
timestamp 1713453518
transform 1 0 1912 0 -1 3370
box -8 -3 16 105
use FILL  FILL_88
timestamp 1713453518
transform 1 0 1904 0 -1 3370
box -8 -3 16 105
use FILL  FILL_89
timestamp 1713453518
transform 1 0 1896 0 -1 3370
box -8 -3 16 105
use FILL  FILL_90
timestamp 1713453518
transform 1 0 1864 0 -1 3370
box -8 -3 16 105
use FILL  FILL_91
timestamp 1713453518
transform 1 0 1856 0 -1 3370
box -8 -3 16 105
use FILL  FILL_92
timestamp 1713453518
transform 1 0 1848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_93
timestamp 1713453518
transform 1 0 1840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_94
timestamp 1713453518
transform 1 0 1832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_95
timestamp 1713453518
transform 1 0 1792 0 -1 3370
box -8 -3 16 105
use FILL  FILL_96
timestamp 1713453518
transform 1 0 1784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_97
timestamp 1713453518
transform 1 0 1776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_98
timestamp 1713453518
transform 1 0 1768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_99
timestamp 1713453518
transform 1 0 1760 0 -1 3370
box -8 -3 16 105
use FILL  FILL_100
timestamp 1713453518
transform 1 0 1752 0 -1 3370
box -8 -3 16 105
use FILL  FILL_101
timestamp 1713453518
transform 1 0 1744 0 -1 3370
box -8 -3 16 105
use FILL  FILL_102
timestamp 1713453518
transform 1 0 1696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_103
timestamp 1713453518
transform 1 0 1688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_104
timestamp 1713453518
transform 1 0 1680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_105
timestamp 1713453518
transform 1 0 1672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_106
timestamp 1713453518
transform 1 0 1664 0 -1 3370
box -8 -3 16 105
use FILL  FILL_107
timestamp 1713453518
transform 1 0 1656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_108
timestamp 1713453518
transform 1 0 1648 0 -1 3370
box -8 -3 16 105
use FILL  FILL_109
timestamp 1713453518
transform 1 0 1600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_110
timestamp 1713453518
transform 1 0 1592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_111
timestamp 1713453518
transform 1 0 1584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_112
timestamp 1713453518
transform 1 0 1576 0 -1 3370
box -8 -3 16 105
use FILL  FILL_113
timestamp 1713453518
transform 1 0 1536 0 -1 3370
box -8 -3 16 105
use FILL  FILL_114
timestamp 1713453518
transform 1 0 1528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_115
timestamp 1713453518
transform 1 0 1520 0 -1 3370
box -8 -3 16 105
use FILL  FILL_116
timestamp 1713453518
transform 1 0 1512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_117
timestamp 1713453518
transform 1 0 1440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_118
timestamp 1713453518
transform 1 0 1432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_119
timestamp 1713453518
transform 1 0 1424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_120
timestamp 1713453518
transform 1 0 1416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_121
timestamp 1713453518
transform 1 0 1408 0 -1 3370
box -8 -3 16 105
use FILL  FILL_122
timestamp 1713453518
transform 1 0 1336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_123
timestamp 1713453518
transform 1 0 1328 0 -1 3370
box -8 -3 16 105
use FILL  FILL_124
timestamp 1713453518
transform 1 0 1304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_125
timestamp 1713453518
transform 1 0 1296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_126
timestamp 1713453518
transform 1 0 1232 0 -1 3370
box -8 -3 16 105
use FILL  FILL_127
timestamp 1713453518
transform 1 0 1224 0 -1 3370
box -8 -3 16 105
use FILL  FILL_128
timestamp 1713453518
transform 1 0 1216 0 -1 3370
box -8 -3 16 105
use FILL  FILL_129
timestamp 1713453518
transform 1 0 1208 0 -1 3370
box -8 -3 16 105
use FILL  FILL_130
timestamp 1713453518
transform 1 0 1152 0 -1 3370
box -8 -3 16 105
use FILL  FILL_131
timestamp 1713453518
transform 1 0 1112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_132
timestamp 1713453518
transform 1 0 1104 0 -1 3370
box -8 -3 16 105
use FILL  FILL_133
timestamp 1713453518
transform 1 0 680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_134
timestamp 1713453518
transform 1 0 600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_135
timestamp 1713453518
transform 1 0 496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_136
timestamp 1713453518
transform 1 0 488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_137
timestamp 1713453518
transform 1 0 264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_138
timestamp 1713453518
transform 1 0 256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_139
timestamp 1713453518
transform 1 0 176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_140
timestamp 1713453518
transform 1 0 168 0 -1 3370
box -8 -3 16 105
use FILL  FILL_141
timestamp 1713453518
transform 1 0 3440 0 1 3170
box -8 -3 16 105
use FILL  FILL_142
timestamp 1713453518
transform 1 0 3432 0 1 3170
box -8 -3 16 105
use FILL  FILL_143
timestamp 1713453518
transform 1 0 3424 0 1 3170
box -8 -3 16 105
use FILL  FILL_144
timestamp 1713453518
transform 1 0 3416 0 1 3170
box -8 -3 16 105
use FILL  FILL_145
timestamp 1713453518
transform 1 0 3408 0 1 3170
box -8 -3 16 105
use FILL  FILL_146
timestamp 1713453518
transform 1 0 3336 0 1 3170
box -8 -3 16 105
use FILL  FILL_147
timestamp 1713453518
transform 1 0 3288 0 1 3170
box -8 -3 16 105
use FILL  FILL_148
timestamp 1713453518
transform 1 0 3280 0 1 3170
box -8 -3 16 105
use FILL  FILL_149
timestamp 1713453518
transform 1 0 3272 0 1 3170
box -8 -3 16 105
use FILL  FILL_150
timestamp 1713453518
transform 1 0 3224 0 1 3170
box -8 -3 16 105
use FILL  FILL_151
timestamp 1713453518
transform 1 0 3216 0 1 3170
box -8 -3 16 105
use FILL  FILL_152
timestamp 1713453518
transform 1 0 3176 0 1 3170
box -8 -3 16 105
use FILL  FILL_153
timestamp 1713453518
transform 1 0 3168 0 1 3170
box -8 -3 16 105
use FILL  FILL_154
timestamp 1713453518
transform 1 0 3160 0 1 3170
box -8 -3 16 105
use FILL  FILL_155
timestamp 1713453518
transform 1 0 3152 0 1 3170
box -8 -3 16 105
use FILL  FILL_156
timestamp 1713453518
transform 1 0 3144 0 1 3170
box -8 -3 16 105
use FILL  FILL_157
timestamp 1713453518
transform 1 0 3112 0 1 3170
box -8 -3 16 105
use FILL  FILL_158
timestamp 1713453518
transform 1 0 3072 0 1 3170
box -8 -3 16 105
use FILL  FILL_159
timestamp 1713453518
transform 1 0 3064 0 1 3170
box -8 -3 16 105
use FILL  FILL_160
timestamp 1713453518
transform 1 0 3056 0 1 3170
box -8 -3 16 105
use FILL  FILL_161
timestamp 1713453518
transform 1 0 3048 0 1 3170
box -8 -3 16 105
use FILL  FILL_162
timestamp 1713453518
transform 1 0 3016 0 1 3170
box -8 -3 16 105
use FILL  FILL_163
timestamp 1713453518
transform 1 0 3008 0 1 3170
box -8 -3 16 105
use FILL  FILL_164
timestamp 1713453518
transform 1 0 3000 0 1 3170
box -8 -3 16 105
use FILL  FILL_165
timestamp 1713453518
transform 1 0 2992 0 1 3170
box -8 -3 16 105
use FILL  FILL_166
timestamp 1713453518
transform 1 0 2984 0 1 3170
box -8 -3 16 105
use FILL  FILL_167
timestamp 1713453518
transform 1 0 2960 0 1 3170
box -8 -3 16 105
use FILL  FILL_168
timestamp 1713453518
transform 1 0 2952 0 1 3170
box -8 -3 16 105
use FILL  FILL_169
timestamp 1713453518
transform 1 0 2944 0 1 3170
box -8 -3 16 105
use FILL  FILL_170
timestamp 1713453518
transform 1 0 2920 0 1 3170
box -8 -3 16 105
use FILL  FILL_171
timestamp 1713453518
transform 1 0 2912 0 1 3170
box -8 -3 16 105
use FILL  FILL_172
timestamp 1713453518
transform 1 0 2904 0 1 3170
box -8 -3 16 105
use FILL  FILL_173
timestamp 1713453518
transform 1 0 2896 0 1 3170
box -8 -3 16 105
use FILL  FILL_174
timestamp 1713453518
transform 1 0 2888 0 1 3170
box -8 -3 16 105
use FILL  FILL_175
timestamp 1713453518
transform 1 0 2880 0 1 3170
box -8 -3 16 105
use FILL  FILL_176
timestamp 1713453518
transform 1 0 2856 0 1 3170
box -8 -3 16 105
use FILL  FILL_177
timestamp 1713453518
transform 1 0 2848 0 1 3170
box -8 -3 16 105
use FILL  FILL_178
timestamp 1713453518
transform 1 0 2816 0 1 3170
box -8 -3 16 105
use FILL  FILL_179
timestamp 1713453518
transform 1 0 2808 0 1 3170
box -8 -3 16 105
use FILL  FILL_180
timestamp 1713453518
transform 1 0 2800 0 1 3170
box -8 -3 16 105
use FILL  FILL_181
timestamp 1713453518
transform 1 0 2792 0 1 3170
box -8 -3 16 105
use FILL  FILL_182
timestamp 1713453518
transform 1 0 2784 0 1 3170
box -8 -3 16 105
use FILL  FILL_183
timestamp 1713453518
transform 1 0 2776 0 1 3170
box -8 -3 16 105
use FILL  FILL_184
timestamp 1713453518
transform 1 0 2768 0 1 3170
box -8 -3 16 105
use FILL  FILL_185
timestamp 1713453518
transform 1 0 2760 0 1 3170
box -8 -3 16 105
use FILL  FILL_186
timestamp 1713453518
transform 1 0 2752 0 1 3170
box -8 -3 16 105
use FILL  FILL_187
timestamp 1713453518
transform 1 0 2704 0 1 3170
box -8 -3 16 105
use FILL  FILL_188
timestamp 1713453518
transform 1 0 2696 0 1 3170
box -8 -3 16 105
use FILL  FILL_189
timestamp 1713453518
transform 1 0 2688 0 1 3170
box -8 -3 16 105
use FILL  FILL_190
timestamp 1713453518
transform 1 0 2680 0 1 3170
box -8 -3 16 105
use FILL  FILL_191
timestamp 1713453518
transform 1 0 2672 0 1 3170
box -8 -3 16 105
use FILL  FILL_192
timestamp 1713453518
transform 1 0 2664 0 1 3170
box -8 -3 16 105
use FILL  FILL_193
timestamp 1713453518
transform 1 0 2656 0 1 3170
box -8 -3 16 105
use FILL  FILL_194
timestamp 1713453518
transform 1 0 2648 0 1 3170
box -8 -3 16 105
use FILL  FILL_195
timestamp 1713453518
transform 1 0 2624 0 1 3170
box -8 -3 16 105
use FILL  FILL_196
timestamp 1713453518
transform 1 0 2616 0 1 3170
box -8 -3 16 105
use FILL  FILL_197
timestamp 1713453518
transform 1 0 2608 0 1 3170
box -8 -3 16 105
use FILL  FILL_198
timestamp 1713453518
transform 1 0 2600 0 1 3170
box -8 -3 16 105
use FILL  FILL_199
timestamp 1713453518
transform 1 0 2568 0 1 3170
box -8 -3 16 105
use FILL  FILL_200
timestamp 1713453518
transform 1 0 2560 0 1 3170
box -8 -3 16 105
use FILL  FILL_201
timestamp 1713453518
transform 1 0 2552 0 1 3170
box -8 -3 16 105
use FILL  FILL_202
timestamp 1713453518
transform 1 0 2544 0 1 3170
box -8 -3 16 105
use FILL  FILL_203
timestamp 1713453518
transform 1 0 2536 0 1 3170
box -8 -3 16 105
use FILL  FILL_204
timestamp 1713453518
transform 1 0 2528 0 1 3170
box -8 -3 16 105
use FILL  FILL_205
timestamp 1713453518
transform 1 0 2520 0 1 3170
box -8 -3 16 105
use FILL  FILL_206
timestamp 1713453518
transform 1 0 2480 0 1 3170
box -8 -3 16 105
use FILL  FILL_207
timestamp 1713453518
transform 1 0 2472 0 1 3170
box -8 -3 16 105
use FILL  FILL_208
timestamp 1713453518
transform 1 0 2464 0 1 3170
box -8 -3 16 105
use FILL  FILL_209
timestamp 1713453518
transform 1 0 2456 0 1 3170
box -8 -3 16 105
use FILL  FILL_210
timestamp 1713453518
transform 1 0 2448 0 1 3170
box -8 -3 16 105
use FILL  FILL_211
timestamp 1713453518
transform 1 0 2440 0 1 3170
box -8 -3 16 105
use FILL  FILL_212
timestamp 1713453518
transform 1 0 2432 0 1 3170
box -8 -3 16 105
use FILL  FILL_213
timestamp 1713453518
transform 1 0 2424 0 1 3170
box -8 -3 16 105
use FILL  FILL_214
timestamp 1713453518
transform 1 0 2416 0 1 3170
box -8 -3 16 105
use FILL  FILL_215
timestamp 1713453518
transform 1 0 2408 0 1 3170
box -8 -3 16 105
use FILL  FILL_216
timestamp 1713453518
transform 1 0 2360 0 1 3170
box -8 -3 16 105
use FILL  FILL_217
timestamp 1713453518
transform 1 0 2352 0 1 3170
box -8 -3 16 105
use FILL  FILL_218
timestamp 1713453518
transform 1 0 2344 0 1 3170
box -8 -3 16 105
use FILL  FILL_219
timestamp 1713453518
transform 1 0 2336 0 1 3170
box -8 -3 16 105
use FILL  FILL_220
timestamp 1713453518
transform 1 0 2328 0 1 3170
box -8 -3 16 105
use FILL  FILL_221
timestamp 1713453518
transform 1 0 2320 0 1 3170
box -8 -3 16 105
use FILL  FILL_222
timestamp 1713453518
transform 1 0 2312 0 1 3170
box -8 -3 16 105
use FILL  FILL_223
timestamp 1713453518
transform 1 0 2304 0 1 3170
box -8 -3 16 105
use FILL  FILL_224
timestamp 1713453518
transform 1 0 2296 0 1 3170
box -8 -3 16 105
use FILL  FILL_225
timestamp 1713453518
transform 1 0 2256 0 1 3170
box -8 -3 16 105
use FILL  FILL_226
timestamp 1713453518
transform 1 0 2248 0 1 3170
box -8 -3 16 105
use FILL  FILL_227
timestamp 1713453518
transform 1 0 2240 0 1 3170
box -8 -3 16 105
use FILL  FILL_228
timestamp 1713453518
transform 1 0 2232 0 1 3170
box -8 -3 16 105
use FILL  FILL_229
timestamp 1713453518
transform 1 0 2224 0 1 3170
box -8 -3 16 105
use FILL  FILL_230
timestamp 1713453518
transform 1 0 2216 0 1 3170
box -8 -3 16 105
use FILL  FILL_231
timestamp 1713453518
transform 1 0 2208 0 1 3170
box -8 -3 16 105
use FILL  FILL_232
timestamp 1713453518
transform 1 0 2200 0 1 3170
box -8 -3 16 105
use FILL  FILL_233
timestamp 1713453518
transform 1 0 2192 0 1 3170
box -8 -3 16 105
use FILL  FILL_234
timestamp 1713453518
transform 1 0 2152 0 1 3170
box -8 -3 16 105
use FILL  FILL_235
timestamp 1713453518
transform 1 0 2144 0 1 3170
box -8 -3 16 105
use FILL  FILL_236
timestamp 1713453518
transform 1 0 2136 0 1 3170
box -8 -3 16 105
use FILL  FILL_237
timestamp 1713453518
transform 1 0 2128 0 1 3170
box -8 -3 16 105
use FILL  FILL_238
timestamp 1713453518
transform 1 0 2120 0 1 3170
box -8 -3 16 105
use FILL  FILL_239
timestamp 1713453518
transform 1 0 2112 0 1 3170
box -8 -3 16 105
use FILL  FILL_240
timestamp 1713453518
transform 1 0 2104 0 1 3170
box -8 -3 16 105
use FILL  FILL_241
timestamp 1713453518
transform 1 0 2096 0 1 3170
box -8 -3 16 105
use FILL  FILL_242
timestamp 1713453518
transform 1 0 2088 0 1 3170
box -8 -3 16 105
use FILL  FILL_243
timestamp 1713453518
transform 1 0 2080 0 1 3170
box -8 -3 16 105
use FILL  FILL_244
timestamp 1713453518
transform 1 0 2032 0 1 3170
box -8 -3 16 105
use FILL  FILL_245
timestamp 1713453518
transform 1 0 2024 0 1 3170
box -8 -3 16 105
use FILL  FILL_246
timestamp 1713453518
transform 1 0 2016 0 1 3170
box -8 -3 16 105
use FILL  FILL_247
timestamp 1713453518
transform 1 0 2008 0 1 3170
box -8 -3 16 105
use FILL  FILL_248
timestamp 1713453518
transform 1 0 2000 0 1 3170
box -8 -3 16 105
use FILL  FILL_249
timestamp 1713453518
transform 1 0 1992 0 1 3170
box -8 -3 16 105
use FILL  FILL_250
timestamp 1713453518
transform 1 0 1984 0 1 3170
box -8 -3 16 105
use FILL  FILL_251
timestamp 1713453518
transform 1 0 1976 0 1 3170
box -8 -3 16 105
use FILL  FILL_252
timestamp 1713453518
transform 1 0 1936 0 1 3170
box -8 -3 16 105
use FILL  FILL_253
timestamp 1713453518
transform 1 0 1928 0 1 3170
box -8 -3 16 105
use FILL  FILL_254
timestamp 1713453518
transform 1 0 1920 0 1 3170
box -8 -3 16 105
use FILL  FILL_255
timestamp 1713453518
transform 1 0 1912 0 1 3170
box -8 -3 16 105
use FILL  FILL_256
timestamp 1713453518
transform 1 0 1904 0 1 3170
box -8 -3 16 105
use FILL  FILL_257
timestamp 1713453518
transform 1 0 1896 0 1 3170
box -8 -3 16 105
use FILL  FILL_258
timestamp 1713453518
transform 1 0 1864 0 1 3170
box -8 -3 16 105
use FILL  FILL_259
timestamp 1713453518
transform 1 0 1856 0 1 3170
box -8 -3 16 105
use FILL  FILL_260
timestamp 1713453518
transform 1 0 1848 0 1 3170
box -8 -3 16 105
use FILL  FILL_261
timestamp 1713453518
transform 1 0 1840 0 1 3170
box -8 -3 16 105
use FILL  FILL_262
timestamp 1713453518
transform 1 0 1832 0 1 3170
box -8 -3 16 105
use FILL  FILL_263
timestamp 1713453518
transform 1 0 1824 0 1 3170
box -8 -3 16 105
use FILL  FILL_264
timestamp 1713453518
transform 1 0 1816 0 1 3170
box -8 -3 16 105
use FILL  FILL_265
timestamp 1713453518
transform 1 0 1808 0 1 3170
box -8 -3 16 105
use FILL  FILL_266
timestamp 1713453518
transform 1 0 1800 0 1 3170
box -8 -3 16 105
use FILL  FILL_267
timestamp 1713453518
transform 1 0 1760 0 1 3170
box -8 -3 16 105
use FILL  FILL_268
timestamp 1713453518
transform 1 0 1752 0 1 3170
box -8 -3 16 105
use FILL  FILL_269
timestamp 1713453518
transform 1 0 1744 0 1 3170
box -8 -3 16 105
use FILL  FILL_270
timestamp 1713453518
transform 1 0 1736 0 1 3170
box -8 -3 16 105
use FILL  FILL_271
timestamp 1713453518
transform 1 0 1728 0 1 3170
box -8 -3 16 105
use FILL  FILL_272
timestamp 1713453518
transform 1 0 1704 0 1 3170
box -8 -3 16 105
use FILL  FILL_273
timestamp 1713453518
transform 1 0 1696 0 1 3170
box -8 -3 16 105
use FILL  FILL_274
timestamp 1713453518
transform 1 0 1688 0 1 3170
box -8 -3 16 105
use FILL  FILL_275
timestamp 1713453518
transform 1 0 1680 0 1 3170
box -8 -3 16 105
use FILL  FILL_276
timestamp 1713453518
transform 1 0 1672 0 1 3170
box -8 -3 16 105
use FILL  FILL_277
timestamp 1713453518
transform 1 0 1664 0 1 3170
box -8 -3 16 105
use FILL  FILL_278
timestamp 1713453518
transform 1 0 1656 0 1 3170
box -8 -3 16 105
use FILL  FILL_279
timestamp 1713453518
transform 1 0 1648 0 1 3170
box -8 -3 16 105
use FILL  FILL_280
timestamp 1713453518
transform 1 0 1600 0 1 3170
box -8 -3 16 105
use FILL  FILL_281
timestamp 1713453518
transform 1 0 1592 0 1 3170
box -8 -3 16 105
use FILL  FILL_282
timestamp 1713453518
transform 1 0 1584 0 1 3170
box -8 -3 16 105
use FILL  FILL_283
timestamp 1713453518
transform 1 0 1576 0 1 3170
box -8 -3 16 105
use FILL  FILL_284
timestamp 1713453518
transform 1 0 1568 0 1 3170
box -8 -3 16 105
use FILL  FILL_285
timestamp 1713453518
transform 1 0 1560 0 1 3170
box -8 -3 16 105
use FILL  FILL_286
timestamp 1713453518
transform 1 0 1552 0 1 3170
box -8 -3 16 105
use FILL  FILL_287
timestamp 1713453518
transform 1 0 1544 0 1 3170
box -8 -3 16 105
use FILL  FILL_288
timestamp 1713453518
transform 1 0 1504 0 1 3170
box -8 -3 16 105
use FILL  FILL_289
timestamp 1713453518
transform 1 0 1496 0 1 3170
box -8 -3 16 105
use FILL  FILL_290
timestamp 1713453518
transform 1 0 1488 0 1 3170
box -8 -3 16 105
use FILL  FILL_291
timestamp 1713453518
transform 1 0 1480 0 1 3170
box -8 -3 16 105
use FILL  FILL_292
timestamp 1713453518
transform 1 0 1472 0 1 3170
box -8 -3 16 105
use FILL  FILL_293
timestamp 1713453518
transform 1 0 1464 0 1 3170
box -8 -3 16 105
use FILL  FILL_294
timestamp 1713453518
transform 1 0 1416 0 1 3170
box -8 -3 16 105
use FILL  FILL_295
timestamp 1713453518
transform 1 0 1408 0 1 3170
box -8 -3 16 105
use FILL  FILL_296
timestamp 1713453518
transform 1 0 1400 0 1 3170
box -8 -3 16 105
use FILL  FILL_297
timestamp 1713453518
transform 1 0 1392 0 1 3170
box -8 -3 16 105
use FILL  FILL_298
timestamp 1713453518
transform 1 0 1368 0 1 3170
box -8 -3 16 105
use FILL  FILL_299
timestamp 1713453518
transform 1 0 1360 0 1 3170
box -8 -3 16 105
use FILL  FILL_300
timestamp 1713453518
transform 1 0 1352 0 1 3170
box -8 -3 16 105
use FILL  FILL_301
timestamp 1713453518
transform 1 0 1344 0 1 3170
box -8 -3 16 105
use FILL  FILL_302
timestamp 1713453518
transform 1 0 1304 0 1 3170
box -8 -3 16 105
use FILL  FILL_303
timestamp 1713453518
transform 1 0 1296 0 1 3170
box -8 -3 16 105
use FILL  FILL_304
timestamp 1713453518
transform 1 0 1288 0 1 3170
box -8 -3 16 105
use FILL  FILL_305
timestamp 1713453518
transform 1 0 1280 0 1 3170
box -8 -3 16 105
use FILL  FILL_306
timestamp 1713453518
transform 1 0 1272 0 1 3170
box -8 -3 16 105
use FILL  FILL_307
timestamp 1713453518
transform 1 0 1240 0 1 3170
box -8 -3 16 105
use FILL  FILL_308
timestamp 1713453518
transform 1 0 1232 0 1 3170
box -8 -3 16 105
use FILL  FILL_309
timestamp 1713453518
transform 1 0 1224 0 1 3170
box -8 -3 16 105
use FILL  FILL_310
timestamp 1713453518
transform 1 0 1192 0 1 3170
box -8 -3 16 105
use FILL  FILL_311
timestamp 1713453518
transform 1 0 1184 0 1 3170
box -8 -3 16 105
use FILL  FILL_312
timestamp 1713453518
transform 1 0 1176 0 1 3170
box -8 -3 16 105
use FILL  FILL_313
timestamp 1713453518
transform 1 0 1168 0 1 3170
box -8 -3 16 105
use FILL  FILL_314
timestamp 1713453518
transform 1 0 1136 0 1 3170
box -8 -3 16 105
use FILL  FILL_315
timestamp 1713453518
transform 1 0 1128 0 1 3170
box -8 -3 16 105
use FILL  FILL_316
timestamp 1713453518
transform 1 0 1120 0 1 3170
box -8 -3 16 105
use FILL  FILL_317
timestamp 1713453518
transform 1 0 1112 0 1 3170
box -8 -3 16 105
use FILL  FILL_318
timestamp 1713453518
transform 1 0 1104 0 1 3170
box -8 -3 16 105
use FILL  FILL_319
timestamp 1713453518
transform 1 0 1064 0 1 3170
box -8 -3 16 105
use FILL  FILL_320
timestamp 1713453518
transform 1 0 1056 0 1 3170
box -8 -3 16 105
use FILL  FILL_321
timestamp 1713453518
transform 1 0 1048 0 1 3170
box -8 -3 16 105
use FILL  FILL_322
timestamp 1713453518
transform 1 0 1040 0 1 3170
box -8 -3 16 105
use FILL  FILL_323
timestamp 1713453518
transform 1 0 1016 0 1 3170
box -8 -3 16 105
use FILL  FILL_324
timestamp 1713453518
transform 1 0 1008 0 1 3170
box -8 -3 16 105
use FILL  FILL_325
timestamp 1713453518
transform 1 0 960 0 1 3170
box -8 -3 16 105
use FILL  FILL_326
timestamp 1713453518
transform 1 0 952 0 1 3170
box -8 -3 16 105
use FILL  FILL_327
timestamp 1713453518
transform 1 0 944 0 1 3170
box -8 -3 16 105
use FILL  FILL_328
timestamp 1713453518
transform 1 0 896 0 1 3170
box -8 -3 16 105
use FILL  FILL_329
timestamp 1713453518
transform 1 0 888 0 1 3170
box -8 -3 16 105
use FILL  FILL_330
timestamp 1713453518
transform 1 0 880 0 1 3170
box -8 -3 16 105
use FILL  FILL_331
timestamp 1713453518
transform 1 0 872 0 1 3170
box -8 -3 16 105
use FILL  FILL_332
timestamp 1713453518
transform 1 0 864 0 1 3170
box -8 -3 16 105
use FILL  FILL_333
timestamp 1713453518
transform 1 0 800 0 1 3170
box -8 -3 16 105
use FILL  FILL_334
timestamp 1713453518
transform 1 0 792 0 1 3170
box -8 -3 16 105
use FILL  FILL_335
timestamp 1713453518
transform 1 0 784 0 1 3170
box -8 -3 16 105
use FILL  FILL_336
timestamp 1713453518
transform 1 0 680 0 1 3170
box -8 -3 16 105
use FILL  FILL_337
timestamp 1713453518
transform 1 0 672 0 1 3170
box -8 -3 16 105
use FILL  FILL_338
timestamp 1713453518
transform 1 0 664 0 1 3170
box -8 -3 16 105
use FILL  FILL_339
timestamp 1713453518
transform 1 0 616 0 1 3170
box -8 -3 16 105
use FILL  FILL_340
timestamp 1713453518
transform 1 0 608 0 1 3170
box -8 -3 16 105
use FILL  FILL_341
timestamp 1713453518
transform 1 0 504 0 1 3170
box -8 -3 16 105
use FILL  FILL_342
timestamp 1713453518
transform 1 0 496 0 1 3170
box -8 -3 16 105
use FILL  FILL_343
timestamp 1713453518
transform 1 0 488 0 1 3170
box -8 -3 16 105
use FILL  FILL_344
timestamp 1713453518
transform 1 0 480 0 1 3170
box -8 -3 16 105
use FILL  FILL_345
timestamp 1713453518
transform 1 0 472 0 1 3170
box -8 -3 16 105
use FILL  FILL_346
timestamp 1713453518
transform 1 0 416 0 1 3170
box -8 -3 16 105
use FILL  FILL_347
timestamp 1713453518
transform 1 0 408 0 1 3170
box -8 -3 16 105
use FILL  FILL_348
timestamp 1713453518
transform 1 0 400 0 1 3170
box -8 -3 16 105
use FILL  FILL_349
timestamp 1713453518
transform 1 0 392 0 1 3170
box -8 -3 16 105
use FILL  FILL_350
timestamp 1713453518
transform 1 0 288 0 1 3170
box -8 -3 16 105
use FILL  FILL_351
timestamp 1713453518
transform 1 0 280 0 1 3170
box -8 -3 16 105
use FILL  FILL_352
timestamp 1713453518
transform 1 0 272 0 1 3170
box -8 -3 16 105
use FILL  FILL_353
timestamp 1713453518
transform 1 0 264 0 1 3170
box -8 -3 16 105
use FILL  FILL_354
timestamp 1713453518
transform 1 0 160 0 1 3170
box -8 -3 16 105
use FILL  FILL_355
timestamp 1713453518
transform 1 0 152 0 1 3170
box -8 -3 16 105
use FILL  FILL_356
timestamp 1713453518
transform 1 0 144 0 1 3170
box -8 -3 16 105
use FILL  FILL_357
timestamp 1713453518
transform 1 0 136 0 1 3170
box -8 -3 16 105
use FILL  FILL_358
timestamp 1713453518
transform 1 0 128 0 1 3170
box -8 -3 16 105
use FILL  FILL_359
timestamp 1713453518
transform 1 0 120 0 1 3170
box -8 -3 16 105
use FILL  FILL_360
timestamp 1713453518
transform 1 0 112 0 1 3170
box -8 -3 16 105
use FILL  FILL_361
timestamp 1713453518
transform 1 0 104 0 1 3170
box -8 -3 16 105
use FILL  FILL_362
timestamp 1713453518
transform 1 0 96 0 1 3170
box -8 -3 16 105
use FILL  FILL_363
timestamp 1713453518
transform 1 0 88 0 1 3170
box -8 -3 16 105
use FILL  FILL_364
timestamp 1713453518
transform 1 0 80 0 1 3170
box -8 -3 16 105
use FILL  FILL_365
timestamp 1713453518
transform 1 0 72 0 1 3170
box -8 -3 16 105
use FILL  FILL_366
timestamp 1713453518
transform 1 0 3440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_367
timestamp 1713453518
transform 1 0 3376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_368
timestamp 1713453518
transform 1 0 3288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_369
timestamp 1713453518
transform 1 0 3224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_370
timestamp 1713453518
transform 1 0 3184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_371
timestamp 1713453518
transform 1 0 3176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_372
timestamp 1713453518
transform 1 0 3168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_373
timestamp 1713453518
transform 1 0 3160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_374
timestamp 1713453518
transform 1 0 3152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_375
timestamp 1713453518
transform 1 0 3088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_376
timestamp 1713453518
transform 1 0 3080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_377
timestamp 1713453518
transform 1 0 3072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_378
timestamp 1713453518
transform 1 0 3064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_379
timestamp 1713453518
transform 1 0 3056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_380
timestamp 1713453518
transform 1 0 3048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_381
timestamp 1713453518
transform 1 0 3000 0 -1 3170
box -8 -3 16 105
use FILL  FILL_382
timestamp 1713453518
transform 1 0 2992 0 -1 3170
box -8 -3 16 105
use FILL  FILL_383
timestamp 1713453518
transform 1 0 2984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_384
timestamp 1713453518
transform 1 0 2976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_385
timestamp 1713453518
transform 1 0 2968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_386
timestamp 1713453518
transform 1 0 2960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_387
timestamp 1713453518
transform 1 0 2912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_388
timestamp 1713453518
transform 1 0 2904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_389
timestamp 1713453518
transform 1 0 2896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_390
timestamp 1713453518
transform 1 0 2888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_391
timestamp 1713453518
transform 1 0 2880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_392
timestamp 1713453518
transform 1 0 2872 0 -1 3170
box -8 -3 16 105
use FILL  FILL_393
timestamp 1713453518
transform 1 0 2864 0 -1 3170
box -8 -3 16 105
use FILL  FILL_394
timestamp 1713453518
transform 1 0 2824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_395
timestamp 1713453518
transform 1 0 2816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_396
timestamp 1713453518
transform 1 0 2808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_397
timestamp 1713453518
transform 1 0 2800 0 -1 3170
box -8 -3 16 105
use FILL  FILL_398
timestamp 1713453518
transform 1 0 2760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_399
timestamp 1713453518
transform 1 0 2752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_400
timestamp 1713453518
transform 1 0 2744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_401
timestamp 1713453518
transform 1 0 2736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_402
timestamp 1713453518
transform 1 0 2728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_403
timestamp 1713453518
transform 1 0 2720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_404
timestamp 1713453518
transform 1 0 2712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_405
timestamp 1713453518
transform 1 0 2672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_406
timestamp 1713453518
transform 1 0 2664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_407
timestamp 1713453518
transform 1 0 2656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_408
timestamp 1713453518
transform 1 0 2648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_409
timestamp 1713453518
transform 1 0 2640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_410
timestamp 1713453518
transform 1 0 2600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_411
timestamp 1713453518
transform 1 0 2592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_412
timestamp 1713453518
transform 1 0 2584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_413
timestamp 1713453518
transform 1 0 2576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_414
timestamp 1713453518
transform 1 0 2568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_415
timestamp 1713453518
transform 1 0 2560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_416
timestamp 1713453518
transform 1 0 2552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_417
timestamp 1713453518
transform 1 0 2544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_418
timestamp 1713453518
transform 1 0 2504 0 -1 3170
box -8 -3 16 105
use FILL  FILL_419
timestamp 1713453518
transform 1 0 2496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_420
timestamp 1713453518
transform 1 0 2488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_421
timestamp 1713453518
transform 1 0 2480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_422
timestamp 1713453518
transform 1 0 2472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_423
timestamp 1713453518
transform 1 0 2464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_424
timestamp 1713453518
transform 1 0 2440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_425
timestamp 1713453518
transform 1 0 2432 0 -1 3170
box -8 -3 16 105
use FILL  FILL_426
timestamp 1713453518
transform 1 0 2424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_427
timestamp 1713453518
transform 1 0 2392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_428
timestamp 1713453518
transform 1 0 2384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_429
timestamp 1713453518
transform 1 0 2376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_430
timestamp 1713453518
transform 1 0 2368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_431
timestamp 1713453518
transform 1 0 2360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_432
timestamp 1713453518
transform 1 0 2352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_433
timestamp 1713453518
transform 1 0 2344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_434
timestamp 1713453518
transform 1 0 2336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_435
timestamp 1713453518
transform 1 0 2288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_436
timestamp 1713453518
transform 1 0 2280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_437
timestamp 1713453518
transform 1 0 2272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_438
timestamp 1713453518
transform 1 0 2264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_439
timestamp 1713453518
transform 1 0 2256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_440
timestamp 1713453518
transform 1 0 2248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_441
timestamp 1713453518
transform 1 0 2240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_442
timestamp 1713453518
transform 1 0 2208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_443
timestamp 1713453518
transform 1 0 2200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_444
timestamp 1713453518
transform 1 0 2192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_445
timestamp 1713453518
transform 1 0 2184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_446
timestamp 1713453518
transform 1 0 2176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_447
timestamp 1713453518
transform 1 0 2168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_448
timestamp 1713453518
transform 1 0 2128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_449
timestamp 1713453518
transform 1 0 2120 0 -1 3170
box -8 -3 16 105
use FILL  FILL_450
timestamp 1713453518
transform 1 0 2112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_451
timestamp 1713453518
transform 1 0 2104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_452
timestamp 1713453518
transform 1 0 2096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_453
timestamp 1713453518
transform 1 0 2088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_454
timestamp 1713453518
transform 1 0 2080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_455
timestamp 1713453518
transform 1 0 2048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_456
timestamp 1713453518
transform 1 0 2040 0 -1 3170
box -8 -3 16 105
use FILL  FILL_457
timestamp 1713453518
transform 1 0 2032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_458
timestamp 1713453518
transform 1 0 2024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_459
timestamp 1713453518
transform 1 0 2016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_460
timestamp 1713453518
transform 1 0 2008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_461
timestamp 1713453518
transform 1 0 1968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_462
timestamp 1713453518
transform 1 0 1960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_463
timestamp 1713453518
transform 1 0 1952 0 -1 3170
box -8 -3 16 105
use FILL  FILL_464
timestamp 1713453518
transform 1 0 1944 0 -1 3170
box -8 -3 16 105
use FILL  FILL_465
timestamp 1713453518
transform 1 0 1936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_466
timestamp 1713453518
transform 1 0 1928 0 -1 3170
box -8 -3 16 105
use FILL  FILL_467
timestamp 1713453518
transform 1 0 1920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_468
timestamp 1713453518
transform 1 0 1912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_469
timestamp 1713453518
transform 1 0 1864 0 -1 3170
box -8 -3 16 105
use FILL  FILL_470
timestamp 1713453518
transform 1 0 1856 0 -1 3170
box -8 -3 16 105
use FILL  FILL_471
timestamp 1713453518
transform 1 0 1848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_472
timestamp 1713453518
transform 1 0 1840 0 -1 3170
box -8 -3 16 105
use FILL  FILL_473
timestamp 1713453518
transform 1 0 1832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_474
timestamp 1713453518
transform 1 0 1824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_475
timestamp 1713453518
transform 1 0 1816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_476
timestamp 1713453518
transform 1 0 1808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_477
timestamp 1713453518
transform 1 0 1800 0 -1 3170
box -8 -3 16 105
use FILL  FILL_478
timestamp 1713453518
transform 1 0 1752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_479
timestamp 1713453518
transform 1 0 1744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_480
timestamp 1713453518
transform 1 0 1736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_481
timestamp 1713453518
transform 1 0 1728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_482
timestamp 1713453518
transform 1 0 1720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_483
timestamp 1713453518
transform 1 0 1712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_484
timestamp 1713453518
transform 1 0 1704 0 -1 3170
box -8 -3 16 105
use FILL  FILL_485
timestamp 1713453518
transform 1 0 1672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_486
timestamp 1713453518
transform 1 0 1664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_487
timestamp 1713453518
transform 1 0 1656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_488
timestamp 1713453518
transform 1 0 1648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_489
timestamp 1713453518
transform 1 0 1624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_490
timestamp 1713453518
transform 1 0 1616 0 -1 3170
box -8 -3 16 105
use FILL  FILL_491
timestamp 1713453518
transform 1 0 1608 0 -1 3170
box -8 -3 16 105
use FILL  FILL_492
timestamp 1713453518
transform 1 0 1584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_493
timestamp 1713453518
transform 1 0 1576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_494
timestamp 1713453518
transform 1 0 1568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_495
timestamp 1713453518
transform 1 0 1560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_496
timestamp 1713453518
transform 1 0 1552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_497
timestamp 1713453518
transform 1 0 1544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_498
timestamp 1713453518
transform 1 0 1504 0 -1 3170
box -8 -3 16 105
use FILL  FILL_499
timestamp 1713453518
transform 1 0 1496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_500
timestamp 1713453518
transform 1 0 1488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_501
timestamp 1713453518
transform 1 0 1480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_502
timestamp 1713453518
transform 1 0 1472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_503
timestamp 1713453518
transform 1 0 1432 0 -1 3170
box -8 -3 16 105
use FILL  FILL_504
timestamp 1713453518
transform 1 0 1424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_505
timestamp 1713453518
transform 1 0 1400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_506
timestamp 1713453518
transform 1 0 1392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_507
timestamp 1713453518
transform 1 0 1352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_508
timestamp 1713453518
transform 1 0 1344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_509
timestamp 1713453518
transform 1 0 1336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_510
timestamp 1713453518
transform 1 0 1328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_511
timestamp 1713453518
transform 1 0 1272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_512
timestamp 1713453518
transform 1 0 1264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_513
timestamp 1713453518
transform 1 0 1256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_514
timestamp 1713453518
transform 1 0 1248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_515
timestamp 1713453518
transform 1 0 1240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_516
timestamp 1713453518
transform 1 0 1232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_517
timestamp 1713453518
transform 1 0 1176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_518
timestamp 1713453518
transform 1 0 1168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_519
timestamp 1713453518
transform 1 0 1160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_520
timestamp 1713453518
transform 1 0 1152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_521
timestamp 1713453518
transform 1 0 1144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_522
timestamp 1713453518
transform 1 0 1088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_523
timestamp 1713453518
transform 1 0 1080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_524
timestamp 1713453518
transform 1 0 976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_525
timestamp 1713453518
transform 1 0 968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_526
timestamp 1713453518
transform 1 0 960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_527
timestamp 1713453518
transform 1 0 952 0 -1 3170
box -8 -3 16 105
use FILL  FILL_528
timestamp 1713453518
transform 1 0 856 0 -1 3170
box -8 -3 16 105
use FILL  FILL_529
timestamp 1713453518
transform 1 0 848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_530
timestamp 1713453518
transform 1 0 840 0 -1 3170
box -8 -3 16 105
use FILL  FILL_531
timestamp 1713453518
transform 1 0 832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_532
timestamp 1713453518
transform 1 0 728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_533
timestamp 1713453518
transform 1 0 720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_534
timestamp 1713453518
transform 1 0 712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_535
timestamp 1713453518
transform 1 0 704 0 -1 3170
box -8 -3 16 105
use FILL  FILL_536
timestamp 1713453518
transform 1 0 696 0 -1 3170
box -8 -3 16 105
use FILL  FILL_537
timestamp 1713453518
transform 1 0 632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_538
timestamp 1713453518
transform 1 0 624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_539
timestamp 1713453518
transform 1 0 584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_540
timestamp 1713453518
transform 1 0 576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_541
timestamp 1713453518
transform 1 0 568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_542
timestamp 1713453518
transform 1 0 560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_543
timestamp 1713453518
transform 1 0 512 0 -1 3170
box -8 -3 16 105
use FILL  FILL_544
timestamp 1713453518
transform 1 0 504 0 -1 3170
box -8 -3 16 105
use FILL  FILL_545
timestamp 1713453518
transform 1 0 496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_546
timestamp 1713453518
transform 1 0 488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_547
timestamp 1713453518
transform 1 0 480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_548
timestamp 1713453518
transform 1 0 376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_549
timestamp 1713453518
transform 1 0 368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_550
timestamp 1713453518
transform 1 0 360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_551
timestamp 1713453518
transform 1 0 352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_552
timestamp 1713453518
transform 1 0 344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_553
timestamp 1713453518
transform 1 0 336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_554
timestamp 1713453518
transform 1 0 328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_555
timestamp 1713453518
transform 1 0 320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_556
timestamp 1713453518
transform 1 0 288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_557
timestamp 1713453518
transform 1 0 280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_558
timestamp 1713453518
transform 1 0 224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_559
timestamp 1713453518
transform 1 0 216 0 -1 3170
box -8 -3 16 105
use FILL  FILL_560
timestamp 1713453518
transform 1 0 208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_561
timestamp 1713453518
transform 1 0 200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_562
timestamp 1713453518
transform 1 0 192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_563
timestamp 1713453518
transform 1 0 184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_564
timestamp 1713453518
transform 1 0 176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_565
timestamp 1713453518
transform 1 0 72 0 -1 3170
box -8 -3 16 105
use FILL  FILL_566
timestamp 1713453518
transform 1 0 3440 0 1 2970
box -8 -3 16 105
use FILL  FILL_567
timestamp 1713453518
transform 1 0 3432 0 1 2970
box -8 -3 16 105
use FILL  FILL_568
timestamp 1713453518
transform 1 0 3344 0 1 2970
box -8 -3 16 105
use FILL  FILL_569
timestamp 1713453518
transform 1 0 3336 0 1 2970
box -8 -3 16 105
use FILL  FILL_570
timestamp 1713453518
transform 1 0 3328 0 1 2970
box -8 -3 16 105
use FILL  FILL_571
timestamp 1713453518
transform 1 0 3296 0 1 2970
box -8 -3 16 105
use FILL  FILL_572
timestamp 1713453518
transform 1 0 3288 0 1 2970
box -8 -3 16 105
use FILL  FILL_573
timestamp 1713453518
transform 1 0 3248 0 1 2970
box -8 -3 16 105
use FILL  FILL_574
timestamp 1713453518
transform 1 0 3240 0 1 2970
box -8 -3 16 105
use FILL  FILL_575
timestamp 1713453518
transform 1 0 3232 0 1 2970
box -8 -3 16 105
use FILL  FILL_576
timestamp 1713453518
transform 1 0 3192 0 1 2970
box -8 -3 16 105
use FILL  FILL_577
timestamp 1713453518
transform 1 0 3184 0 1 2970
box -8 -3 16 105
use FILL  FILL_578
timestamp 1713453518
transform 1 0 3176 0 1 2970
box -8 -3 16 105
use FILL  FILL_579
timestamp 1713453518
transform 1 0 3144 0 1 2970
box -8 -3 16 105
use FILL  FILL_580
timestamp 1713453518
transform 1 0 3136 0 1 2970
box -8 -3 16 105
use FILL  FILL_581
timestamp 1713453518
transform 1 0 3128 0 1 2970
box -8 -3 16 105
use FILL  FILL_582
timestamp 1713453518
transform 1 0 3120 0 1 2970
box -8 -3 16 105
use FILL  FILL_583
timestamp 1713453518
transform 1 0 3112 0 1 2970
box -8 -3 16 105
use FILL  FILL_584
timestamp 1713453518
transform 1 0 3056 0 1 2970
box -8 -3 16 105
use FILL  FILL_585
timestamp 1713453518
transform 1 0 3048 0 1 2970
box -8 -3 16 105
use FILL  FILL_586
timestamp 1713453518
transform 1 0 3040 0 1 2970
box -8 -3 16 105
use FILL  FILL_587
timestamp 1713453518
transform 1 0 3032 0 1 2970
box -8 -3 16 105
use FILL  FILL_588
timestamp 1713453518
transform 1 0 3024 0 1 2970
box -8 -3 16 105
use FILL  FILL_589
timestamp 1713453518
transform 1 0 2992 0 1 2970
box -8 -3 16 105
use FILL  FILL_590
timestamp 1713453518
transform 1 0 2984 0 1 2970
box -8 -3 16 105
use FILL  FILL_591
timestamp 1713453518
transform 1 0 2944 0 1 2970
box -8 -3 16 105
use FILL  FILL_592
timestamp 1713453518
transform 1 0 2936 0 1 2970
box -8 -3 16 105
use FILL  FILL_593
timestamp 1713453518
transform 1 0 2928 0 1 2970
box -8 -3 16 105
use FILL  FILL_594
timestamp 1713453518
transform 1 0 2920 0 1 2970
box -8 -3 16 105
use FILL  FILL_595
timestamp 1713453518
transform 1 0 2912 0 1 2970
box -8 -3 16 105
use FILL  FILL_596
timestamp 1713453518
transform 1 0 2904 0 1 2970
box -8 -3 16 105
use FILL  FILL_597
timestamp 1713453518
transform 1 0 2832 0 1 2970
box -8 -3 16 105
use FILL  FILL_598
timestamp 1713453518
transform 1 0 2824 0 1 2970
box -8 -3 16 105
use FILL  FILL_599
timestamp 1713453518
transform 1 0 2816 0 1 2970
box -8 -3 16 105
use FILL  FILL_600
timestamp 1713453518
transform 1 0 2808 0 1 2970
box -8 -3 16 105
use FILL  FILL_601
timestamp 1713453518
transform 1 0 2800 0 1 2970
box -8 -3 16 105
use FILL  FILL_602
timestamp 1713453518
transform 1 0 2792 0 1 2970
box -8 -3 16 105
use FILL  FILL_603
timestamp 1713453518
transform 1 0 2768 0 1 2970
box -8 -3 16 105
use FILL  FILL_604
timestamp 1713453518
transform 1 0 2760 0 1 2970
box -8 -3 16 105
use FILL  FILL_605
timestamp 1713453518
transform 1 0 2720 0 1 2970
box -8 -3 16 105
use FILL  FILL_606
timestamp 1713453518
transform 1 0 2712 0 1 2970
box -8 -3 16 105
use FILL  FILL_607
timestamp 1713453518
transform 1 0 2704 0 1 2970
box -8 -3 16 105
use FILL  FILL_608
timestamp 1713453518
transform 1 0 2696 0 1 2970
box -8 -3 16 105
use FILL  FILL_609
timestamp 1713453518
transform 1 0 2688 0 1 2970
box -8 -3 16 105
use FILL  FILL_610
timestamp 1713453518
transform 1 0 2680 0 1 2970
box -8 -3 16 105
use FILL  FILL_611
timestamp 1713453518
transform 1 0 2672 0 1 2970
box -8 -3 16 105
use FILL  FILL_612
timestamp 1713453518
transform 1 0 2664 0 1 2970
box -8 -3 16 105
use FILL  FILL_613
timestamp 1713453518
transform 1 0 2656 0 1 2970
box -8 -3 16 105
use FILL  FILL_614
timestamp 1713453518
transform 1 0 2608 0 1 2970
box -8 -3 16 105
use FILL  FILL_615
timestamp 1713453518
transform 1 0 2600 0 1 2970
box -8 -3 16 105
use FILL  FILL_616
timestamp 1713453518
transform 1 0 2592 0 1 2970
box -8 -3 16 105
use FILL  FILL_617
timestamp 1713453518
transform 1 0 2584 0 1 2970
box -8 -3 16 105
use FILL  FILL_618
timestamp 1713453518
transform 1 0 2576 0 1 2970
box -8 -3 16 105
use FILL  FILL_619
timestamp 1713453518
transform 1 0 2568 0 1 2970
box -8 -3 16 105
use FILL  FILL_620
timestamp 1713453518
transform 1 0 2560 0 1 2970
box -8 -3 16 105
use FILL  FILL_621
timestamp 1713453518
transform 1 0 2552 0 1 2970
box -8 -3 16 105
use FILL  FILL_622
timestamp 1713453518
transform 1 0 2520 0 1 2970
box -8 -3 16 105
use FILL  FILL_623
timestamp 1713453518
transform 1 0 2512 0 1 2970
box -8 -3 16 105
use FILL  FILL_624
timestamp 1713453518
transform 1 0 2504 0 1 2970
box -8 -3 16 105
use FILL  FILL_625
timestamp 1713453518
transform 1 0 2496 0 1 2970
box -8 -3 16 105
use FILL  FILL_626
timestamp 1713453518
transform 1 0 2488 0 1 2970
box -8 -3 16 105
use FILL  FILL_627
timestamp 1713453518
transform 1 0 2480 0 1 2970
box -8 -3 16 105
use FILL  FILL_628
timestamp 1713453518
transform 1 0 2448 0 1 2970
box -8 -3 16 105
use FILL  FILL_629
timestamp 1713453518
transform 1 0 2440 0 1 2970
box -8 -3 16 105
use FILL  FILL_630
timestamp 1713453518
transform 1 0 2432 0 1 2970
box -8 -3 16 105
use FILL  FILL_631
timestamp 1713453518
transform 1 0 2424 0 1 2970
box -8 -3 16 105
use FILL  FILL_632
timestamp 1713453518
transform 1 0 2416 0 1 2970
box -8 -3 16 105
use FILL  FILL_633
timestamp 1713453518
transform 1 0 2384 0 1 2970
box -8 -3 16 105
use FILL  FILL_634
timestamp 1713453518
transform 1 0 2376 0 1 2970
box -8 -3 16 105
use FILL  FILL_635
timestamp 1713453518
transform 1 0 2368 0 1 2970
box -8 -3 16 105
use FILL  FILL_636
timestamp 1713453518
transform 1 0 2360 0 1 2970
box -8 -3 16 105
use FILL  FILL_637
timestamp 1713453518
transform 1 0 2352 0 1 2970
box -8 -3 16 105
use FILL  FILL_638
timestamp 1713453518
transform 1 0 2344 0 1 2970
box -8 -3 16 105
use FILL  FILL_639
timestamp 1713453518
transform 1 0 2336 0 1 2970
box -8 -3 16 105
use FILL  FILL_640
timestamp 1713453518
transform 1 0 2288 0 1 2970
box -8 -3 16 105
use FILL  FILL_641
timestamp 1713453518
transform 1 0 2280 0 1 2970
box -8 -3 16 105
use FILL  FILL_642
timestamp 1713453518
transform 1 0 2272 0 1 2970
box -8 -3 16 105
use FILL  FILL_643
timestamp 1713453518
transform 1 0 2264 0 1 2970
box -8 -3 16 105
use FILL  FILL_644
timestamp 1713453518
transform 1 0 2256 0 1 2970
box -8 -3 16 105
use FILL  FILL_645
timestamp 1713453518
transform 1 0 2248 0 1 2970
box -8 -3 16 105
use FILL  FILL_646
timestamp 1713453518
transform 1 0 2240 0 1 2970
box -8 -3 16 105
use FILL  FILL_647
timestamp 1713453518
transform 1 0 2232 0 1 2970
box -8 -3 16 105
use FILL  FILL_648
timestamp 1713453518
transform 1 0 2224 0 1 2970
box -8 -3 16 105
use FILL  FILL_649
timestamp 1713453518
transform 1 0 2184 0 1 2970
box -8 -3 16 105
use FILL  FILL_650
timestamp 1713453518
transform 1 0 2176 0 1 2970
box -8 -3 16 105
use FILL  FILL_651
timestamp 1713453518
transform 1 0 2168 0 1 2970
box -8 -3 16 105
use FILL  FILL_652
timestamp 1713453518
transform 1 0 2160 0 1 2970
box -8 -3 16 105
use FILL  FILL_653
timestamp 1713453518
transform 1 0 2152 0 1 2970
box -8 -3 16 105
use FILL  FILL_654
timestamp 1713453518
transform 1 0 2144 0 1 2970
box -8 -3 16 105
use FILL  FILL_655
timestamp 1713453518
transform 1 0 2136 0 1 2970
box -8 -3 16 105
use FILL  FILL_656
timestamp 1713453518
transform 1 0 2128 0 1 2970
box -8 -3 16 105
use FILL  FILL_657
timestamp 1713453518
transform 1 0 2120 0 1 2970
box -8 -3 16 105
use FILL  FILL_658
timestamp 1713453518
transform 1 0 2072 0 1 2970
box -8 -3 16 105
use FILL  FILL_659
timestamp 1713453518
transform 1 0 2064 0 1 2970
box -8 -3 16 105
use FILL  FILL_660
timestamp 1713453518
transform 1 0 2056 0 1 2970
box -8 -3 16 105
use FILL  FILL_661
timestamp 1713453518
transform 1 0 2048 0 1 2970
box -8 -3 16 105
use FILL  FILL_662
timestamp 1713453518
transform 1 0 2040 0 1 2970
box -8 -3 16 105
use FILL  FILL_663
timestamp 1713453518
transform 1 0 2032 0 1 2970
box -8 -3 16 105
use FILL  FILL_664
timestamp 1713453518
transform 1 0 2024 0 1 2970
box -8 -3 16 105
use FILL  FILL_665
timestamp 1713453518
transform 1 0 2016 0 1 2970
box -8 -3 16 105
use FILL  FILL_666
timestamp 1713453518
transform 1 0 1984 0 1 2970
box -8 -3 16 105
use FILL  FILL_667
timestamp 1713453518
transform 1 0 1976 0 1 2970
box -8 -3 16 105
use FILL  FILL_668
timestamp 1713453518
transform 1 0 1968 0 1 2970
box -8 -3 16 105
use FILL  FILL_669
timestamp 1713453518
transform 1 0 1960 0 1 2970
box -8 -3 16 105
use FILL  FILL_670
timestamp 1713453518
transform 1 0 1952 0 1 2970
box -8 -3 16 105
use FILL  FILL_671
timestamp 1713453518
transform 1 0 1944 0 1 2970
box -8 -3 16 105
use FILL  FILL_672
timestamp 1713453518
transform 1 0 1912 0 1 2970
box -8 -3 16 105
use FILL  FILL_673
timestamp 1713453518
transform 1 0 1904 0 1 2970
box -8 -3 16 105
use FILL  FILL_674
timestamp 1713453518
transform 1 0 1896 0 1 2970
box -8 -3 16 105
use FILL  FILL_675
timestamp 1713453518
transform 1 0 1888 0 1 2970
box -8 -3 16 105
use FILL  FILL_676
timestamp 1713453518
transform 1 0 1880 0 1 2970
box -8 -3 16 105
use FILL  FILL_677
timestamp 1713453518
transform 1 0 1872 0 1 2970
box -8 -3 16 105
use FILL  FILL_678
timestamp 1713453518
transform 1 0 1848 0 1 2970
box -8 -3 16 105
use FILL  FILL_679
timestamp 1713453518
transform 1 0 1840 0 1 2970
box -8 -3 16 105
use FILL  FILL_680
timestamp 1713453518
transform 1 0 1832 0 1 2970
box -8 -3 16 105
use FILL  FILL_681
timestamp 1713453518
transform 1 0 1824 0 1 2970
box -8 -3 16 105
use FILL  FILL_682
timestamp 1713453518
transform 1 0 1816 0 1 2970
box -8 -3 16 105
use FILL  FILL_683
timestamp 1713453518
transform 1 0 1808 0 1 2970
box -8 -3 16 105
use FILL  FILL_684
timestamp 1713453518
transform 1 0 1768 0 1 2970
box -8 -3 16 105
use FILL  FILL_685
timestamp 1713453518
transform 1 0 1760 0 1 2970
box -8 -3 16 105
use FILL  FILL_686
timestamp 1713453518
transform 1 0 1752 0 1 2970
box -8 -3 16 105
use FILL  FILL_687
timestamp 1713453518
transform 1 0 1744 0 1 2970
box -8 -3 16 105
use FILL  FILL_688
timestamp 1713453518
transform 1 0 1736 0 1 2970
box -8 -3 16 105
use FILL  FILL_689
timestamp 1713453518
transform 1 0 1728 0 1 2970
box -8 -3 16 105
use FILL  FILL_690
timestamp 1713453518
transform 1 0 1720 0 1 2970
box -8 -3 16 105
use FILL  FILL_691
timestamp 1713453518
transform 1 0 1712 0 1 2970
box -8 -3 16 105
use FILL  FILL_692
timestamp 1713453518
transform 1 0 1704 0 1 2970
box -8 -3 16 105
use FILL  FILL_693
timestamp 1713453518
transform 1 0 1656 0 1 2970
box -8 -3 16 105
use FILL  FILL_694
timestamp 1713453518
transform 1 0 1648 0 1 2970
box -8 -3 16 105
use FILL  FILL_695
timestamp 1713453518
transform 1 0 1640 0 1 2970
box -8 -3 16 105
use FILL  FILL_696
timestamp 1713453518
transform 1 0 1632 0 1 2970
box -8 -3 16 105
use FILL  FILL_697
timestamp 1713453518
transform 1 0 1624 0 1 2970
box -8 -3 16 105
use FILL  FILL_698
timestamp 1713453518
transform 1 0 1616 0 1 2970
box -8 -3 16 105
use FILL  FILL_699
timestamp 1713453518
transform 1 0 1608 0 1 2970
box -8 -3 16 105
use FILL  FILL_700
timestamp 1713453518
transform 1 0 1600 0 1 2970
box -8 -3 16 105
use FILL  FILL_701
timestamp 1713453518
transform 1 0 1560 0 1 2970
box -8 -3 16 105
use FILL  FILL_702
timestamp 1713453518
transform 1 0 1552 0 1 2970
box -8 -3 16 105
use FILL  FILL_703
timestamp 1713453518
transform 1 0 1544 0 1 2970
box -8 -3 16 105
use FILL  FILL_704
timestamp 1713453518
transform 1 0 1536 0 1 2970
box -8 -3 16 105
use FILL  FILL_705
timestamp 1713453518
transform 1 0 1496 0 1 2970
box -8 -3 16 105
use FILL  FILL_706
timestamp 1713453518
transform 1 0 1488 0 1 2970
box -8 -3 16 105
use FILL  FILL_707
timestamp 1713453518
transform 1 0 1480 0 1 2970
box -8 -3 16 105
use FILL  FILL_708
timestamp 1713453518
transform 1 0 1472 0 1 2970
box -8 -3 16 105
use FILL  FILL_709
timestamp 1713453518
transform 1 0 1464 0 1 2970
box -8 -3 16 105
use FILL  FILL_710
timestamp 1713453518
transform 1 0 1424 0 1 2970
box -8 -3 16 105
use FILL  FILL_711
timestamp 1713453518
transform 1 0 1416 0 1 2970
box -8 -3 16 105
use FILL  FILL_712
timestamp 1713453518
transform 1 0 1408 0 1 2970
box -8 -3 16 105
use FILL  FILL_713
timestamp 1713453518
transform 1 0 1400 0 1 2970
box -8 -3 16 105
use FILL  FILL_714
timestamp 1713453518
transform 1 0 1392 0 1 2970
box -8 -3 16 105
use FILL  FILL_715
timestamp 1713453518
transform 1 0 1352 0 1 2970
box -8 -3 16 105
use FILL  FILL_716
timestamp 1713453518
transform 1 0 1344 0 1 2970
box -8 -3 16 105
use FILL  FILL_717
timestamp 1713453518
transform 1 0 1336 0 1 2970
box -8 -3 16 105
use FILL  FILL_718
timestamp 1713453518
transform 1 0 1328 0 1 2970
box -8 -3 16 105
use FILL  FILL_719
timestamp 1713453518
transform 1 0 1288 0 1 2970
box -8 -3 16 105
use FILL  FILL_720
timestamp 1713453518
transform 1 0 1280 0 1 2970
box -8 -3 16 105
use FILL  FILL_721
timestamp 1713453518
transform 1 0 1272 0 1 2970
box -8 -3 16 105
use FILL  FILL_722
timestamp 1713453518
transform 1 0 1240 0 1 2970
box -8 -3 16 105
use FILL  FILL_723
timestamp 1713453518
transform 1 0 1232 0 1 2970
box -8 -3 16 105
use FILL  FILL_724
timestamp 1713453518
transform 1 0 1224 0 1 2970
box -8 -3 16 105
use FILL  FILL_725
timestamp 1713453518
transform 1 0 1192 0 1 2970
box -8 -3 16 105
use FILL  FILL_726
timestamp 1713453518
transform 1 0 1184 0 1 2970
box -8 -3 16 105
use FILL  FILL_727
timestamp 1713453518
transform 1 0 1176 0 1 2970
box -8 -3 16 105
use FILL  FILL_728
timestamp 1713453518
transform 1 0 1168 0 1 2970
box -8 -3 16 105
use FILL  FILL_729
timestamp 1713453518
transform 1 0 1160 0 1 2970
box -8 -3 16 105
use FILL  FILL_730
timestamp 1713453518
transform 1 0 1104 0 1 2970
box -8 -3 16 105
use FILL  FILL_731
timestamp 1713453518
transform 1 0 1096 0 1 2970
box -8 -3 16 105
use FILL  FILL_732
timestamp 1713453518
transform 1 0 1088 0 1 2970
box -8 -3 16 105
use FILL  FILL_733
timestamp 1713453518
transform 1 0 1080 0 1 2970
box -8 -3 16 105
use FILL  FILL_734
timestamp 1713453518
transform 1 0 1072 0 1 2970
box -8 -3 16 105
use FILL  FILL_735
timestamp 1713453518
transform 1 0 1000 0 1 2970
box -8 -3 16 105
use FILL  FILL_736
timestamp 1713453518
transform 1 0 992 0 1 2970
box -8 -3 16 105
use FILL  FILL_737
timestamp 1713453518
transform 1 0 984 0 1 2970
box -8 -3 16 105
use FILL  FILL_738
timestamp 1713453518
transform 1 0 976 0 1 2970
box -8 -3 16 105
use FILL  FILL_739
timestamp 1713453518
transform 1 0 872 0 1 2970
box -8 -3 16 105
use FILL  FILL_740
timestamp 1713453518
transform 1 0 864 0 1 2970
box -8 -3 16 105
use FILL  FILL_741
timestamp 1713453518
transform 1 0 856 0 1 2970
box -8 -3 16 105
use FILL  FILL_742
timestamp 1713453518
transform 1 0 848 0 1 2970
box -8 -3 16 105
use FILL  FILL_743
timestamp 1713453518
transform 1 0 800 0 1 2970
box -8 -3 16 105
use FILL  FILL_744
timestamp 1713453518
transform 1 0 792 0 1 2970
box -8 -3 16 105
use FILL  FILL_745
timestamp 1713453518
transform 1 0 744 0 1 2970
box -8 -3 16 105
use FILL  FILL_746
timestamp 1713453518
transform 1 0 736 0 1 2970
box -8 -3 16 105
use FILL  FILL_747
timestamp 1713453518
transform 1 0 728 0 1 2970
box -8 -3 16 105
use FILL  FILL_748
timestamp 1713453518
transform 1 0 720 0 1 2970
box -8 -3 16 105
use FILL  FILL_749
timestamp 1713453518
transform 1 0 712 0 1 2970
box -8 -3 16 105
use FILL  FILL_750
timestamp 1713453518
transform 1 0 704 0 1 2970
box -8 -3 16 105
use FILL  FILL_751
timestamp 1713453518
transform 1 0 632 0 1 2970
box -8 -3 16 105
use FILL  FILL_752
timestamp 1713453518
transform 1 0 624 0 1 2970
box -8 -3 16 105
use FILL  FILL_753
timestamp 1713453518
transform 1 0 616 0 1 2970
box -8 -3 16 105
use FILL  FILL_754
timestamp 1713453518
transform 1 0 608 0 1 2970
box -8 -3 16 105
use FILL  FILL_755
timestamp 1713453518
transform 1 0 568 0 1 2970
box -8 -3 16 105
use FILL  FILL_756
timestamp 1713453518
transform 1 0 560 0 1 2970
box -8 -3 16 105
use FILL  FILL_757
timestamp 1713453518
transform 1 0 512 0 1 2970
box -8 -3 16 105
use FILL  FILL_758
timestamp 1713453518
transform 1 0 504 0 1 2970
box -8 -3 16 105
use FILL  FILL_759
timestamp 1713453518
transform 1 0 496 0 1 2970
box -8 -3 16 105
use FILL  FILL_760
timestamp 1713453518
transform 1 0 488 0 1 2970
box -8 -3 16 105
use FILL  FILL_761
timestamp 1713453518
transform 1 0 440 0 1 2970
box -8 -3 16 105
use FILL  FILL_762
timestamp 1713453518
transform 1 0 432 0 1 2970
box -8 -3 16 105
use FILL  FILL_763
timestamp 1713453518
transform 1 0 424 0 1 2970
box -8 -3 16 105
use FILL  FILL_764
timestamp 1713453518
transform 1 0 416 0 1 2970
box -8 -3 16 105
use FILL  FILL_765
timestamp 1713453518
transform 1 0 408 0 1 2970
box -8 -3 16 105
use FILL  FILL_766
timestamp 1713453518
transform 1 0 400 0 1 2970
box -8 -3 16 105
use FILL  FILL_767
timestamp 1713453518
transform 1 0 392 0 1 2970
box -8 -3 16 105
use FILL  FILL_768
timestamp 1713453518
transform 1 0 288 0 1 2970
box -8 -3 16 105
use FILL  FILL_769
timestamp 1713453518
transform 1 0 280 0 1 2970
box -8 -3 16 105
use FILL  FILL_770
timestamp 1713453518
transform 1 0 272 0 1 2970
box -8 -3 16 105
use FILL  FILL_771
timestamp 1713453518
transform 1 0 264 0 1 2970
box -8 -3 16 105
use FILL  FILL_772
timestamp 1713453518
transform 1 0 256 0 1 2970
box -8 -3 16 105
use FILL  FILL_773
timestamp 1713453518
transform 1 0 248 0 1 2970
box -8 -3 16 105
use FILL  FILL_774
timestamp 1713453518
transform 1 0 184 0 1 2970
box -8 -3 16 105
use FILL  FILL_775
timestamp 1713453518
transform 1 0 176 0 1 2970
box -8 -3 16 105
use FILL  FILL_776
timestamp 1713453518
transform 1 0 168 0 1 2970
box -8 -3 16 105
use FILL  FILL_777
timestamp 1713453518
transform 1 0 160 0 1 2970
box -8 -3 16 105
use FILL  FILL_778
timestamp 1713453518
transform 1 0 152 0 1 2970
box -8 -3 16 105
use FILL  FILL_779
timestamp 1713453518
transform 1 0 128 0 1 2970
box -8 -3 16 105
use FILL  FILL_780
timestamp 1713453518
transform 1 0 120 0 1 2970
box -8 -3 16 105
use FILL  FILL_781
timestamp 1713453518
transform 1 0 112 0 1 2970
box -8 -3 16 105
use FILL  FILL_782
timestamp 1713453518
transform 1 0 104 0 1 2970
box -8 -3 16 105
use FILL  FILL_783
timestamp 1713453518
transform 1 0 96 0 1 2970
box -8 -3 16 105
use FILL  FILL_784
timestamp 1713453518
transform 1 0 88 0 1 2970
box -8 -3 16 105
use FILL  FILL_785
timestamp 1713453518
transform 1 0 80 0 1 2970
box -8 -3 16 105
use FILL  FILL_786
timestamp 1713453518
transform 1 0 72 0 1 2970
box -8 -3 16 105
use FILL  FILL_787
timestamp 1713453518
transform 1 0 3440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_788
timestamp 1713453518
transform 1 0 3432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_789
timestamp 1713453518
transform 1 0 3408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_790
timestamp 1713453518
transform 1 0 3400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_791
timestamp 1713453518
transform 1 0 3352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_792
timestamp 1713453518
transform 1 0 3344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_793
timestamp 1713453518
transform 1 0 3272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_794
timestamp 1713453518
transform 1 0 3264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_795
timestamp 1713453518
transform 1 0 3256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_796
timestamp 1713453518
transform 1 0 3248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_797
timestamp 1713453518
transform 1 0 3240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_798
timestamp 1713453518
transform 1 0 3176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_799
timestamp 1713453518
transform 1 0 3168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_800
timestamp 1713453518
transform 1 0 3160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_801
timestamp 1713453518
transform 1 0 3152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_802
timestamp 1713453518
transform 1 0 3144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_803
timestamp 1713453518
transform 1 0 3104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_804
timestamp 1713453518
transform 1 0 3064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_805
timestamp 1713453518
transform 1 0 3024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_806
timestamp 1713453518
transform 1 0 3016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_807
timestamp 1713453518
transform 1 0 2992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_808
timestamp 1713453518
transform 1 0 2984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_809
timestamp 1713453518
transform 1 0 2936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_810
timestamp 1713453518
transform 1 0 2928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_811
timestamp 1713453518
transform 1 0 2896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_812
timestamp 1713453518
transform 1 0 2888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_813
timestamp 1713453518
transform 1 0 2880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_814
timestamp 1713453518
transform 1 0 2872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_815
timestamp 1713453518
transform 1 0 2808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_816
timestamp 1713453518
transform 1 0 2800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_817
timestamp 1713453518
transform 1 0 2792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_818
timestamp 1713453518
transform 1 0 2784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_819
timestamp 1713453518
transform 1 0 2744 0 -1 2970
box -8 -3 16 105
use FILL  FILL_820
timestamp 1713453518
transform 1 0 2736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_821
timestamp 1713453518
transform 1 0 2728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_822
timestamp 1713453518
transform 1 0 2720 0 -1 2970
box -8 -3 16 105
use FILL  FILL_823
timestamp 1713453518
transform 1 0 2680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_824
timestamp 1713453518
transform 1 0 2672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_825
timestamp 1713453518
transform 1 0 2664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_826
timestamp 1713453518
transform 1 0 2656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_827
timestamp 1713453518
transform 1 0 2648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_828
timestamp 1713453518
transform 1 0 2600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_829
timestamp 1713453518
transform 1 0 2592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_830
timestamp 1713453518
transform 1 0 2584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_831
timestamp 1713453518
transform 1 0 2576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_832
timestamp 1713453518
transform 1 0 2568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_833
timestamp 1713453518
transform 1 0 2528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_834
timestamp 1713453518
transform 1 0 2520 0 -1 2970
box -8 -3 16 105
use FILL  FILL_835
timestamp 1713453518
transform 1 0 2512 0 -1 2970
box -8 -3 16 105
use FILL  FILL_836
timestamp 1713453518
transform 1 0 2504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_837
timestamp 1713453518
transform 1 0 2496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_838
timestamp 1713453518
transform 1 0 2464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_839
timestamp 1713453518
transform 1 0 2456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_840
timestamp 1713453518
transform 1 0 2448 0 -1 2970
box -8 -3 16 105
use FILL  FILL_841
timestamp 1713453518
transform 1 0 2440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_842
timestamp 1713453518
transform 1 0 2400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_843
timestamp 1713453518
transform 1 0 2392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_844
timestamp 1713453518
transform 1 0 2384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_845
timestamp 1713453518
transform 1 0 2376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_846
timestamp 1713453518
transform 1 0 2368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_847
timestamp 1713453518
transform 1 0 2360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_848
timestamp 1713453518
transform 1 0 2352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_849
timestamp 1713453518
transform 1 0 2304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_850
timestamp 1713453518
transform 1 0 2296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_851
timestamp 1713453518
transform 1 0 2288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_852
timestamp 1713453518
transform 1 0 2280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_853
timestamp 1713453518
transform 1 0 2272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_854
timestamp 1713453518
transform 1 0 2264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_855
timestamp 1713453518
transform 1 0 2256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_856
timestamp 1713453518
transform 1 0 2248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_857
timestamp 1713453518
transform 1 0 2200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_858
timestamp 1713453518
transform 1 0 2192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_859
timestamp 1713453518
transform 1 0 2184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_860
timestamp 1713453518
transform 1 0 2176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_861
timestamp 1713453518
transform 1 0 2168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_862
timestamp 1713453518
transform 1 0 2160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_863
timestamp 1713453518
transform 1 0 2152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_864
timestamp 1713453518
transform 1 0 2144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_865
timestamp 1713453518
transform 1 0 2096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_866
timestamp 1713453518
transform 1 0 2088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_867
timestamp 1713453518
transform 1 0 2080 0 -1 2970
box -8 -3 16 105
use FILL  FILL_868
timestamp 1713453518
transform 1 0 2072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_869
timestamp 1713453518
transform 1 0 2064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_870
timestamp 1713453518
transform 1 0 2056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_871
timestamp 1713453518
transform 1 0 2048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_872
timestamp 1713453518
transform 1 0 2000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_873
timestamp 1713453518
transform 1 0 1992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_874
timestamp 1713453518
transform 1 0 1984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_875
timestamp 1713453518
transform 1 0 1976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_876
timestamp 1713453518
transform 1 0 1968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_877
timestamp 1713453518
transform 1 0 1960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_878
timestamp 1713453518
transform 1 0 1952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_879
timestamp 1713453518
transform 1 0 1944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_880
timestamp 1713453518
transform 1 0 1896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_881
timestamp 1713453518
transform 1 0 1888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_882
timestamp 1713453518
transform 1 0 1880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_883
timestamp 1713453518
transform 1 0 1872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_884
timestamp 1713453518
transform 1 0 1864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_885
timestamp 1713453518
transform 1 0 1856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_886
timestamp 1713453518
transform 1 0 1848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_887
timestamp 1713453518
transform 1 0 1808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_888
timestamp 1713453518
transform 1 0 1800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_889
timestamp 1713453518
transform 1 0 1792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_890
timestamp 1713453518
transform 1 0 1784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_891
timestamp 1713453518
transform 1 0 1776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_892
timestamp 1713453518
transform 1 0 1768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_893
timestamp 1713453518
transform 1 0 1760 0 -1 2970
box -8 -3 16 105
use FILL  FILL_894
timestamp 1713453518
transform 1 0 1752 0 -1 2970
box -8 -3 16 105
use FILL  FILL_895
timestamp 1713453518
transform 1 0 1704 0 -1 2970
box -8 -3 16 105
use FILL  FILL_896
timestamp 1713453518
transform 1 0 1696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_897
timestamp 1713453518
transform 1 0 1688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_898
timestamp 1713453518
transform 1 0 1680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_899
timestamp 1713453518
transform 1 0 1672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_900
timestamp 1713453518
transform 1 0 1664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_901
timestamp 1713453518
transform 1 0 1656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_902
timestamp 1713453518
transform 1 0 1648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_903
timestamp 1713453518
transform 1 0 1600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_904
timestamp 1713453518
transform 1 0 1592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_905
timestamp 1713453518
transform 1 0 1584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_906
timestamp 1713453518
transform 1 0 1576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_907
timestamp 1713453518
transform 1 0 1568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_908
timestamp 1713453518
transform 1 0 1560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_909
timestamp 1713453518
transform 1 0 1552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_910
timestamp 1713453518
transform 1 0 1544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_911
timestamp 1713453518
transform 1 0 1496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_912
timestamp 1713453518
transform 1 0 1488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_913
timestamp 1713453518
transform 1 0 1480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_914
timestamp 1713453518
transform 1 0 1472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_915
timestamp 1713453518
transform 1 0 1464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_916
timestamp 1713453518
transform 1 0 1456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_917
timestamp 1713453518
transform 1 0 1416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_918
timestamp 1713453518
transform 1 0 1408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_919
timestamp 1713453518
transform 1 0 1400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_920
timestamp 1713453518
transform 1 0 1336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_921
timestamp 1713453518
transform 1 0 1328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_922
timestamp 1713453518
transform 1 0 1320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_923
timestamp 1713453518
transform 1 0 1312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_924
timestamp 1713453518
transform 1 0 1240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_925
timestamp 1713453518
transform 1 0 1232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_926
timestamp 1713453518
transform 1 0 1224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_927
timestamp 1713453518
transform 1 0 1216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_928
timestamp 1713453518
transform 1 0 1208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_929
timestamp 1713453518
transform 1 0 1168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_930
timestamp 1713453518
transform 1 0 1128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_931
timestamp 1713453518
transform 1 0 1120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_932
timestamp 1713453518
transform 1 0 1112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_933
timestamp 1713453518
transform 1 0 1104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_934
timestamp 1713453518
transform 1 0 1032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_935
timestamp 1713453518
transform 1 0 928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_936
timestamp 1713453518
transform 1 0 920 0 -1 2970
box -8 -3 16 105
use FILL  FILL_937
timestamp 1713453518
transform 1 0 784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_938
timestamp 1713453518
transform 1 0 776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_939
timestamp 1713453518
transform 1 0 768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_940
timestamp 1713453518
transform 1 0 760 0 -1 2970
box -8 -3 16 105
use FILL  FILL_941
timestamp 1713453518
transform 1 0 696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_942
timestamp 1713453518
transform 1 0 656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_943
timestamp 1713453518
transform 1 0 648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_944
timestamp 1713453518
transform 1 0 608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_945
timestamp 1713453518
transform 1 0 600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_946
timestamp 1713453518
transform 1 0 592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_947
timestamp 1713453518
transform 1 0 520 0 -1 2970
box -8 -3 16 105
use FILL  FILL_948
timestamp 1713453518
transform 1 0 512 0 -1 2970
box -8 -3 16 105
use FILL  FILL_949
timestamp 1713453518
transform 1 0 504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_950
timestamp 1713453518
transform 1 0 496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_951
timestamp 1713453518
transform 1 0 392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_952
timestamp 1713453518
transform 1 0 384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_953
timestamp 1713453518
transform 1 0 376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_954
timestamp 1713453518
transform 1 0 272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_955
timestamp 1713453518
transform 1 0 264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_956
timestamp 1713453518
transform 1 0 184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_957
timestamp 1713453518
transform 1 0 176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_958
timestamp 1713453518
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_959
timestamp 1713453518
transform 1 0 3384 0 1 2770
box -8 -3 16 105
use FILL  FILL_960
timestamp 1713453518
transform 1 0 3336 0 1 2770
box -8 -3 16 105
use FILL  FILL_961
timestamp 1713453518
transform 1 0 3280 0 1 2770
box -8 -3 16 105
use FILL  FILL_962
timestamp 1713453518
transform 1 0 3256 0 1 2770
box -8 -3 16 105
use FILL  FILL_963
timestamp 1713453518
transform 1 0 3224 0 1 2770
box -8 -3 16 105
use FILL  FILL_964
timestamp 1713453518
transform 1 0 3216 0 1 2770
box -8 -3 16 105
use FILL  FILL_965
timestamp 1713453518
transform 1 0 3144 0 1 2770
box -8 -3 16 105
use FILL  FILL_966
timestamp 1713453518
transform 1 0 3136 0 1 2770
box -8 -3 16 105
use FILL  FILL_967
timestamp 1713453518
transform 1 0 3128 0 1 2770
box -8 -3 16 105
use FILL  FILL_968
timestamp 1713453518
transform 1 0 3056 0 1 2770
box -8 -3 16 105
use FILL  FILL_969
timestamp 1713453518
transform 1 0 3048 0 1 2770
box -8 -3 16 105
use FILL  FILL_970
timestamp 1713453518
transform 1 0 3040 0 1 2770
box -8 -3 16 105
use FILL  FILL_971
timestamp 1713453518
transform 1 0 2976 0 1 2770
box -8 -3 16 105
use FILL  FILL_972
timestamp 1713453518
transform 1 0 2896 0 1 2770
box -8 -3 16 105
use FILL  FILL_973
timestamp 1713453518
transform 1 0 2888 0 1 2770
box -8 -3 16 105
use FILL  FILL_974
timestamp 1713453518
transform 1 0 2880 0 1 2770
box -8 -3 16 105
use FILL  FILL_975
timestamp 1713453518
transform 1 0 2800 0 1 2770
box -8 -3 16 105
use FILL  FILL_976
timestamp 1713453518
transform 1 0 2792 0 1 2770
box -8 -3 16 105
use FILL  FILL_977
timestamp 1713453518
transform 1 0 2736 0 1 2770
box -8 -3 16 105
use FILL  FILL_978
timestamp 1713453518
transform 1 0 2728 0 1 2770
box -8 -3 16 105
use FILL  FILL_979
timestamp 1713453518
transform 1 0 2696 0 1 2770
box -8 -3 16 105
use FILL  FILL_980
timestamp 1713453518
transform 1 0 2688 0 1 2770
box -8 -3 16 105
use FILL  FILL_981
timestamp 1713453518
transform 1 0 2664 0 1 2770
box -8 -3 16 105
use FILL  FILL_982
timestamp 1713453518
transform 1 0 2632 0 1 2770
box -8 -3 16 105
use FILL  FILL_983
timestamp 1713453518
transform 1 0 2624 0 1 2770
box -8 -3 16 105
use FILL  FILL_984
timestamp 1713453518
transform 1 0 2616 0 1 2770
box -8 -3 16 105
use FILL  FILL_985
timestamp 1713453518
transform 1 0 2608 0 1 2770
box -8 -3 16 105
use FILL  FILL_986
timestamp 1713453518
transform 1 0 2600 0 1 2770
box -8 -3 16 105
use FILL  FILL_987
timestamp 1713453518
transform 1 0 2592 0 1 2770
box -8 -3 16 105
use FILL  FILL_988
timestamp 1713453518
transform 1 0 2560 0 1 2770
box -8 -3 16 105
use FILL  FILL_989
timestamp 1713453518
transform 1 0 2552 0 1 2770
box -8 -3 16 105
use FILL  FILL_990
timestamp 1713453518
transform 1 0 2544 0 1 2770
box -8 -3 16 105
use FILL  FILL_991
timestamp 1713453518
transform 1 0 2496 0 1 2770
box -8 -3 16 105
use FILL  FILL_992
timestamp 1713453518
transform 1 0 2488 0 1 2770
box -8 -3 16 105
use FILL  FILL_993
timestamp 1713453518
transform 1 0 2480 0 1 2770
box -8 -3 16 105
use FILL  FILL_994
timestamp 1713453518
transform 1 0 2472 0 1 2770
box -8 -3 16 105
use FILL  FILL_995
timestamp 1713453518
transform 1 0 2464 0 1 2770
box -8 -3 16 105
use FILL  FILL_996
timestamp 1713453518
transform 1 0 2456 0 1 2770
box -8 -3 16 105
use FILL  FILL_997
timestamp 1713453518
transform 1 0 2448 0 1 2770
box -8 -3 16 105
use FILL  FILL_998
timestamp 1713453518
transform 1 0 2408 0 1 2770
box -8 -3 16 105
use FILL  FILL_999
timestamp 1713453518
transform 1 0 2400 0 1 2770
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1713453518
transform 1 0 2392 0 1 2770
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1713453518
transform 1 0 2384 0 1 2770
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1713453518
transform 1 0 2376 0 1 2770
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1713453518
transform 1 0 2368 0 1 2770
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1713453518
transform 1 0 2328 0 1 2770
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1713453518
transform 1 0 2320 0 1 2770
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1713453518
transform 1 0 2312 0 1 2770
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1713453518
transform 1 0 2304 0 1 2770
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1713453518
transform 1 0 2296 0 1 2770
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1713453518
transform 1 0 2288 0 1 2770
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1713453518
transform 1 0 2280 0 1 2770
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1713453518
transform 1 0 2272 0 1 2770
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1713453518
transform 1 0 2224 0 1 2770
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1713453518
transform 1 0 2216 0 1 2770
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1713453518
transform 1 0 2208 0 1 2770
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1713453518
transform 1 0 2200 0 1 2770
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1713453518
transform 1 0 2192 0 1 2770
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1713453518
transform 1 0 2184 0 1 2770
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1713453518
transform 1 0 2176 0 1 2770
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1713453518
transform 1 0 2168 0 1 2770
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1713453518
transform 1 0 2160 0 1 2770
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1713453518
transform 1 0 2112 0 1 2770
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1713453518
transform 1 0 2104 0 1 2770
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1713453518
transform 1 0 2096 0 1 2770
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1713453518
transform 1 0 2088 0 1 2770
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1713453518
transform 1 0 2080 0 1 2770
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1713453518
transform 1 0 2072 0 1 2770
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1713453518
transform 1 0 2064 0 1 2770
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1713453518
transform 1 0 2040 0 1 2770
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1713453518
transform 1 0 2032 0 1 2770
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1713453518
transform 1 0 2024 0 1 2770
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1713453518
transform 1 0 2016 0 1 2770
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1713453518
transform 1 0 1984 0 1 2770
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1713453518
transform 1 0 1976 0 1 2770
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1713453518
transform 1 0 1968 0 1 2770
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1713453518
transform 1 0 1960 0 1 2770
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1713453518
transform 1 0 1952 0 1 2770
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1713453518
transform 1 0 1944 0 1 2770
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1713453518
transform 1 0 1912 0 1 2770
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1713453518
transform 1 0 1904 0 1 2770
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1713453518
transform 1 0 1896 0 1 2770
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1713453518
transform 1 0 1888 0 1 2770
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1713453518
transform 1 0 1880 0 1 2770
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1713453518
transform 1 0 1872 0 1 2770
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1713453518
transform 1 0 1864 0 1 2770
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1713453518
transform 1 0 1832 0 1 2770
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1713453518
transform 1 0 1824 0 1 2770
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1713453518
transform 1 0 1816 0 1 2770
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1713453518
transform 1 0 1808 0 1 2770
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1713453518
transform 1 0 1784 0 1 2770
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1713453518
transform 1 0 1776 0 1 2770
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1713453518
transform 1 0 1768 0 1 2770
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1713453518
transform 1 0 1760 0 1 2770
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1713453518
transform 1 0 1752 0 1 2770
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1713453518
transform 1 0 1720 0 1 2770
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1713453518
transform 1 0 1712 0 1 2770
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1713453518
transform 1 0 1704 0 1 2770
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1713453518
transform 1 0 1696 0 1 2770
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1713453518
transform 1 0 1688 0 1 2770
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1713453518
transform 1 0 1680 0 1 2770
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1713453518
transform 1 0 1648 0 1 2770
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1713453518
transform 1 0 1640 0 1 2770
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1713453518
transform 1 0 1632 0 1 2770
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1713453518
transform 1 0 1624 0 1 2770
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1713453518
transform 1 0 1616 0 1 2770
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1713453518
transform 1 0 1608 0 1 2770
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1713453518
transform 1 0 1600 0 1 2770
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1713453518
transform 1 0 1568 0 1 2770
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1713453518
transform 1 0 1560 0 1 2770
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1713453518
transform 1 0 1552 0 1 2770
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1713453518
transform 1 0 1544 0 1 2770
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1713453518
transform 1 0 1504 0 1 2770
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1713453518
transform 1 0 1496 0 1 2770
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1713453518
transform 1 0 1488 0 1 2770
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1713453518
transform 1 0 1480 0 1 2770
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1713453518
transform 1 0 1440 0 1 2770
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1713453518
transform 1 0 1432 0 1 2770
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1713453518
transform 1 0 1424 0 1 2770
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1713453518
transform 1 0 1392 0 1 2770
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1713453518
transform 1 0 1384 0 1 2770
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1713453518
transform 1 0 1360 0 1 2770
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1713453518
transform 1 0 1352 0 1 2770
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1713453518
transform 1 0 1344 0 1 2770
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1713453518
transform 1 0 1304 0 1 2770
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1713453518
transform 1 0 1296 0 1 2770
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1713453518
transform 1 0 1288 0 1 2770
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1713453518
transform 1 0 1248 0 1 2770
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1713453518
transform 1 0 1240 0 1 2770
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1713453518
transform 1 0 1232 0 1 2770
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1713453518
transform 1 0 1224 0 1 2770
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1713453518
transform 1 0 1216 0 1 2770
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1713453518
transform 1 0 1160 0 1 2770
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1713453518
transform 1 0 1152 0 1 2770
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1713453518
transform 1 0 1144 0 1 2770
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1713453518
transform 1 0 1136 0 1 2770
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1713453518
transform 1 0 1128 0 1 2770
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1713453518
transform 1 0 1096 0 1 2770
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1713453518
transform 1 0 1088 0 1 2770
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1713453518
transform 1 0 1064 0 1 2770
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1713453518
transform 1 0 1056 0 1 2770
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1713453518
transform 1 0 1016 0 1 2770
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1713453518
transform 1 0 1008 0 1 2770
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1713453518
transform 1 0 1000 0 1 2770
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1713453518
transform 1 0 992 0 1 2770
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1713453518
transform 1 0 984 0 1 2770
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1713453518
transform 1 0 976 0 1 2770
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1713453518
transform 1 0 968 0 1 2770
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1713453518
transform 1 0 960 0 1 2770
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1713453518
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1713453518
transform 1 0 888 0 1 2770
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1713453518
transform 1 0 880 0 1 2770
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1713453518
transform 1 0 872 0 1 2770
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1713453518
transform 1 0 864 0 1 2770
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1713453518
transform 1 0 824 0 1 2770
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1713453518
transform 1 0 816 0 1 2770
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1713453518
transform 1 0 808 0 1 2770
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1713453518
transform 1 0 736 0 1 2770
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1713453518
transform 1 0 728 0 1 2770
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1713453518
transform 1 0 720 0 1 2770
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1713453518
transform 1 0 712 0 1 2770
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1713453518
transform 1 0 664 0 1 2770
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1713453518
transform 1 0 616 0 1 2770
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1713453518
transform 1 0 608 0 1 2770
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1713453518
transform 1 0 600 0 1 2770
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1713453518
transform 1 0 592 0 1 2770
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1713453518
transform 1 0 544 0 1 2770
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1713453518
transform 1 0 536 0 1 2770
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1713453518
transform 1 0 488 0 1 2770
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1713453518
transform 1 0 480 0 1 2770
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1713453518
transform 1 0 432 0 1 2770
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1713453518
transform 1 0 424 0 1 2770
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1713453518
transform 1 0 416 0 1 2770
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1713453518
transform 1 0 408 0 1 2770
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1713453518
transform 1 0 304 0 1 2770
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1713453518
transform 1 0 296 0 1 2770
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1713453518
transform 1 0 288 0 1 2770
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1713453518
transform 1 0 280 0 1 2770
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1713453518
transform 1 0 200 0 1 2770
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1713453518
transform 1 0 192 0 1 2770
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1713453518
transform 1 0 184 0 1 2770
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1713453518
transform 1 0 176 0 1 2770
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1713453518
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1713453518
transform 1 0 3440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1713453518
transform 1 0 3392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1713453518
transform 1 0 3320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1713453518
transform 1 0 3312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1713453518
transform 1 0 3304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1713453518
transform 1 0 3248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1713453518
transform 1 0 3240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1713453518
transform 1 0 3232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1713453518
transform 1 0 3192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1713453518
transform 1 0 3184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1713453518
transform 1 0 3144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1713453518
transform 1 0 3136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1713453518
transform 1 0 3088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1713453518
transform 1 0 3080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1713453518
transform 1 0 3072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1713453518
transform 1 0 3016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1713453518
transform 1 0 2984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1713453518
transform 1 0 2976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1713453518
transform 1 0 2968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1713453518
transform 1 0 2888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1713453518
transform 1 0 2880 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1713453518
transform 1 0 2872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1713453518
transform 1 0 2824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1713453518
transform 1 0 2752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1713453518
transform 1 0 2744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1713453518
transform 1 0 2736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1713453518
transform 1 0 2696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1713453518
transform 1 0 2688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1713453518
transform 1 0 2640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1713453518
transform 1 0 2632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1713453518
transform 1 0 2600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1713453518
transform 1 0 2592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1713453518
transform 1 0 2584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1713453518
transform 1 0 2576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1713453518
transform 1 0 2568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1713453518
transform 1 0 2520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1713453518
transform 1 0 2512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1713453518
transform 1 0 2504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1713453518
transform 1 0 2496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1713453518
transform 1 0 2488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1713453518
transform 1 0 2480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1713453518
transform 1 0 2472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1713453518
transform 1 0 2464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1713453518
transform 1 0 2416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1713453518
transform 1 0 2408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1713453518
transform 1 0 2400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1713453518
transform 1 0 2392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1713453518
transform 1 0 2384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1713453518
transform 1 0 2376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1713453518
transform 1 0 2368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1713453518
transform 1 0 2360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1713453518
transform 1 0 2312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1713453518
transform 1 0 2304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1713453518
transform 1 0 2296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1713453518
transform 1 0 2288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1713453518
transform 1 0 2280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1713453518
transform 1 0 2272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1713453518
transform 1 0 2264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1713453518
transform 1 0 2232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1713453518
transform 1 0 2224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1713453518
transform 1 0 2200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1713453518
transform 1 0 2192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1713453518
transform 1 0 2184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1713453518
transform 1 0 2176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1713453518
transform 1 0 2128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1713453518
transform 1 0 2120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1713453518
transform 1 0 2112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1713453518
transform 1 0 2104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1713453518
transform 1 0 2096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1713453518
transform 1 0 2064 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1713453518
transform 1 0 2056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1713453518
transform 1 0 2048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1713453518
transform 1 0 2040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1713453518
transform 1 0 2032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1713453518
transform 1 0 2024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1713453518
transform 1 0 2016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1713453518
transform 1 0 1968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1713453518
transform 1 0 1960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1713453518
transform 1 0 1952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1713453518
transform 1 0 1944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1713453518
transform 1 0 1936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1713453518
transform 1 0 1928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1713453518
transform 1 0 1920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1713453518
transform 1 0 1880 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1713453518
transform 1 0 1872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1713453518
transform 1 0 1864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1713453518
transform 1 0 1856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1713453518
transform 1 0 1848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1713453518
transform 1 0 1840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1713453518
transform 1 0 1800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1713453518
transform 1 0 1792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1713453518
transform 1 0 1784 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1713453518
transform 1 0 1776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1713453518
transform 1 0 1768 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1713453518
transform 1 0 1760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1713453518
transform 1 0 1752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1713453518
transform 1 0 1704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1713453518
transform 1 0 1696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1713453518
transform 1 0 1688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1713453518
transform 1 0 1680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1713453518
transform 1 0 1672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1713453518
transform 1 0 1664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1713453518
transform 1 0 1656 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1713453518
transform 1 0 1648 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1713453518
transform 1 0 1616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1713453518
transform 1 0 1608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1713453518
transform 1 0 1576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1713453518
transform 1 0 1568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1713453518
transform 1 0 1560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1713453518
transform 1 0 1552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1713453518
transform 1 0 1520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1713453518
transform 1 0 1512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1713453518
transform 1 0 1504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1713453518
transform 1 0 1472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1713453518
transform 1 0 1464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1713453518
transform 1 0 1456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1713453518
transform 1 0 1408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1713453518
transform 1 0 1400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1713453518
transform 1 0 1392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1713453518
transform 1 0 1384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1713453518
transform 1 0 1336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1713453518
transform 1 0 1328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1713453518
transform 1 0 1304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1713453518
transform 1 0 1296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1713453518
transform 1 0 1288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1713453518
transform 1 0 1280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1713453518
transform 1 0 1232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1713453518
transform 1 0 1224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1713453518
transform 1 0 1192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1713453518
transform 1 0 1184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1713453518
transform 1 0 1176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1713453518
transform 1 0 1144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1713453518
transform 1 0 1136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1713453518
transform 1 0 1128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1713453518
transform 1 0 1120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1713453518
transform 1 0 1056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1713453518
transform 1 0 1048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1713453518
transform 1 0 1040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1713453518
transform 1 0 936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1713453518
transform 1 0 928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1713453518
transform 1 0 920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1713453518
transform 1 0 912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1713453518
transform 1 0 904 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1713453518
transform 1 0 840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1713453518
transform 1 0 832 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1713453518
transform 1 0 792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1713453518
transform 1 0 784 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1713453518
transform 1 0 776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1713453518
transform 1 0 728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1713453518
transform 1 0 720 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1713453518
transform 1 0 712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1713453518
transform 1 0 664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1713453518
transform 1 0 656 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1713453518
transform 1 0 648 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1713453518
transform 1 0 640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1713453518
transform 1 0 576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1713453518
transform 1 0 568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1713453518
transform 1 0 560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1713453518
transform 1 0 552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1713453518
transform 1 0 480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1713453518
transform 1 0 472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1713453518
transform 1 0 464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1713453518
transform 1 0 456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1713453518
transform 1 0 352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1713453518
transform 1 0 344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1713453518
transform 1 0 336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1713453518
transform 1 0 328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1713453518
transform 1 0 320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1713453518
transform 1 0 240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1713453518
transform 1 0 232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1713453518
transform 1 0 224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1713453518
transform 1 0 216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1713453518
transform 1 0 208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1713453518
transform 1 0 200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1713453518
transform 1 0 96 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1713453518
transform 1 0 88 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1713453518
transform 1 0 80 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1713453518
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1713453518
transform 1 0 3440 0 1 2570
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1713453518
transform 1 0 3432 0 1 2570
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1713453518
transform 1 0 3384 0 1 2570
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1713453518
transform 1 0 3376 0 1 2570
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1713453518
transform 1 0 3368 0 1 2570
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1713453518
transform 1 0 3312 0 1 2570
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1713453518
transform 1 0 3304 0 1 2570
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1713453518
transform 1 0 3256 0 1 2570
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1713453518
transform 1 0 3248 0 1 2570
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1713453518
transform 1 0 3240 0 1 2570
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1713453518
transform 1 0 3232 0 1 2570
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1713453518
transform 1 0 3200 0 1 2570
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1713453518
transform 1 0 3168 0 1 2570
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1713453518
transform 1 0 3160 0 1 2570
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1713453518
transform 1 0 3152 0 1 2570
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1713453518
transform 1 0 3144 0 1 2570
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1713453518
transform 1 0 3136 0 1 2570
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1713453518
transform 1 0 3128 0 1 2570
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1713453518
transform 1 0 3064 0 1 2570
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1713453518
transform 1 0 3056 0 1 2570
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1713453518
transform 1 0 3048 0 1 2570
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1713453518
transform 1 0 3040 0 1 2570
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1713453518
transform 1 0 2992 0 1 2570
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1713453518
transform 1 0 2984 0 1 2570
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1713453518
transform 1 0 2976 0 1 2570
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1713453518
transform 1 0 2968 0 1 2570
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1713453518
transform 1 0 2904 0 1 2570
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1713453518
transform 1 0 2896 0 1 2570
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1713453518
transform 1 0 2888 0 1 2570
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1713453518
transform 1 0 2880 0 1 2570
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1713453518
transform 1 0 2848 0 1 2570
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1713453518
transform 1 0 2808 0 1 2570
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1713453518
transform 1 0 2800 0 1 2570
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1713453518
transform 1 0 2760 0 1 2570
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1713453518
transform 1 0 2752 0 1 2570
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1713453518
transform 1 0 2744 0 1 2570
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1713453518
transform 1 0 2736 0 1 2570
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1713453518
transform 1 0 2728 0 1 2570
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1713453518
transform 1 0 2696 0 1 2570
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1713453518
transform 1 0 2640 0 1 2570
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1713453518
transform 1 0 2632 0 1 2570
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1713453518
transform 1 0 2624 0 1 2570
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1713453518
transform 1 0 2616 0 1 2570
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1713453518
transform 1 0 2608 0 1 2570
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1713453518
transform 1 0 2600 0 1 2570
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1713453518
transform 1 0 2560 0 1 2570
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1713453518
transform 1 0 2552 0 1 2570
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1713453518
transform 1 0 2544 0 1 2570
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1713453518
transform 1 0 2536 0 1 2570
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1713453518
transform 1 0 2504 0 1 2570
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1713453518
transform 1 0 2496 0 1 2570
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1713453518
transform 1 0 2488 0 1 2570
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1713453518
transform 1 0 2480 0 1 2570
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1713453518
transform 1 0 2432 0 1 2570
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1713453518
transform 1 0 2424 0 1 2570
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1713453518
transform 1 0 2416 0 1 2570
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1713453518
transform 1 0 2408 0 1 2570
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1713453518
transform 1 0 2400 0 1 2570
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1713453518
transform 1 0 2392 0 1 2570
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1713453518
transform 1 0 2384 0 1 2570
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1713453518
transform 1 0 2336 0 1 2570
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1713453518
transform 1 0 2328 0 1 2570
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1713453518
transform 1 0 2320 0 1 2570
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1713453518
transform 1 0 2296 0 1 2570
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1713453518
transform 1 0 2288 0 1 2570
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1713453518
transform 1 0 2280 0 1 2570
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1713453518
transform 1 0 2272 0 1 2570
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1713453518
transform 1 0 2240 0 1 2570
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1713453518
transform 1 0 2232 0 1 2570
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1713453518
transform 1 0 2224 0 1 2570
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1713453518
transform 1 0 2184 0 1 2570
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1713453518
transform 1 0 2176 0 1 2570
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1713453518
transform 1 0 2168 0 1 2570
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1713453518
transform 1 0 2160 0 1 2570
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1713453518
transform 1 0 2152 0 1 2570
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1713453518
transform 1 0 2144 0 1 2570
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1713453518
transform 1 0 2104 0 1 2570
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1713453518
transform 1 0 2096 0 1 2570
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1713453518
transform 1 0 2088 0 1 2570
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1713453518
transform 1 0 2080 0 1 2570
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1713453518
transform 1 0 2048 0 1 2570
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1713453518
transform 1 0 2040 0 1 2570
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1713453518
transform 1 0 2032 0 1 2570
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1713453518
transform 1 0 2024 0 1 2570
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1713453518
transform 1 0 1984 0 1 2570
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1713453518
transform 1 0 1976 0 1 2570
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1713453518
transform 1 0 1968 0 1 2570
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1713453518
transform 1 0 1960 0 1 2570
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1713453518
transform 1 0 1952 0 1 2570
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1713453518
transform 1 0 1944 0 1 2570
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1713453518
transform 1 0 1896 0 1 2570
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1713453518
transform 1 0 1888 0 1 2570
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1713453518
transform 1 0 1880 0 1 2570
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1713453518
transform 1 0 1872 0 1 2570
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1713453518
transform 1 0 1864 0 1 2570
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1713453518
transform 1 0 1856 0 1 2570
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1713453518
transform 1 0 1824 0 1 2570
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1713453518
transform 1 0 1816 0 1 2570
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1713453518
transform 1 0 1808 0 1 2570
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1713453518
transform 1 0 1784 0 1 2570
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1713453518
transform 1 0 1776 0 1 2570
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1713453518
transform 1 0 1768 0 1 2570
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1713453518
transform 1 0 1760 0 1 2570
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1713453518
transform 1 0 1752 0 1 2570
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1713453518
transform 1 0 1744 0 1 2570
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1713453518
transform 1 0 1712 0 1 2570
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1713453518
transform 1 0 1704 0 1 2570
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1713453518
transform 1 0 1696 0 1 2570
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1713453518
transform 1 0 1688 0 1 2570
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1713453518
transform 1 0 1648 0 1 2570
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1713453518
transform 1 0 1640 0 1 2570
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1713453518
transform 1 0 1632 0 1 2570
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1713453518
transform 1 0 1624 0 1 2570
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1713453518
transform 1 0 1616 0 1 2570
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1713453518
transform 1 0 1576 0 1 2570
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1713453518
transform 1 0 1568 0 1 2570
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1713453518
transform 1 0 1560 0 1 2570
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1713453518
transform 1 0 1552 0 1 2570
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1713453518
transform 1 0 1544 0 1 2570
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1713453518
transform 1 0 1512 0 1 2570
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1713453518
transform 1 0 1504 0 1 2570
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1713453518
transform 1 0 1496 0 1 2570
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1713453518
transform 1 0 1456 0 1 2570
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1713453518
transform 1 0 1448 0 1 2570
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1713453518
transform 1 0 1440 0 1 2570
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1713453518
transform 1 0 1432 0 1 2570
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1713453518
transform 1 0 1400 0 1 2570
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1713453518
transform 1 0 1392 0 1 2570
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1713453518
transform 1 0 1384 0 1 2570
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1713453518
transform 1 0 1344 0 1 2570
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1713453518
transform 1 0 1336 0 1 2570
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1713453518
transform 1 0 1328 0 1 2570
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1713453518
transform 1 0 1320 0 1 2570
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1713453518
transform 1 0 1280 0 1 2570
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1713453518
transform 1 0 1272 0 1 2570
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1713453518
transform 1 0 1232 0 1 2570
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1713453518
transform 1 0 1224 0 1 2570
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1713453518
transform 1 0 1216 0 1 2570
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1713453518
transform 1 0 1208 0 1 2570
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1713453518
transform 1 0 1160 0 1 2570
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1713453518
transform 1 0 1152 0 1 2570
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1713453518
transform 1 0 1144 0 1 2570
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1713453518
transform 1 0 1112 0 1 2570
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1713453518
transform 1 0 1104 0 1 2570
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1713453518
transform 1 0 1096 0 1 2570
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1713453518
transform 1 0 1088 0 1 2570
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1713453518
transform 1 0 1016 0 1 2570
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1713453518
transform 1 0 1008 0 1 2570
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1713453518
transform 1 0 1000 0 1 2570
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1713453518
transform 1 0 896 0 1 2570
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1713453518
transform 1 0 888 0 1 2570
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1713453518
transform 1 0 880 0 1 2570
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1713453518
transform 1 0 816 0 1 2570
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1713453518
transform 1 0 808 0 1 2570
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1713453518
transform 1 0 728 0 1 2570
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1713453518
transform 1 0 720 0 1 2570
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1713453518
transform 1 0 624 0 1 2570
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1713453518
transform 1 0 616 0 1 2570
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1713453518
transform 1 0 608 0 1 2570
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1713453518
transform 1 0 600 0 1 2570
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1713453518
transform 1 0 528 0 1 2570
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1713453518
transform 1 0 520 0 1 2570
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1713453518
transform 1 0 472 0 1 2570
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1713453518
transform 1 0 464 0 1 2570
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1713453518
transform 1 0 360 0 1 2570
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1713453518
transform 1 0 352 0 1 2570
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1713453518
transform 1 0 344 0 1 2570
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1713453518
transform 1 0 336 0 1 2570
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1713453518
transform 1 0 328 0 1 2570
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1713453518
transform 1 0 264 0 1 2570
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1713453518
transform 1 0 208 0 1 2570
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1713453518
transform 1 0 200 0 1 2570
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1713453518
transform 1 0 192 0 1 2570
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1713453518
transform 1 0 184 0 1 2570
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1713453518
transform 1 0 80 0 1 2570
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1713453518
transform 1 0 72 0 1 2570
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1713453518
transform 1 0 3440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1713453518
transform 1 0 3376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1713453518
transform 1 0 3368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1713453518
transform 1 0 3360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1713453518
transform 1 0 3264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1713453518
transform 1 0 3256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1713453518
transform 1 0 3248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1713453518
transform 1 0 3240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1713453518
transform 1 0 3184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1713453518
transform 1 0 3176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1713453518
transform 1 0 3168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1713453518
transform 1 0 3160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1713453518
transform 1 0 3152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1713453518
transform 1 0 3144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1713453518
transform 1 0 3088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1713453518
transform 1 0 3080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1713453518
transform 1 0 3072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1713453518
transform 1 0 3048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1713453518
transform 1 0 3040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1713453518
transform 1 0 3032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1713453518
transform 1 0 3024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1713453518
transform 1 0 2960 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1713453518
transform 1 0 2952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1713453518
transform 1 0 2944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1713453518
transform 1 0 2896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1713453518
transform 1 0 2888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1713453518
transform 1 0 2856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1713453518
transform 1 0 2848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1713453518
transform 1 0 2840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1713453518
transform 1 0 2800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1713453518
transform 1 0 2792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1713453518
transform 1 0 2784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1713453518
transform 1 0 2736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1713453518
transform 1 0 2728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1713453518
transform 1 0 2720 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1713453518
transform 1 0 2712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1713453518
transform 1 0 2672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1713453518
transform 1 0 2664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1713453518
transform 1 0 2632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1713453518
transform 1 0 2624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1713453518
transform 1 0 2616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1713453518
transform 1 0 2608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1713453518
transform 1 0 2600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1713453518
transform 1 0 2552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1713453518
transform 1 0 2544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1713453518
transform 1 0 2536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1713453518
transform 1 0 2528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1713453518
transform 1 0 2520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1713453518
transform 1 0 2512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1713453518
transform 1 0 2504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1713453518
transform 1 0 2496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1713453518
transform 1 0 2456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1713453518
transform 1 0 2448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1713453518
transform 1 0 2440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1713453518
transform 1 0 2432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1713453518
transform 1 0 2392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1713453518
transform 1 0 2384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1713453518
transform 1 0 2376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1713453518
transform 1 0 2368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1713453518
transform 1 0 2360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1713453518
transform 1 0 2352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1713453518
transform 1 0 2344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1713453518
transform 1 0 2336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1713453518
transform 1 0 2288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1713453518
transform 1 0 2280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1713453518
transform 1 0 2272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1713453518
transform 1 0 2264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1713453518
transform 1 0 2256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1713453518
transform 1 0 2248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1713453518
transform 1 0 2240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1713453518
transform 1 0 2192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1713453518
transform 1 0 2184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1713453518
transform 1 0 2176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1713453518
transform 1 0 2168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1713453518
transform 1 0 2160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1713453518
transform 1 0 2120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1713453518
transform 1 0 2112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1713453518
transform 1 0 2104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1713453518
transform 1 0 2072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1713453518
transform 1 0 2064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1713453518
transform 1 0 2056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1713453518
transform 1 0 2048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1713453518
transform 1 0 2040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1713453518
transform 1 0 2032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1713453518
transform 1 0 2024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1713453518
transform 1 0 1976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1713453518
transform 1 0 1968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1713453518
transform 1 0 1960 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1713453518
transform 1 0 1952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1713453518
transform 1 0 1944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1713453518
transform 1 0 1920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1713453518
transform 1 0 1912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1713453518
transform 1 0 1904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1713453518
transform 1 0 1872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1713453518
transform 1 0 1864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1713453518
transform 1 0 1856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1713453518
transform 1 0 1848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1713453518
transform 1 0 1808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1713453518
transform 1 0 1800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1713453518
transform 1 0 1792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1713453518
transform 1 0 1784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1713453518
transform 1 0 1744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1713453518
transform 1 0 1736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1713453518
transform 1 0 1728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1713453518
transform 1 0 1696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1713453518
transform 1 0 1688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1713453518
transform 1 0 1680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1713453518
transform 1 0 1672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1713453518
transform 1 0 1664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1713453518
transform 1 0 1624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1713453518
transform 1 0 1616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1713453518
transform 1 0 1608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1713453518
transform 1 0 1600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1713453518
transform 1 0 1560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1713453518
transform 1 0 1552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1713453518
transform 1 0 1544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1713453518
transform 1 0 1536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1713453518
transform 1 0 1528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1713453518
transform 1 0 1472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1713453518
transform 1 0 1464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1713453518
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1713453518
transform 1 0 1448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1713453518
transform 1 0 1440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1713453518
transform 1 0 1392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1713453518
transform 1 0 1368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1713453518
transform 1 0 1360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1713453518
transform 1 0 1336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1713453518
transform 1 0 1328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1713453518
transform 1 0 1320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1713453518
transform 1 0 1312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1713453518
transform 1 0 1272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1713453518
transform 1 0 1232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1713453518
transform 1 0 1224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1713453518
transform 1 0 1216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1713453518
transform 1 0 1208 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1713453518
transform 1 0 1200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1713453518
transform 1 0 1152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1713453518
transform 1 0 1144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1713453518
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1713453518
transform 1 0 1104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1713453518
transform 1 0 1096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1713453518
transform 1 0 1088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1713453518
transform 1 0 1080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1713453518
transform 1 0 1008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1713453518
transform 1 0 1000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1713453518
transform 1 0 992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1713453518
transform 1 0 984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1713453518
transform 1 0 880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1713453518
transform 1 0 872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1713453518
transform 1 0 864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1713453518
transform 1 0 856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1713453518
transform 1 0 848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1713453518
transform 1 0 784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1713453518
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1713453518
transform 1 0 744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1713453518
transform 1 0 736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1713453518
transform 1 0 728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1713453518
transform 1 0 688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1713453518
transform 1 0 640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1713453518
transform 1 0 632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1713453518
transform 1 0 624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1713453518
transform 1 0 616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1713453518
transform 1 0 608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1713453518
transform 1 0 552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1713453518
transform 1 0 512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1713453518
transform 1 0 504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1713453518
transform 1 0 496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1713453518
transform 1 0 488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1713453518
transform 1 0 416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1713453518
transform 1 0 408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1713453518
transform 1 0 304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1713453518
transform 1 0 296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1713453518
transform 1 0 288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1713453518
transform 1 0 280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1713453518
transform 1 0 272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1713453518
transform 1 0 192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1713453518
transform 1 0 184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1713453518
transform 1 0 176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1713453518
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1713453518
transform 1 0 3440 0 1 2370
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1713453518
transform 1 0 3432 0 1 2370
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1713453518
transform 1 0 3424 0 1 2370
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1713453518
transform 1 0 3384 0 1 2370
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1713453518
transform 1 0 3360 0 1 2370
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1713453518
transform 1 0 3336 0 1 2370
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1713453518
transform 1 0 3328 0 1 2370
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1713453518
transform 1 0 3320 0 1 2370
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1713453518
transform 1 0 3288 0 1 2370
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1713453518
transform 1 0 3280 0 1 2370
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1713453518
transform 1 0 3272 0 1 2370
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1713453518
transform 1 0 3240 0 1 2370
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1713453518
transform 1 0 3232 0 1 2370
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1713453518
transform 1 0 3224 0 1 2370
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1713453518
transform 1 0 3192 0 1 2370
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1713453518
transform 1 0 3184 0 1 2370
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1713453518
transform 1 0 3176 0 1 2370
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1713453518
transform 1 0 3168 0 1 2370
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1713453518
transform 1 0 3120 0 1 2370
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1713453518
transform 1 0 3112 0 1 2370
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1713453518
transform 1 0 3104 0 1 2370
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1713453518
transform 1 0 3096 0 1 2370
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1713453518
transform 1 0 3088 0 1 2370
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1713453518
transform 1 0 3080 0 1 2370
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1713453518
transform 1 0 3048 0 1 2370
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1713453518
transform 1 0 3040 0 1 2370
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1713453518
transform 1 0 3032 0 1 2370
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1713453518
transform 1 0 2984 0 1 2370
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1713453518
transform 1 0 2976 0 1 2370
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1713453518
transform 1 0 2968 0 1 2370
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1713453518
transform 1 0 2960 0 1 2370
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1713453518
transform 1 0 2952 0 1 2370
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1713453518
transform 1 0 2904 0 1 2370
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1713453518
transform 1 0 2896 0 1 2370
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1713453518
transform 1 0 2864 0 1 2370
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1713453518
transform 1 0 2856 0 1 2370
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1713453518
transform 1 0 2848 0 1 2370
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1713453518
transform 1 0 2840 0 1 2370
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1713453518
transform 1 0 2832 0 1 2370
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1713453518
transform 1 0 2824 0 1 2370
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1713453518
transform 1 0 2816 0 1 2370
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1713453518
transform 1 0 2752 0 1 2370
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1713453518
transform 1 0 2744 0 1 2370
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1713453518
transform 1 0 2736 0 1 2370
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1713453518
transform 1 0 2728 0 1 2370
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1713453518
transform 1 0 2720 0 1 2370
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1713453518
transform 1 0 2712 0 1 2370
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1713453518
transform 1 0 2704 0 1 2370
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1713453518
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1713453518
transform 1 0 2632 0 1 2370
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1713453518
transform 1 0 2624 0 1 2370
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1713453518
transform 1 0 2616 0 1 2370
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1713453518
transform 1 0 2608 0 1 2370
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1713453518
transform 1 0 2600 0 1 2370
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1713453518
transform 1 0 2560 0 1 2370
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1713453518
transform 1 0 2552 0 1 2370
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1713453518
transform 1 0 2544 0 1 2370
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1713453518
transform 1 0 2536 0 1 2370
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1713453518
transform 1 0 2496 0 1 2370
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1713453518
transform 1 0 2488 0 1 2370
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1713453518
transform 1 0 2480 0 1 2370
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1713453518
transform 1 0 2472 0 1 2370
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1713453518
transform 1 0 2464 0 1 2370
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1713453518
transform 1 0 2456 0 1 2370
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1713453518
transform 1 0 2448 0 1 2370
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1713453518
transform 1 0 2440 0 1 2370
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1713453518
transform 1 0 2392 0 1 2370
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1713453518
transform 1 0 2384 0 1 2370
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1713453518
transform 1 0 2376 0 1 2370
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1713453518
transform 1 0 2368 0 1 2370
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1713453518
transform 1 0 2360 0 1 2370
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1713453518
transform 1 0 2352 0 1 2370
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1713453518
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1713453518
transform 1 0 2336 0 1 2370
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1713453518
transform 1 0 2328 0 1 2370
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1713453518
transform 1 0 2280 0 1 2370
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1713453518
transform 1 0 2272 0 1 2370
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1713453518
transform 1 0 2264 0 1 2370
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1713453518
transform 1 0 2256 0 1 2370
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1713453518
transform 1 0 2248 0 1 2370
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1713453518
transform 1 0 2240 0 1 2370
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1713453518
transform 1 0 2216 0 1 2370
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1713453518
transform 1 0 2208 0 1 2370
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1713453518
transform 1 0 2200 0 1 2370
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1713453518
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1713453518
transform 1 0 2152 0 1 2370
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1713453518
transform 1 0 2144 0 1 2370
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1713453518
transform 1 0 2136 0 1 2370
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1713453518
transform 1 0 2128 0 1 2370
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1713453518
transform 1 0 2120 0 1 2370
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1713453518
transform 1 0 2112 0 1 2370
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1713453518
transform 1 0 2064 0 1 2370
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1713453518
transform 1 0 2056 0 1 2370
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1713453518
transform 1 0 2048 0 1 2370
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1713453518
transform 1 0 2040 0 1 2370
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1713453518
transform 1 0 2032 0 1 2370
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1713453518
transform 1 0 2008 0 1 2370
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1713453518
transform 1 0 2000 0 1 2370
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1713453518
transform 1 0 1992 0 1 2370
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1713453518
transform 1 0 1984 0 1 2370
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1713453518
transform 1 0 1936 0 1 2370
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1713453518
transform 1 0 1928 0 1 2370
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1713453518
transform 1 0 1920 0 1 2370
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1713453518
transform 1 0 1912 0 1 2370
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1713453518
transform 1 0 1904 0 1 2370
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1713453518
transform 1 0 1896 0 1 2370
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1713453518
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1713453518
transform 1 0 1856 0 1 2370
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1713453518
transform 1 0 1848 0 1 2370
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1713453518
transform 1 0 1816 0 1 2370
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1713453518
transform 1 0 1808 0 1 2370
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1713453518
transform 1 0 1800 0 1 2370
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1713453518
transform 1 0 1792 0 1 2370
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1713453518
transform 1 0 1784 0 1 2370
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1713453518
transform 1 0 1776 0 1 2370
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1713453518
transform 1 0 1736 0 1 2370
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1713453518
transform 1 0 1728 0 1 2370
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1713453518
transform 1 0 1720 0 1 2370
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1713453518
transform 1 0 1688 0 1 2370
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1713453518
transform 1 0 1680 0 1 2370
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1713453518
transform 1 0 1672 0 1 2370
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1713453518
transform 1 0 1664 0 1 2370
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1713453518
transform 1 0 1656 0 1 2370
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1713453518
transform 1 0 1608 0 1 2370
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1713453518
transform 1 0 1600 0 1 2370
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1713453518
transform 1 0 1592 0 1 2370
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1713453518
transform 1 0 1584 0 1 2370
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1713453518
transform 1 0 1552 0 1 2370
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1713453518
transform 1 0 1544 0 1 2370
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1713453518
transform 1 0 1536 0 1 2370
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1713453518
transform 1 0 1496 0 1 2370
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1713453518
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1713453518
transform 1 0 1480 0 1 2370
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1713453518
transform 1 0 1472 0 1 2370
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1713453518
transform 1 0 1424 0 1 2370
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1713453518
transform 1 0 1416 0 1 2370
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1713453518
transform 1 0 1408 0 1 2370
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1713453518
transform 1 0 1400 0 1 2370
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1713453518
transform 1 0 1392 0 1 2370
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1713453518
transform 1 0 1352 0 1 2370
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1713453518
transform 1 0 1344 0 1 2370
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1713453518
transform 1 0 1336 0 1 2370
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1713453518
transform 1 0 1288 0 1 2370
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1713453518
transform 1 0 1280 0 1 2370
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1713453518
transform 1 0 1272 0 1 2370
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1713453518
transform 1 0 1264 0 1 2370
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1713453518
transform 1 0 1256 0 1 2370
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1713453518
transform 1 0 1248 0 1 2370
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1713453518
transform 1 0 1208 0 1 2370
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1713453518
transform 1 0 1200 0 1 2370
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1713453518
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1713453518
transform 1 0 1152 0 1 2370
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1713453518
transform 1 0 1144 0 1 2370
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1713453518
transform 1 0 1136 0 1 2370
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1713453518
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1713453518
transform 1 0 1056 0 1 2370
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1713453518
transform 1 0 1048 0 1 2370
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1713453518
transform 1 0 1040 0 1 2370
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1713453518
transform 1 0 1032 0 1 2370
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1713453518
transform 1 0 928 0 1 2370
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1713453518
transform 1 0 920 0 1 2370
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1713453518
transform 1 0 912 0 1 2370
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1713453518
transform 1 0 904 0 1 2370
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1713453518
transform 1 0 896 0 1 2370
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1713453518
transform 1 0 888 0 1 2370
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1713453518
transform 1 0 880 0 1 2370
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1713453518
transform 1 0 816 0 1 2370
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1713453518
transform 1 0 808 0 1 2370
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1713453518
transform 1 0 800 0 1 2370
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1713453518
transform 1 0 792 0 1 2370
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1713453518
transform 1 0 744 0 1 2370
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1713453518
transform 1 0 704 0 1 2370
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1713453518
transform 1 0 696 0 1 2370
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1713453518
transform 1 0 688 0 1 2370
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1713453518
transform 1 0 680 0 1 2370
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1713453518
transform 1 0 672 0 1 2370
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1713453518
transform 1 0 632 0 1 2370
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1713453518
transform 1 0 624 0 1 2370
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1713453518
transform 1 0 616 0 1 2370
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1713453518
transform 1 0 560 0 1 2370
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1713453518
transform 1 0 552 0 1 2370
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1713453518
transform 1 0 544 0 1 2370
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1713453518
transform 1 0 536 0 1 2370
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1713453518
transform 1 0 488 0 1 2370
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1713453518
transform 1 0 456 0 1 2370
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1713453518
transform 1 0 448 0 1 2370
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1713453518
transform 1 0 440 0 1 2370
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1713453518
transform 1 0 432 0 1 2370
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1713453518
transform 1 0 384 0 1 2370
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1713453518
transform 1 0 376 0 1 2370
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1713453518
transform 1 0 368 0 1 2370
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1713453518
transform 1 0 360 0 1 2370
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1713453518
transform 1 0 352 0 1 2370
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1713453518
transform 1 0 344 0 1 2370
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1713453518
transform 1 0 240 0 1 2370
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1713453518
transform 1 0 232 0 1 2370
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1713453518
transform 1 0 224 0 1 2370
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1713453518
transform 1 0 216 0 1 2370
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1713453518
transform 1 0 208 0 1 2370
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1713453518
transform 1 0 176 0 1 2370
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1713453518
transform 1 0 168 0 1 2370
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1713453518
transform 1 0 160 0 1 2370
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1713453518
transform 1 0 152 0 1 2370
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1713453518
transform 1 0 144 0 1 2370
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1713453518
transform 1 0 136 0 1 2370
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1713453518
transform 1 0 128 0 1 2370
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1713453518
transform 1 0 120 0 1 2370
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1713453518
transform 1 0 112 0 1 2370
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1713453518
transform 1 0 104 0 1 2370
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1713453518
transform 1 0 96 0 1 2370
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1713453518
transform 1 0 88 0 1 2370
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1713453518
transform 1 0 80 0 1 2370
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1713453518
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1713453518
transform 1 0 3440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1713453518
transform 1 0 3432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1713453518
transform 1 0 3384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1713453518
transform 1 0 3376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1713453518
transform 1 0 3368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1713453518
transform 1 0 3360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1713453518
transform 1 0 3352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1713453518
transform 1 0 3344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1713453518
transform 1 0 3288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1713453518
transform 1 0 3280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1713453518
transform 1 0 3272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1713453518
transform 1 0 3248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1713453518
transform 1 0 3240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1713453518
transform 1 0 3232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1713453518
transform 1 0 3224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1713453518
transform 1 0 3192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1713453518
transform 1 0 3184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1713453518
transform 1 0 3176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1713453518
transform 1 0 3136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1713453518
transform 1 0 3128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1713453518
transform 1 0 3120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1713453518
transform 1 0 3112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1713453518
transform 1 0 3104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1713453518
transform 1 0 3096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1713453518
transform 1 0 3048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1713453518
transform 1 0 3040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1713453518
transform 1 0 3032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1713453518
transform 1 0 3024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1713453518
transform 1 0 2992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1713453518
transform 1 0 2984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1713453518
transform 1 0 2976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1713453518
transform 1 0 2968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1713453518
transform 1 0 2928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1713453518
transform 1 0 2920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1713453518
transform 1 0 2912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1713453518
transform 1 0 2904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1713453518
transform 1 0 2864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1713453518
transform 1 0 2856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1713453518
transform 1 0 2848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1713453518
transform 1 0 2840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1713453518
transform 1 0 2808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1713453518
transform 1 0 2800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1713453518
transform 1 0 2792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1713453518
transform 1 0 2784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1713453518
transform 1 0 2744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1713453518
transform 1 0 2736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1713453518
transform 1 0 2728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1713453518
transform 1 0 2720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1713453518
transform 1 0 2672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1713453518
transform 1 0 2664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1713453518
transform 1 0 2656 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1713453518
transform 1 0 2648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1713453518
transform 1 0 2640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1713453518
transform 1 0 2592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1713453518
transform 1 0 2584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1713453518
transform 1 0 2576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1713453518
transform 1 0 2568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1713453518
transform 1 0 2544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1713453518
transform 1 0 2536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1713453518
transform 1 0 2496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1713453518
transform 1 0 2488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1713453518
transform 1 0 2480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1713453518
transform 1 0 2472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1713453518
transform 1 0 2464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1713453518
transform 1 0 2432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1713453518
transform 1 0 2424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1713453518
transform 1 0 2416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1713453518
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1713453518
transform 1 0 2376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1713453518
transform 1 0 2368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1713453518
transform 1 0 2360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1713453518
transform 1 0 2352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1713453518
transform 1 0 2344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1713453518
transform 1 0 2336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1713453518
transform 1 0 2288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1713453518
transform 1 0 2280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1713453518
transform 1 0 2272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1713453518
transform 1 0 2264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1713453518
transform 1 0 2256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1713453518
transform 1 0 2248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1713453518
transform 1 0 2240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1713453518
transform 1 0 2232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1713453518
transform 1 0 2192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1713453518
transform 1 0 2184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1713453518
transform 1 0 2176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1713453518
transform 1 0 2168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1713453518
transform 1 0 2160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1713453518
transform 1 0 2128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1713453518
transform 1 0 2120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1713453518
transform 1 0 2112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1713453518
transform 1 0 2104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1713453518
transform 1 0 2096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1713453518
transform 1 0 2056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1713453518
transform 1 0 2048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1713453518
transform 1 0 2040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1713453518
transform 1 0 2032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1713453518
transform 1 0 2024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1713453518
transform 1 0 2016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1713453518
transform 1 0 1984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1713453518
transform 1 0 1976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1713453518
transform 1 0 1968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1713453518
transform 1 0 1960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1713453518
transform 1 0 1952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1713453518
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1713453518
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1713453518
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1713453518
transform 1 0 1888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1713453518
transform 1 0 1880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1713453518
transform 1 0 1856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1713453518
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1713453518
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1713453518
transform 1 0 1832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1713453518
transform 1 0 1824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1713453518
transform 1 0 1816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1713453518
transform 1 0 1776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1713453518
transform 1 0 1768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1713453518
transform 1 0 1760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1713453518
transform 1 0 1752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1713453518
transform 1 0 1744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1713453518
transform 1 0 1736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1713453518
transform 1 0 1728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1713453518
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1713453518
transform 1 0 1680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1713453518
transform 1 0 1672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1713453518
transform 1 0 1664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1713453518
transform 1 0 1656 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1713453518
transform 1 0 1648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1713453518
transform 1 0 1640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1713453518
transform 1 0 1592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1713453518
transform 1 0 1584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1713453518
transform 1 0 1576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1713453518
transform 1 0 1544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1713453518
transform 1 0 1536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1713453518
transform 1 0 1528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1713453518
transform 1 0 1520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1713453518
transform 1 0 1512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1713453518
transform 1 0 1464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1713453518
transform 1 0 1456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1713453518
transform 1 0 1448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1713453518
transform 1 0 1440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1713453518
transform 1 0 1416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1713453518
transform 1 0 1408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1713453518
transform 1 0 1376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1713453518
transform 1 0 1344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1713453518
transform 1 0 1336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1713453518
transform 1 0 1328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1713453518
transform 1 0 1320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1713453518
transform 1 0 1312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1713453518
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1713453518
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1713453518
transform 1 0 1224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1713453518
transform 1 0 1216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1713453518
transform 1 0 1208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1713453518
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1713453518
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1713453518
transform 1 0 1136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1713453518
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1713453518
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1713453518
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1713453518
transform 1 0 1104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1713453518
transform 1 0 1032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1713453518
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1713453518
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1713453518
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1713453518
transform 1 0 904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1713453518
transform 1 0 896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1713453518
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1713453518
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1713453518
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1713453518
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1713453518
transform 1 0 728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1713453518
transform 1 0 720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1713453518
transform 1 0 712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1713453518
transform 1 0 704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1713453518
transform 1 0 624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1713453518
transform 1 0 616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1713453518
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1713453518
transform 1 0 464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1713453518
transform 1 0 456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1713453518
transform 1 0 448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1713453518
transform 1 0 368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1713453518
transform 1 0 360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1713453518
transform 1 0 352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1713453518
transform 1 0 248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1713453518
transform 1 0 240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1713453518
transform 1 0 232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1713453518
transform 1 0 176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1713453518
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1713453518
transform 1 0 3440 0 1 2170
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1713453518
transform 1 0 3432 0 1 2170
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1713453518
transform 1 0 3424 0 1 2170
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1713453518
transform 1 0 3416 0 1 2170
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1713453518
transform 1 0 3352 0 1 2170
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1713453518
transform 1 0 3344 0 1 2170
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1713453518
transform 1 0 3336 0 1 2170
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1713453518
transform 1 0 3328 0 1 2170
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1713453518
transform 1 0 3264 0 1 2170
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1713453518
transform 1 0 3256 0 1 2170
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1713453518
transform 1 0 3248 0 1 2170
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1713453518
transform 1 0 3240 0 1 2170
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1713453518
transform 1 0 3232 0 1 2170
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1713453518
transform 1 0 3224 0 1 2170
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1713453518
transform 1 0 3184 0 1 2170
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1713453518
transform 1 0 3176 0 1 2170
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1713453518
transform 1 0 3168 0 1 2170
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1713453518
transform 1 0 3160 0 1 2170
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1713453518
transform 1 0 3120 0 1 2170
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1713453518
transform 1 0 3112 0 1 2170
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1713453518
transform 1 0 3104 0 1 2170
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1713453518
transform 1 0 3096 0 1 2170
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1713453518
transform 1 0 3088 0 1 2170
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1713453518
transform 1 0 3048 0 1 2170
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1713453518
transform 1 0 3040 0 1 2170
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1713453518
transform 1 0 3032 0 1 2170
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1713453518
transform 1 0 2992 0 1 2170
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1713453518
transform 1 0 2984 0 1 2170
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1713453518
transform 1 0 2976 0 1 2170
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1713453518
transform 1 0 2968 0 1 2170
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1713453518
transform 1 0 2928 0 1 2170
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1713453518
transform 1 0 2920 0 1 2170
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1713453518
transform 1 0 2912 0 1 2170
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1713453518
transform 1 0 2904 0 1 2170
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1713453518
transform 1 0 2856 0 1 2170
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1713453518
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1713453518
transform 1 0 2840 0 1 2170
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1713453518
transform 1 0 2832 0 1 2170
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1713453518
transform 1 0 2824 0 1 2170
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1713453518
transform 1 0 2800 0 1 2170
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1713453518
transform 1 0 2792 0 1 2170
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1713453518
transform 1 0 2752 0 1 2170
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1713453518
transform 1 0 2744 0 1 2170
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1713453518
transform 1 0 2736 0 1 2170
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1713453518
transform 1 0 2728 0 1 2170
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1713453518
transform 1 0 2720 0 1 2170
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1713453518
transform 1 0 2712 0 1 2170
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1713453518
transform 1 0 2680 0 1 2170
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1713453518
transform 1 0 2672 0 1 2170
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1713453518
transform 1 0 2664 0 1 2170
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1713453518
transform 1 0 2624 0 1 2170
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1713453518
transform 1 0 2616 0 1 2170
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1713453518
transform 1 0 2608 0 1 2170
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1713453518
transform 1 0 2600 0 1 2170
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1713453518
transform 1 0 2592 0 1 2170
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1713453518
transform 1 0 2584 0 1 2170
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1713453518
transform 1 0 2576 0 1 2170
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1713453518
transform 1 0 2528 0 1 2170
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1713453518
transform 1 0 2520 0 1 2170
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1713453518
transform 1 0 2512 0 1 2170
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1713453518
transform 1 0 2504 0 1 2170
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1713453518
transform 1 0 2496 0 1 2170
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1713453518
transform 1 0 2488 0 1 2170
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1713453518
transform 1 0 2480 0 1 2170
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1713453518
transform 1 0 2432 0 1 2170
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1713453518
transform 1 0 2424 0 1 2170
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1713453518
transform 1 0 2416 0 1 2170
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1713453518
transform 1 0 2408 0 1 2170
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1713453518
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1713453518
transform 1 0 2360 0 1 2170
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1713453518
transform 1 0 2352 0 1 2170
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1713453518
transform 1 0 2344 0 1 2170
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1713453518
transform 1 0 2336 0 1 2170
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1713453518
transform 1 0 2288 0 1 2170
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1713453518
transform 1 0 2280 0 1 2170
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1713453518
transform 1 0 2272 0 1 2170
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1713453518
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1713453518
transform 1 0 2256 0 1 2170
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1713453518
transform 1 0 2216 0 1 2170
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1713453518
transform 1 0 2208 0 1 2170
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1713453518
transform 1 0 2200 0 1 2170
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1713453518
transform 1 0 2192 0 1 2170
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1713453518
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1713453518
transform 1 0 2176 0 1 2170
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1713453518
transform 1 0 2168 0 1 2170
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1713453518
transform 1 0 2120 0 1 2170
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1713453518
transform 1 0 2112 0 1 2170
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1713453518
transform 1 0 2104 0 1 2170
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1713453518
transform 1 0 2096 0 1 2170
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1713453518
transform 1 0 2088 0 1 2170
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1713453518
transform 1 0 2080 0 1 2170
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1713453518
transform 1 0 2072 0 1 2170
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1713453518
transform 1 0 2064 0 1 2170
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1713453518
transform 1 0 2016 0 1 2170
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1713453518
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1713453518
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1713453518
transform 1 0 1992 0 1 2170
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1713453518
transform 1 0 1984 0 1 2170
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1713453518
transform 1 0 1976 0 1 2170
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1713453518
transform 1 0 1968 0 1 2170
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1713453518
transform 1 0 1960 0 1 2170
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1713453518
transform 1 0 1912 0 1 2170
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1713453518
transform 1 0 1904 0 1 2170
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1713453518
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1713453518
transform 1 0 1888 0 1 2170
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1713453518
transform 1 0 1880 0 1 2170
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1713453518
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1713453518
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1713453518
transform 1 0 1832 0 1 2170
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1713453518
transform 1 0 1824 0 1 2170
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1713453518
transform 1 0 1816 0 1 2170
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1713453518
transform 1 0 1776 0 1 2170
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1713453518
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1713453518
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1713453518
transform 1 0 1752 0 1 2170
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1713453518
transform 1 0 1744 0 1 2170
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1713453518
transform 1 0 1704 0 1 2170
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1713453518
transform 1 0 1696 0 1 2170
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1713453518
transform 1 0 1688 0 1 2170
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1713453518
transform 1 0 1680 0 1 2170
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1713453518
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1713453518
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1713453518
transform 1 0 1624 0 1 2170
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1713453518
transform 1 0 1616 0 1 2170
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1713453518
transform 1 0 1608 0 1 2170
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1713453518
transform 1 0 1600 0 1 2170
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1713453518
transform 1 0 1592 0 1 2170
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1713453518
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1713453518
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1713453518
transform 1 0 1520 0 1 2170
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1713453518
transform 1 0 1512 0 1 2170
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1713453518
transform 1 0 1504 0 1 2170
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1713453518
transform 1 0 1496 0 1 2170
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1713453518
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1713453518
transform 1 0 1424 0 1 2170
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1713453518
transform 1 0 1416 0 1 2170
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1713453518
transform 1 0 1408 0 1 2170
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1713453518
transform 1 0 1400 0 1 2170
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1713453518
transform 1 0 1392 0 1 2170
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1713453518
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1713453518
transform 1 0 1344 0 1 2170
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1713453518
transform 1 0 1336 0 1 2170
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1713453518
transform 1 0 1296 0 1 2170
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1713453518
transform 1 0 1288 0 1 2170
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1713453518
transform 1 0 1280 0 1 2170
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1713453518
transform 1 0 1272 0 1 2170
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1713453518
transform 1 0 1264 0 1 2170
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1713453518
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1713453518
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1713453518
transform 1 0 1208 0 1 2170
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1713453518
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1713453518
transform 1 0 1160 0 1 2170
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1713453518
transform 1 0 1152 0 1 2170
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1713453518
transform 1 0 1144 0 1 2170
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1713453518
transform 1 0 1136 0 1 2170
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1713453518
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1713453518
transform 1 0 1072 0 1 2170
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1713453518
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1713453518
transform 1 0 1056 0 1 2170
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1713453518
transform 1 0 1048 0 1 2170
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1713453518
transform 1 0 976 0 1 2170
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1713453518
transform 1 0 968 0 1 2170
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1713453518
transform 1 0 960 0 1 2170
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1713453518
transform 1 0 952 0 1 2170
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1713453518
transform 1 0 848 0 1 2170
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1713453518
transform 1 0 840 0 1 2170
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1713453518
transform 1 0 832 0 1 2170
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1713453518
transform 1 0 824 0 1 2170
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1713453518
transform 1 0 760 0 1 2170
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1713453518
transform 1 0 752 0 1 2170
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1713453518
transform 1 0 744 0 1 2170
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1713453518
transform 1 0 680 0 1 2170
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1713453518
transform 1 0 672 0 1 2170
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1713453518
transform 1 0 664 0 1 2170
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1713453518
transform 1 0 656 0 1 2170
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1713453518
transform 1 0 648 0 1 2170
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1713453518
transform 1 0 552 0 1 2170
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1713453518
transform 1 0 544 0 1 2170
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1713453518
transform 1 0 536 0 1 2170
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1713453518
transform 1 0 528 0 1 2170
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1713453518
transform 1 0 520 0 1 2170
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1713453518
transform 1 0 432 0 1 2170
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1713453518
transform 1 0 424 0 1 2170
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1713453518
transform 1 0 416 0 1 2170
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1713453518
transform 1 0 408 0 1 2170
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1713453518
transform 1 0 304 0 1 2170
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1713453518
transform 1 0 296 0 1 2170
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1713453518
transform 1 0 288 0 1 2170
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1713453518
transform 1 0 280 0 1 2170
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1713453518
transform 1 0 200 0 1 2170
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1713453518
transform 1 0 192 0 1 2170
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1713453518
transform 1 0 184 0 1 2170
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1713453518
transform 1 0 176 0 1 2170
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1713453518
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1713453518
transform 1 0 3440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1713453518
transform 1 0 3432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1713453518
transform 1 0 3384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1713453518
transform 1 0 3376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1713453518
transform 1 0 3368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1713453518
transform 1 0 3360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1713453518
transform 1 0 3352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1713453518
transform 1 0 3296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1713453518
transform 1 0 3288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1713453518
transform 1 0 3280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1713453518
transform 1 0 3272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1713453518
transform 1 0 3264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1713453518
transform 1 0 3232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1713453518
transform 1 0 3224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1713453518
transform 1 0 3216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1713453518
transform 1 0 3176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1713453518
transform 1 0 3168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1713453518
transform 1 0 3160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1713453518
transform 1 0 3152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1713453518
transform 1 0 3144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1713453518
transform 1 0 3104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1713453518
transform 1 0 3096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1713453518
transform 1 0 3088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1713453518
transform 1 0 3056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1713453518
transform 1 0 3048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1713453518
transform 1 0 3040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1713453518
transform 1 0 3032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1713453518
transform 1 0 2984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1713453518
transform 1 0 2976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1713453518
transform 1 0 2968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1713453518
transform 1 0 2944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1713453518
transform 1 0 2936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1713453518
transform 1 0 2912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1713453518
transform 1 0 2904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1713453518
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1713453518
transform 1 0 2856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1713453518
transform 1 0 2848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1713453518
transform 1 0 2840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1713453518
transform 1 0 2800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1713453518
transform 1 0 2792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1713453518
transform 1 0 2784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1713453518
transform 1 0 2776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1713453518
transform 1 0 2768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1713453518
transform 1 0 2728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1713453518
transform 1 0 2720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1713453518
transform 1 0 2712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1713453518
transform 1 0 2680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1713453518
transform 1 0 2672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1713453518
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1713453518
transform 1 0 2640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1713453518
transform 1 0 2632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1713453518
transform 1 0 2624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1713453518
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1713453518
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1713453518
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1713453518
transform 1 0 2536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1713453518
transform 1 0 2528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1713453518
transform 1 0 2520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1713453518
transform 1 0 2512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1713453518
transform 1 0 2504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1713453518
transform 1 0 2440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1713453518
transform 1 0 2432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1713453518
transform 1 0 2424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1713453518
transform 1 0 2416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1713453518
transform 1 0 2408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1713453518
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1713453518
transform 1 0 2392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1713453518
transform 1 0 2344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1713453518
transform 1 0 2336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1713453518
transform 1 0 2328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1713453518
transform 1 0 2320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1713453518
transform 1 0 2312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1713453518
transform 1 0 2304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1713453518
transform 1 0 2264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1713453518
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1713453518
transform 1 0 2248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1713453518
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1713453518
transform 1 0 2208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1713453518
transform 1 0 2200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1713453518
transform 1 0 2192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1713453518
transform 1 0 2184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1713453518
transform 1 0 2176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1713453518
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1713453518
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1713453518
transform 1 0 2112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1713453518
transform 1 0 2104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1713453518
transform 1 0 2096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1713453518
transform 1 0 2088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1713453518
transform 1 0 2056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1713453518
transform 1 0 2048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1713453518
transform 1 0 2040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1713453518
transform 1 0 2008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1713453518
transform 1 0 2000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1713453518
transform 1 0 1992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1713453518
transform 1 0 1984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1713453518
transform 1 0 1976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1713453518
transform 1 0 1968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1713453518
transform 1 0 1928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1713453518
transform 1 0 1920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1713453518
transform 1 0 1912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1713453518
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1713453518
transform 1 0 1896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1713453518
transform 1 0 1872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1713453518
transform 1 0 1864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1713453518
transform 1 0 1832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1713453518
transform 1 0 1824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1713453518
transform 1 0 1816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1713453518
transform 1 0 1808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1713453518
transform 1 0 1800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1713453518
transform 1 0 1760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1713453518
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1713453518
transform 1 0 1744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1713453518
transform 1 0 1736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1713453518
transform 1 0 1728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1713453518
transform 1 0 1720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1713453518
transform 1 0 1712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1713453518
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1713453518
transform 1 0 1648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1713453518
transform 1 0 1640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1713453518
transform 1 0 1632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1713453518
transform 1 0 1624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1713453518
transform 1 0 1616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1713453518
transform 1 0 1592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1713453518
transform 1 0 1560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1713453518
transform 1 0 1552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1713453518
transform 1 0 1544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1713453518
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1713453518
transform 1 0 1496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1713453518
transform 1 0 1488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1713453518
transform 1 0 1464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1713453518
transform 1 0 1456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1713453518
transform 1 0 1448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1713453518
transform 1 0 1440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1713453518
transform 1 0 1432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1713453518
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1713453518
transform 1 0 1384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1713453518
transform 1 0 1352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1713453518
transform 1 0 1344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1713453518
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1713453518
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1713453518
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1713453518
transform 1 0 1288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1713453518
transform 1 0 1256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1713453518
transform 1 0 1248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1713453518
transform 1 0 1240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1713453518
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1713453518
transform 1 0 1224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1713453518
transform 1 0 1176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1713453518
transform 1 0 1168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1713453518
transform 1 0 1160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1713453518
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1713453518
transform 1 0 1120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1713453518
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1713453518
transform 1 0 1072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1713453518
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1713453518
transform 1 0 1056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1713453518
transform 1 0 992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1713453518
transform 1 0 984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1713453518
transform 1 0 976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1713453518
transform 1 0 872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1713453518
transform 1 0 864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1713453518
transform 1 0 856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1713453518
transform 1 0 848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1713453518
transform 1 0 840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1713453518
transform 1 0 776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1713453518
transform 1 0 768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1713453518
transform 1 0 760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1713453518
transform 1 0 752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1713453518
transform 1 0 680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1713453518
transform 1 0 672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1713453518
transform 1 0 664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1713453518
transform 1 0 656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1713453518
transform 1 0 648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1713453518
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1713453518
transform 1 0 560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1713453518
transform 1 0 552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1713453518
transform 1 0 544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1713453518
transform 1 0 520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1713453518
transform 1 0 512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1713453518
transform 1 0 504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1713453518
transform 1 0 432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1713453518
transform 1 0 424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1713453518
transform 1 0 416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1713453518
transform 1 0 312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1713453518
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1713453518
transform 1 0 296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1713453518
transform 1 0 288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1713453518
transform 1 0 208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1713453518
transform 1 0 200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1713453518
transform 1 0 192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1713453518
transform 1 0 184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1713453518
transform 1 0 80 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1713453518
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1713453518
transform 1 0 3440 0 1 1970
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1713453518
transform 1 0 3432 0 1 1970
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1713453518
transform 1 0 3424 0 1 1970
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1713453518
transform 1 0 3360 0 1 1970
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1713453518
transform 1 0 3352 0 1 1970
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1713453518
transform 1 0 3344 0 1 1970
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1713453518
transform 1 0 3336 0 1 1970
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1713453518
transform 1 0 3288 0 1 1970
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1713453518
transform 1 0 3280 0 1 1970
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1713453518
transform 1 0 3272 0 1 1970
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1713453518
transform 1 0 3240 0 1 1970
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1713453518
transform 1 0 3232 0 1 1970
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1713453518
transform 1 0 3224 0 1 1970
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1713453518
transform 1 0 3216 0 1 1970
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1713453518
transform 1 0 3208 0 1 1970
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1713453518
transform 1 0 3200 0 1 1970
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1713453518
transform 1 0 3160 0 1 1970
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1713453518
transform 1 0 3152 0 1 1970
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1713453518
transform 1 0 3144 0 1 1970
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1713453518
transform 1 0 3136 0 1 1970
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1713453518
transform 1 0 3128 0 1 1970
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1713453518
transform 1 0 3120 0 1 1970
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1713453518
transform 1 0 3080 0 1 1970
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1713453518
transform 1 0 3072 0 1 1970
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1713453518
transform 1 0 3064 0 1 1970
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1713453518
transform 1 0 3032 0 1 1970
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1713453518
transform 1 0 3024 0 1 1970
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1713453518
transform 1 0 3016 0 1 1970
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1713453518
transform 1 0 3008 0 1 1970
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1713453518
transform 1 0 3000 0 1 1970
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1713453518
transform 1 0 2992 0 1 1970
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1713453518
transform 1 0 2944 0 1 1970
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1713453518
transform 1 0 2936 0 1 1970
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1713453518
transform 1 0 2928 0 1 1970
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1713453518
transform 1 0 2920 0 1 1970
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1713453518
transform 1 0 2912 0 1 1970
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1713453518
transform 1 0 2904 0 1 1970
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1713453518
transform 1 0 2848 0 1 1970
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1713453518
transform 1 0 2840 0 1 1970
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1713453518
transform 1 0 2832 0 1 1970
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1713453518
transform 1 0 2824 0 1 1970
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1713453518
transform 1 0 2816 0 1 1970
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1713453518
transform 1 0 2808 0 1 1970
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1713453518
transform 1 0 2752 0 1 1970
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1713453518
transform 1 0 2744 0 1 1970
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1713453518
transform 1 0 2736 0 1 1970
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1713453518
transform 1 0 2728 0 1 1970
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1713453518
transform 1 0 2720 0 1 1970
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1713453518
transform 1 0 2688 0 1 1970
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1713453518
transform 1 0 2680 0 1 1970
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1713453518
transform 1 0 2640 0 1 1970
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1713453518
transform 1 0 2632 0 1 1970
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1713453518
transform 1 0 2624 0 1 1970
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1713453518
transform 1 0 2616 0 1 1970
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1713453518
transform 1 0 2608 0 1 1970
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1713453518
transform 1 0 2576 0 1 1970
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1713453518
transform 1 0 2568 0 1 1970
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1713453518
transform 1 0 2560 0 1 1970
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1713453518
transform 1 0 2552 0 1 1970
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1713453518
transform 1 0 2504 0 1 1970
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1713453518
transform 1 0 2496 0 1 1970
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1713453518
transform 1 0 2488 0 1 1970
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1713453518
transform 1 0 2480 0 1 1970
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1713453518
transform 1 0 2472 0 1 1970
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1713453518
transform 1 0 2432 0 1 1970
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1713453518
transform 1 0 2424 0 1 1970
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1713453518
transform 1 0 2416 0 1 1970
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1713453518
transform 1 0 2408 0 1 1970
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1713453518
transform 1 0 2400 0 1 1970
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1713453518
transform 1 0 2392 0 1 1970
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1713453518
transform 1 0 2384 0 1 1970
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1713453518
transform 1 0 2336 0 1 1970
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1713453518
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1713453518
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1713453518
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1713453518
transform 1 0 2304 0 1 1970
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1713453518
transform 1 0 2296 0 1 1970
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1713453518
transform 1 0 2288 0 1 1970
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1713453518
transform 1 0 2280 0 1 1970
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1713453518
transform 1 0 2272 0 1 1970
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1713453518
transform 1 0 2224 0 1 1970
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1713453518
transform 1 0 2216 0 1 1970
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1713453518
transform 1 0 2208 0 1 1970
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1713453518
transform 1 0 2200 0 1 1970
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1713453518
transform 1 0 2192 0 1 1970
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1713453518
transform 1 0 2184 0 1 1970
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1713453518
transform 1 0 2176 0 1 1970
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1713453518
transform 1 0 2168 0 1 1970
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1713453518
transform 1 0 2128 0 1 1970
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1713453518
transform 1 0 2120 0 1 1970
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1713453518
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1713453518
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1713453518
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1713453518
transform 1 0 2088 0 1 1970
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1713453518
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1713453518
transform 1 0 2040 0 1 1970
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1713453518
transform 1 0 2032 0 1 1970
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1713453518
transform 1 0 2024 0 1 1970
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1713453518
transform 1 0 2016 0 1 1970
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1713453518
transform 1 0 2008 0 1 1970
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1713453518
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1713453518
transform 1 0 1960 0 1 1970
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1713453518
transform 1 0 1952 0 1 1970
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1713453518
transform 1 0 1944 0 1 1970
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1713453518
transform 1 0 1936 0 1 1970
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1713453518
transform 1 0 1928 0 1 1970
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1713453518
transform 1 0 1920 0 1 1970
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1713453518
transform 1 0 1880 0 1 1970
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1713453518
transform 1 0 1872 0 1 1970
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1713453518
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1713453518
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1713453518
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1713453518
transform 1 0 1816 0 1 1970
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1713453518
transform 1 0 1808 0 1 1970
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1713453518
transform 1 0 1800 0 1 1970
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1713453518
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1713453518
transform 1 0 1784 0 1 1970
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1713453518
transform 1 0 1776 0 1 1970
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1713453518
transform 1 0 1736 0 1 1970
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1713453518
transform 1 0 1728 0 1 1970
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1713453518
transform 1 0 1720 0 1 1970
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1713453518
transform 1 0 1712 0 1 1970
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1713453518
transform 1 0 1704 0 1 1970
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1713453518
transform 1 0 1696 0 1 1970
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1713453518
transform 1 0 1648 0 1 1970
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1713453518
transform 1 0 1640 0 1 1970
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1713453518
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1713453518
transform 1 0 1584 0 1 1970
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1713453518
transform 1 0 1576 0 1 1970
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1713453518
transform 1 0 1568 0 1 1970
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1713453518
transform 1 0 1560 0 1 1970
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1713453518
transform 1 0 1552 0 1 1970
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1713453518
transform 1 0 1512 0 1 1970
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1713453518
transform 1 0 1504 0 1 1970
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1713453518
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1713453518
transform 1 0 1448 0 1 1970
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1713453518
transform 1 0 1440 0 1 1970
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1713453518
transform 1 0 1432 0 1 1970
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1713453518
transform 1 0 1424 0 1 1970
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1713453518
transform 1 0 1384 0 1 1970
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1713453518
transform 1 0 1376 0 1 1970
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1713453518
transform 1 0 1368 0 1 1970
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1713453518
transform 1 0 1360 0 1 1970
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1713453518
transform 1 0 1352 0 1 1970
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1713453518
transform 1 0 1344 0 1 1970
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1713453518
transform 1 0 1296 0 1 1970
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1713453518
transform 1 0 1288 0 1 1970
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1713453518
transform 1 0 1280 0 1 1970
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1713453518
transform 1 0 1232 0 1 1970
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1713453518
transform 1 0 1224 0 1 1970
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1713453518
transform 1 0 1216 0 1 1970
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1713453518
transform 1 0 1208 0 1 1970
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1713453518
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1713453518
transform 1 0 1152 0 1 1970
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1713453518
transform 1 0 1144 0 1 1970
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1713453518
transform 1 0 1136 0 1 1970
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1713453518
transform 1 0 1128 0 1 1970
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1713453518
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1713453518
transform 1 0 1064 0 1 1970
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1713453518
transform 1 0 1056 0 1 1970
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1713453518
transform 1 0 1016 0 1 1970
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1713453518
transform 1 0 1008 0 1 1970
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1713453518
transform 1 0 1000 0 1 1970
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1713453518
transform 1 0 992 0 1 1970
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1713453518
transform 1 0 888 0 1 1970
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1713453518
transform 1 0 880 0 1 1970
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1713453518
transform 1 0 872 0 1 1970
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1713453518
transform 1 0 864 0 1 1970
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1713453518
transform 1 0 856 0 1 1970
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1713453518
transform 1 0 792 0 1 1970
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1713453518
transform 1 0 752 0 1 1970
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1713453518
transform 1 0 744 0 1 1970
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1713453518
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1713453518
transform 1 0 696 0 1 1970
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1713453518
transform 1 0 656 0 1 1970
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1713453518
transform 1 0 648 0 1 1970
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1713453518
transform 1 0 640 0 1 1970
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1713453518
transform 1 0 600 0 1 1970
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1713453518
transform 1 0 592 0 1 1970
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1713453518
transform 1 0 552 0 1 1970
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1713453518
transform 1 0 544 0 1 1970
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1713453518
transform 1 0 536 0 1 1970
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1713453518
transform 1 0 528 0 1 1970
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1713453518
transform 1 0 480 0 1 1970
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1713453518
transform 1 0 432 0 1 1970
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1713453518
transform 1 0 424 0 1 1970
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1713453518
transform 1 0 416 0 1 1970
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1713453518
transform 1 0 408 0 1 1970
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1713453518
transform 1 0 304 0 1 1970
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1713453518
transform 1 0 296 0 1 1970
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1713453518
transform 1 0 288 0 1 1970
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1713453518
transform 1 0 208 0 1 1970
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1713453518
transform 1 0 200 0 1 1970
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1713453518
transform 1 0 192 0 1 1970
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1713453518
transform 1 0 184 0 1 1970
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1713453518
transform 1 0 80 0 1 1970
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1713453518
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1713453518
transform 1 0 3440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1713453518
transform 1 0 3432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1713453518
transform 1 0 3384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1713453518
transform 1 0 3376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1713453518
transform 1 0 3368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1713453518
transform 1 0 3360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1713453518
transform 1 0 3352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1713453518
transform 1 0 3344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1713453518
transform 1 0 3288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1713453518
transform 1 0 3280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1713453518
transform 1 0 3272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1713453518
transform 1 0 3264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1713453518
transform 1 0 3240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1713453518
transform 1 0 3232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1713453518
transform 1 0 3224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1713453518
transform 1 0 3192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1713453518
transform 1 0 3184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1713453518
transform 1 0 3176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1713453518
transform 1 0 3168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1713453518
transform 1 0 3128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1713453518
transform 1 0 3120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1713453518
transform 1 0 3112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1713453518
transform 1 0 3104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1713453518
transform 1 0 3096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1713453518
transform 1 0 3056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1713453518
transform 1 0 3048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1713453518
transform 1 0 3040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1713453518
transform 1 0 3032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1713453518
transform 1 0 3000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1713453518
transform 1 0 2992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1713453518
transform 1 0 2984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1713453518
transform 1 0 2976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1713453518
transform 1 0 2936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1713453518
transform 1 0 2928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1713453518
transform 1 0 2920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1713453518
transform 1 0 2912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1713453518
transform 1 0 2904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1713453518
transform 1 0 2864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1713453518
transform 1 0 2856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1713453518
transform 1 0 2848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1713453518
transform 1 0 2808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1713453518
transform 1 0 2800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1713453518
transform 1 0 2792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1713453518
transform 1 0 2784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1713453518
transform 1 0 2776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1713453518
transform 1 0 2728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1713453518
transform 1 0 2720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1713453518
transform 1 0 2712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1713453518
transform 1 0 2680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1713453518
transform 1 0 2672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1713453518
transform 1 0 2632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1713453518
transform 1 0 2624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1713453518
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1713453518
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1713453518
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1713453518
transform 1 0 2560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1713453518
transform 1 0 2552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1713453518
transform 1 0 2544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1713453518
transform 1 0 2496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1713453518
transform 1 0 2488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1713453518
transform 1 0 2480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1713453518
transform 1 0 2472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1713453518
transform 1 0 2464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1713453518
transform 1 0 2456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1713453518
transform 1 0 2448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1713453518
transform 1 0 2384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1713453518
transform 1 0 2376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1713453518
transform 1 0 2368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1713453518
transform 1 0 2360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1713453518
transform 1 0 2352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1713453518
transform 1 0 2312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1713453518
transform 1 0 2304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1713453518
transform 1 0 2296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1713453518
transform 1 0 2288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1713453518
transform 1 0 2280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1713453518
transform 1 0 2272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1713453518
transform 1 0 2240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1713453518
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1713453518
transform 1 0 2200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1713453518
transform 1 0 2192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1713453518
transform 1 0 2184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1713453518
transform 1 0 2176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1713453518
transform 1 0 2168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1713453518
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1713453518
transform 1 0 2112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1713453518
transform 1 0 2104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1713453518
transform 1 0 2096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1713453518
transform 1 0 2088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1713453518
transform 1 0 2080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1713453518
transform 1 0 2072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1713453518
transform 1 0 2064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1713453518
transform 1 0 2016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1713453518
transform 1 0 2008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1713453518
transform 1 0 2000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1713453518
transform 1 0 1992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1713453518
transform 1 0 1984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1713453518
transform 1 0 1976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1713453518
transform 1 0 1968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1713453518
transform 1 0 1944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1713453518
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1713453518
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1713453518
transform 1 0 1896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1713453518
transform 1 0 1888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1713453518
transform 1 0 1880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1713453518
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1713453518
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1713453518
transform 1 0 1824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1713453518
transform 1 0 1816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1713453518
transform 1 0 1808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1713453518
transform 1 0 1800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1713453518
transform 1 0 1792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1713453518
transform 1 0 1752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1713453518
transform 1 0 1744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1713453518
transform 1 0 1736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1713453518
transform 1 0 1728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1713453518
transform 1 0 1720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1713453518
transform 1 0 1688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1713453518
transform 1 0 1680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1713453518
transform 1 0 1672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1713453518
transform 1 0 1664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1713453518
transform 1 0 1656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1713453518
transform 1 0 1648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1713453518
transform 1 0 1616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1713453518
transform 1 0 1608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1713453518
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1713453518
transform 1 0 1576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1713453518
transform 1 0 1568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1713453518
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1713453518
transform 1 0 1520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1713453518
transform 1 0 1512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1713453518
transform 1 0 1504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1713453518
transform 1 0 1496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1713453518
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1713453518
transform 1 0 1432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1713453518
transform 1 0 1424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1713453518
transform 1 0 1416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1713453518
transform 1 0 1408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1713453518
transform 1 0 1400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1713453518
transform 1 0 1392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1713453518
transform 1 0 1336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1713453518
transform 1 0 1328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1713453518
transform 1 0 1320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1713453518
transform 1 0 1312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1713453518
transform 1 0 1304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1713453518
transform 1 0 1296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1713453518
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1713453518
transform 1 0 1240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1713453518
transform 1 0 1232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1713453518
transform 1 0 1224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1713453518
transform 1 0 1216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1713453518
transform 1 0 1208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1713453518
transform 1 0 1160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1713453518
transform 1 0 1152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1713453518
transform 1 0 1144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1713453518
transform 1 0 1136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1713453518
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1713453518
transform 1 0 1120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1713453518
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1713453518
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1713453518
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1713453518
transform 1 0 1008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1713453518
transform 1 0 1000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1713453518
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1713453518
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1713453518
transform 1 0 880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1713453518
transform 1 0 808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1713453518
transform 1 0 800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1713453518
transform 1 0 792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1713453518
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1713453518
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1713453518
transform 1 0 688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1713453518
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1713453518
transform 1 0 608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1713453518
transform 1 0 600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1713453518
transform 1 0 552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1713453518
transform 1 0 544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1713453518
transform 1 0 488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1713453518
transform 1 0 480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1713453518
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1713453518
transform 1 0 408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1713453518
transform 1 0 400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1713453518
transform 1 0 296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1713453518
transform 1 0 288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1713453518
transform 1 0 280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1713453518
transform 1 0 200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1713453518
transform 1 0 192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1713453518
transform 1 0 184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1713453518
transform 1 0 176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1713453518
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1713453518
transform 1 0 3440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1713453518
transform 1 0 3400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1713453518
transform 1 0 3392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1713453518
transform 1 0 3384 0 1 1770
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1713453518
transform 1 0 3376 0 1 1770
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1713453518
transform 1 0 3368 0 1 1770
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1713453518
transform 1 0 3320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1713453518
transform 1 0 3312 0 1 1770
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1713453518
transform 1 0 3304 0 1 1770
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1713453518
transform 1 0 3272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1713453518
transform 1 0 3264 0 1 1770
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1713453518
transform 1 0 3256 0 1 1770
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1713453518
transform 1 0 3248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1713453518
transform 1 0 3224 0 1 1770
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1713453518
transform 1 0 3200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1713453518
transform 1 0 3192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1713453518
transform 1 0 3184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1713453518
transform 1 0 3152 0 1 1770
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1713453518
transform 1 0 3144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1713453518
transform 1 0 3136 0 1 1770
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1713453518
transform 1 0 3128 0 1 1770
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1713453518
transform 1 0 3096 0 1 1770
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1713453518
transform 1 0 3056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1713453518
transform 1 0 3048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1713453518
transform 1 0 3040 0 1 1770
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1713453518
transform 1 0 3032 0 1 1770
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1713453518
transform 1 0 3024 0 1 1770
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1713453518
transform 1 0 3016 0 1 1770
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1713453518
transform 1 0 3008 0 1 1770
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1713453518
transform 1 0 2952 0 1 1770
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1713453518
transform 1 0 2944 0 1 1770
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1713453518
transform 1 0 2936 0 1 1770
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1713453518
transform 1 0 2928 0 1 1770
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1713453518
transform 1 0 2920 0 1 1770
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1713453518
transform 1 0 2880 0 1 1770
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1713453518
transform 1 0 2872 0 1 1770
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1713453518
transform 1 0 2824 0 1 1770
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1713453518
transform 1 0 2816 0 1 1770
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1713453518
transform 1 0 2808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1713453518
transform 1 0 2800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1713453518
transform 1 0 2792 0 1 1770
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1713453518
transform 1 0 2784 0 1 1770
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1713453518
transform 1 0 2744 0 1 1770
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1713453518
transform 1 0 2720 0 1 1770
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1713453518
transform 1 0 2712 0 1 1770
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1713453518
transform 1 0 2704 0 1 1770
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1713453518
transform 1 0 2680 0 1 1770
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1713453518
transform 1 0 2672 0 1 1770
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1713453518
transform 1 0 2664 0 1 1770
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1713453518
transform 1 0 2616 0 1 1770
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1713453518
transform 1 0 2608 0 1 1770
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1713453518
transform 1 0 2600 0 1 1770
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1713453518
transform 1 0 2592 0 1 1770
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1713453518
transform 1 0 2584 0 1 1770
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1713453518
transform 1 0 2552 0 1 1770
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1713453518
transform 1 0 2544 0 1 1770
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1713453518
transform 1 0 2536 0 1 1770
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1713453518
transform 1 0 2488 0 1 1770
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1713453518
transform 1 0 2480 0 1 1770
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1713453518
transform 1 0 2472 0 1 1770
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1713453518
transform 1 0 2464 0 1 1770
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1713453518
transform 1 0 2456 0 1 1770
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1713453518
transform 1 0 2432 0 1 1770
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1713453518
transform 1 0 2400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1713453518
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1713453518
transform 1 0 2384 0 1 1770
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1713453518
transform 1 0 2344 0 1 1770
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1713453518
transform 1 0 2336 0 1 1770
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1713453518
transform 1 0 2328 0 1 1770
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1713453518
transform 1 0 2320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1713453518
transform 1 0 2312 0 1 1770
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1713453518
transform 1 0 2280 0 1 1770
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1713453518
transform 1 0 2272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1713453518
transform 1 0 2264 0 1 1770
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1713453518
transform 1 0 2232 0 1 1770
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1713453518
transform 1 0 2224 0 1 1770
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1713453518
transform 1 0 2216 0 1 1770
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1713453518
transform 1 0 2208 0 1 1770
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1713453518
transform 1 0 2200 0 1 1770
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1713453518
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1713453518
transform 1 0 2184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1713453518
transform 1 0 2136 0 1 1770
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1713453518
transform 1 0 2128 0 1 1770
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1713453518
transform 1 0 2120 0 1 1770
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1713453518
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1713453518
transform 1 0 2104 0 1 1770
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1713453518
transform 1 0 2096 0 1 1770
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1713453518
transform 1 0 2088 0 1 1770
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1713453518
transform 1 0 2048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1713453518
transform 1 0 2040 0 1 1770
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1713453518
transform 1 0 2032 0 1 1770
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1713453518
transform 1 0 2024 0 1 1770
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1713453518
transform 1 0 2016 0 1 1770
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1713453518
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1713453518
transform 1 0 1968 0 1 1770
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1713453518
transform 1 0 1960 0 1 1770
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1713453518
transform 1 0 1952 0 1 1770
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1713453518
transform 1 0 1912 0 1 1770
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1713453518
transform 1 0 1904 0 1 1770
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1713453518
transform 1 0 1896 0 1 1770
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1713453518
transform 1 0 1888 0 1 1770
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1713453518
transform 1 0 1880 0 1 1770
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1713453518
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1713453518
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1713453518
transform 1 0 1824 0 1 1770
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1713453518
transform 1 0 1816 0 1 1770
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1713453518
transform 1 0 1808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1713453518
transform 1 0 1800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1713453518
transform 1 0 1792 0 1 1770
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1713453518
transform 1 0 1760 0 1 1770
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1713453518
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1713453518
transform 1 0 1744 0 1 1770
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1713453518
transform 1 0 1736 0 1 1770
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1713453518
transform 1 0 1728 0 1 1770
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1713453518
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1713453518
transform 1 0 1688 0 1 1770
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1713453518
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1713453518
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1713453518
transform 1 0 1664 0 1 1770
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1713453518
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1713453518
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1713453518
transform 1 0 1608 0 1 1770
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1713453518
transform 1 0 1600 0 1 1770
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1713453518
transform 1 0 1552 0 1 1770
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1713453518
transform 1 0 1544 0 1 1770
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1713453518
transform 1 0 1536 0 1 1770
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1713453518
transform 1 0 1528 0 1 1770
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1713453518
transform 1 0 1488 0 1 1770
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1713453518
transform 1 0 1480 0 1 1770
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1713453518
transform 1 0 1448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1713453518
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1713453518
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1713453518
transform 1 0 1424 0 1 1770
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1713453518
transform 1 0 1376 0 1 1770
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1713453518
transform 1 0 1368 0 1 1770
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1713453518
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1713453518
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1713453518
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1713453518
transform 1 0 1288 0 1 1770
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1713453518
transform 1 0 1280 0 1 1770
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1713453518
transform 1 0 1272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1713453518
transform 1 0 1240 0 1 1770
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1713453518
transform 1 0 1232 0 1 1770
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1713453518
transform 1 0 1224 0 1 1770
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1713453518
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1713453518
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1713453518
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1713453518
transform 1 0 1136 0 1 1770
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1713453518
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1713453518
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1713453518
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1713453518
transform 1 0 936 0 1 1770
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1713453518
transform 1 0 928 0 1 1770
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1713453518
transform 1 0 880 0 1 1770
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1713453518
transform 1 0 872 0 1 1770
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1713453518
transform 1 0 768 0 1 1770
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1713453518
transform 1 0 760 0 1 1770
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1713453518
transform 1 0 752 0 1 1770
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1713453518
transform 1 0 744 0 1 1770
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1713453518
transform 1 0 736 0 1 1770
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1713453518
transform 1 0 656 0 1 1770
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1713453518
transform 1 0 648 0 1 1770
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1713453518
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1713453518
transform 1 0 632 0 1 1770
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1713453518
transform 1 0 624 0 1 1770
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1713453518
transform 1 0 552 0 1 1770
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1713453518
transform 1 0 544 0 1 1770
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1713453518
transform 1 0 536 0 1 1770
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1713453518
transform 1 0 528 0 1 1770
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1713453518
transform 1 0 464 0 1 1770
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1713453518
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1713453518
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1713453518
transform 1 0 440 0 1 1770
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1713453518
transform 1 0 392 0 1 1770
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1713453518
transform 1 0 384 0 1 1770
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1713453518
transform 1 0 376 0 1 1770
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1713453518
transform 1 0 320 0 1 1770
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1713453518
transform 1 0 312 0 1 1770
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1713453518
transform 1 0 304 0 1 1770
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1713453518
transform 1 0 200 0 1 1770
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1713453518
transform 1 0 192 0 1 1770
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1713453518
transform 1 0 184 0 1 1770
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1713453518
transform 1 0 176 0 1 1770
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1713453518
transform 1 0 168 0 1 1770
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1713453518
transform 1 0 136 0 1 1770
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1713453518
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1713453518
transform 1 0 120 0 1 1770
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1713453518
transform 1 0 112 0 1 1770
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1713453518
transform 1 0 104 0 1 1770
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1713453518
transform 1 0 96 0 1 1770
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1713453518
transform 1 0 88 0 1 1770
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1713453518
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1713453518
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1713453518
transform 1 0 3440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1713453518
transform 1 0 3432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1713453518
transform 1 0 3408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1713453518
transform 1 0 3400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1713453518
transform 1 0 3352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1713453518
transform 1 0 3344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1713453518
transform 1 0 3336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1713453518
transform 1 0 3328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1713453518
transform 1 0 3320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1713453518
transform 1 0 3288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1713453518
transform 1 0 3280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1713453518
transform 1 0 3248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1713453518
transform 1 0 3240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1713453518
transform 1 0 3232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1713453518
transform 1 0 3224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1713453518
transform 1 0 3216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1713453518
transform 1 0 3208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1713453518
transform 1 0 3168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1713453518
transform 1 0 3160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1713453518
transform 1 0 3152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1713453518
transform 1 0 3144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1713453518
transform 1 0 3136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1713453518
transform 1 0 3128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1713453518
transform 1 0 3096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1713453518
transform 1 0 3088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1713453518
transform 1 0 3080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1713453518
transform 1 0 3072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1713453518
transform 1 0 3024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1713453518
transform 1 0 3016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1713453518
transform 1 0 3008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1713453518
transform 1 0 3000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1713453518
transform 1 0 2992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1713453518
transform 1 0 2984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1713453518
transform 1 0 2944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1713453518
transform 1 0 2912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1713453518
transform 1 0 2904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1713453518
transform 1 0 2896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1713453518
transform 1 0 2864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1713453518
transform 1 0 2856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1713453518
transform 1 0 2848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1713453518
transform 1 0 2840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1713453518
transform 1 0 2832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1713453518
transform 1 0 2824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1713453518
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1713453518
transform 1 0 2744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1713453518
transform 1 0 2736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1713453518
transform 1 0 2728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1713453518
transform 1 0 2720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1713453518
transform 1 0 2680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1713453518
transform 1 0 2640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1713453518
transform 1 0 2632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1713453518
transform 1 0 2624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1713453518
transform 1 0 2616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1713453518
transform 1 0 2608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1713453518
transform 1 0 2600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1713453518
transform 1 0 2544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1713453518
transform 1 0 2536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1713453518
transform 1 0 2528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1713453518
transform 1 0 2520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1713453518
transform 1 0 2472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1713453518
transform 1 0 2464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1713453518
transform 1 0 2456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1713453518
transform 1 0 2448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1713453518
transform 1 0 2400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1713453518
transform 1 0 2392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1713453518
transform 1 0 2384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1713453518
transform 1 0 2376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1713453518
transform 1 0 2336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1713453518
transform 1 0 2328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1713453518
transform 1 0 2320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1713453518
transform 1 0 2312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1713453518
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1713453518
transform 1 0 2272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1713453518
transform 1 0 2264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1713453518
transform 1 0 2256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1713453518
transform 1 0 2216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1713453518
transform 1 0 2208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1713453518
transform 1 0 2200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1713453518
transform 1 0 2192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1713453518
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1713453518
transform 1 0 2176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1713453518
transform 1 0 2128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1713453518
transform 1 0 2120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1713453518
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1713453518
transform 1 0 2104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1713453518
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1713453518
transform 1 0 2048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1713453518
transform 1 0 2040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3130
timestamp 1713453518
transform 1 0 2032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1713453518
transform 1 0 2024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1713453518
transform 1 0 2016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1713453518
transform 1 0 1976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1713453518
transform 1 0 1968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1713453518
transform 1 0 1960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3136
timestamp 1713453518
transform 1 0 1952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1713453518
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1713453518
transform 1 0 1912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1713453518
transform 1 0 1904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1713453518
transform 1 0 1896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1713453518
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1713453518
transform 1 0 1856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1713453518
transform 1 0 1848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1713453518
transform 1 0 1840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1713453518
transform 1 0 1832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1713453518
transform 1 0 1792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1713453518
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1713453518
transform 1 0 1776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1713453518
transform 1 0 1768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1713453518
transform 1 0 1760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1713453518
transform 1 0 1752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1713453518
transform 1 0 1720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1713453518
transform 1 0 1712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1713453518
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1713453518
transform 1 0 1672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1713453518
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1713453518
transform 1 0 1656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1713453518
transform 1 0 1648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1713453518
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1713453518
transform 1 0 1600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1713453518
transform 1 0 1592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1713453518
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1713453518
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1713453518
transform 1 0 1536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1713453518
transform 1 0 1528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1713453518
transform 1 0 1480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1713453518
transform 1 0 1472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1713453518
transform 1 0 1464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1713453518
transform 1 0 1432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1713453518
transform 1 0 1424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1713453518
transform 1 0 1416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1713453518
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1713453518
transform 1 0 1360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1713453518
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1713453518
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1713453518
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1713453518
transform 1 0 1328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1713453518
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1713453518
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1713453518
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1713453518
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1713453518
transform 1 0 1224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1713453518
transform 1 0 1216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1713453518
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1713453518
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1713453518
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1713453518
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1713453518
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1713453518
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1713453518
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1713453518
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1713453518
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1713453518
transform 1 0 1040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1713453518
transform 1 0 936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1713453518
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1713453518
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1713453518
transform 1 0 832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1713453518
transform 1 0 824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1713453518
transform 1 0 816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1713453518
transform 1 0 712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1713453518
transform 1 0 704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1713453518
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1713453518
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1713453518
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1713453518
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1713453518
transform 1 0 576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1713453518
transform 1 0 568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1713453518
transform 1 0 560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1713453518
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1713453518
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1713453518
transform 1 0 472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1713453518
transform 1 0 400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1713453518
transform 1 0 392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1713453518
transform 1 0 384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1713453518
transform 1 0 376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1713453518
transform 1 0 368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1713453518
transform 1 0 296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1713453518
transform 1 0 288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1713453518
transform 1 0 280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1713453518
transform 1 0 272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1713453518
transform 1 0 264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1713453518
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1713453518
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1713453518
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1713453518
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1713453518
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1713453518
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1713453518
transform 1 0 3440 0 1 1570
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1713453518
transform 1 0 3400 0 1 1570
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1713453518
transform 1 0 3392 0 1 1570
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1713453518
transform 1 0 3384 0 1 1570
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1713453518
transform 1 0 3376 0 1 1570
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1713453518
transform 1 0 3328 0 1 1570
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1713453518
transform 1 0 3320 0 1 1570
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1713453518
transform 1 0 3288 0 1 1570
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1713453518
transform 1 0 3280 0 1 1570
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1713453518
transform 1 0 3272 0 1 1570
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1713453518
transform 1 0 3240 0 1 1570
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1713453518
transform 1 0 3232 0 1 1570
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1713453518
transform 1 0 3224 0 1 1570
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1713453518
transform 1 0 3184 0 1 1570
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1713453518
transform 1 0 3176 0 1 1570
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1713453518
transform 1 0 3168 0 1 1570
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1713453518
transform 1 0 3160 0 1 1570
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1713453518
transform 1 0 3152 0 1 1570
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1713453518
transform 1 0 3112 0 1 1570
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1713453518
transform 1 0 3088 0 1 1570
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1713453518
transform 1 0 3080 0 1 1570
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1713453518
transform 1 0 3072 0 1 1570
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1713453518
transform 1 0 3064 0 1 1570
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1713453518
transform 1 0 3032 0 1 1570
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1713453518
transform 1 0 3024 0 1 1570
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1713453518
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1713453518
transform 1 0 2976 0 1 1570
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1713453518
transform 1 0 2968 0 1 1570
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1713453518
transform 1 0 2960 0 1 1570
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1713453518
transform 1 0 2952 0 1 1570
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1713453518
transform 1 0 2912 0 1 1570
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1713453518
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1713453518
transform 1 0 2864 0 1 1570
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1713453518
transform 1 0 2856 0 1 1570
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1713453518
transform 1 0 2848 0 1 1570
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1713453518
transform 1 0 2816 0 1 1570
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1713453518
transform 1 0 2808 0 1 1570
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1713453518
transform 1 0 2760 0 1 1570
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1713453518
transform 1 0 2752 0 1 1570
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1713453518
transform 1 0 2744 0 1 1570
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1713453518
transform 1 0 2736 0 1 1570
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1713453518
transform 1 0 2728 0 1 1570
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1713453518
transform 1 0 2688 0 1 1570
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1713453518
transform 1 0 2656 0 1 1570
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1713453518
transform 1 0 2632 0 1 1570
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1713453518
transform 1 0 2624 0 1 1570
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1713453518
transform 1 0 2616 0 1 1570
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1713453518
transform 1 0 2608 0 1 1570
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1713453518
transform 1 0 2600 0 1 1570
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1713453518
transform 1 0 2536 0 1 1570
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1713453518
transform 1 0 2528 0 1 1570
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1713453518
transform 1 0 2520 0 1 1570
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1713453518
transform 1 0 2480 0 1 1570
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1713453518
transform 1 0 2472 0 1 1570
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1713453518
transform 1 0 2464 0 1 1570
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1713453518
transform 1 0 2456 0 1 1570
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1713453518
transform 1 0 2384 0 1 1570
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1713453518
transform 1 0 2376 0 1 1570
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1713453518
transform 1 0 2368 0 1 1570
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1713453518
transform 1 0 2360 0 1 1570
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1713453518
transform 1 0 2352 0 1 1570
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1713453518
transform 1 0 2344 0 1 1570
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1713453518
transform 1 0 2280 0 1 1570
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1713453518
transform 1 0 2272 0 1 1570
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1713453518
transform 1 0 2264 0 1 1570
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1713453518
transform 1 0 2256 0 1 1570
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1713453518
transform 1 0 2248 0 1 1570
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1713453518
transform 1 0 2240 0 1 1570
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1713453518
transform 1 0 2168 0 1 1570
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1713453518
transform 1 0 2160 0 1 1570
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1713453518
transform 1 0 2152 0 1 1570
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1713453518
transform 1 0 2144 0 1 1570
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1713453518
transform 1 0 2096 0 1 1570
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1713453518
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1713453518
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1713453518
transform 1 0 2040 0 1 1570
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1713453518
transform 1 0 2032 0 1 1570
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1713453518
transform 1 0 2024 0 1 1570
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1713453518
transform 1 0 2016 0 1 1570
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1713453518
transform 1 0 1976 0 1 1570
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1713453518
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1713453518
transform 1 0 1928 0 1 1570
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1713453518
transform 1 0 1920 0 1 1570
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1713453518
transform 1 0 1912 0 1 1570
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1713453518
transform 1 0 1904 0 1 1570
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1713453518
transform 1 0 1856 0 1 1570
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1713453518
transform 1 0 1848 0 1 1570
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1713453518
transform 1 0 1840 0 1 1570
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1713453518
transform 1 0 1832 0 1 1570
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1713453518
transform 1 0 1824 0 1 1570
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1713453518
transform 1 0 1816 0 1 1570
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1713453518
transform 1 0 1808 0 1 1570
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1713453518
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1713453518
transform 1 0 1736 0 1 1570
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1713453518
transform 1 0 1728 0 1 1570
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1713453518
transform 1 0 1720 0 1 1570
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1713453518
transform 1 0 1712 0 1 1570
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1713453518
transform 1 0 1704 0 1 1570
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1713453518
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1713453518
transform 1 0 1640 0 1 1570
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1713453518
transform 1 0 1632 0 1 1570
box -8 -3 16 105
use FILL  FILL_3329
timestamp 1713453518
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1713453518
transform 1 0 1616 0 1 1570
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1713453518
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1713453518
transform 1 0 1560 0 1 1570
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1713453518
transform 1 0 1552 0 1 1570
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1713453518
transform 1 0 1512 0 1 1570
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1713453518
transform 1 0 1504 0 1 1570
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1713453518
transform 1 0 1496 0 1 1570
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1713453518
transform 1 0 1456 0 1 1570
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1713453518
transform 1 0 1448 0 1 1570
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1713453518
transform 1 0 1440 0 1 1570
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1713453518
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1713453518
transform 1 0 1384 0 1 1570
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1713453518
transform 1 0 1376 0 1 1570
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1713453518
transform 1 0 1352 0 1 1570
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1713453518
transform 1 0 1344 0 1 1570
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1713453518
transform 1 0 1336 0 1 1570
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1713453518
transform 1 0 1328 0 1 1570
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1713453518
transform 1 0 1272 0 1 1570
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1713453518
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1713453518
transform 1 0 1256 0 1 1570
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1713453518
transform 1 0 1248 0 1 1570
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1713453518
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1713453518
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1713453518
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1713453518
transform 1 0 1144 0 1 1570
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1713453518
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1713453518
transform 1 0 1128 0 1 1570
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1713453518
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1713453518
transform 1 0 1056 0 1 1570
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1713453518
transform 1 0 1048 0 1 1570
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1713453518
transform 1 0 1040 0 1 1570
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1713453518
transform 1 0 1032 0 1 1570
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1713453518
transform 1 0 976 0 1 1570
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1713453518
transform 1 0 968 0 1 1570
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1713453518
transform 1 0 960 0 1 1570
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1713453518
transform 1 0 888 0 1 1570
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1713453518
transform 1 0 880 0 1 1570
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1713453518
transform 1 0 872 0 1 1570
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1713453518
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1713453518
transform 1 0 760 0 1 1570
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1713453518
transform 1 0 752 0 1 1570
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1713453518
transform 1 0 744 0 1 1570
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1713453518
transform 1 0 664 0 1 1570
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1713453518
transform 1 0 656 0 1 1570
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1713453518
transform 1 0 648 0 1 1570
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1713453518
transform 1 0 568 0 1 1570
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1713453518
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1713453518
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1713453518
transform 1 0 544 0 1 1570
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1713453518
transform 1 0 504 0 1 1570
box -8 -3 16 105
use FILL  FILL_3380
timestamp 1713453518
transform 1 0 496 0 1 1570
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1713453518
transform 1 0 432 0 1 1570
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1713453518
transform 1 0 424 0 1 1570
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1713453518
transform 1 0 416 0 1 1570
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1713453518
transform 1 0 408 0 1 1570
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1713453518
transform 1 0 360 0 1 1570
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1713453518
transform 1 0 304 0 1 1570
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1713453518
transform 1 0 296 0 1 1570
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1713453518
transform 1 0 288 0 1 1570
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1713453518
transform 1 0 184 0 1 1570
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1713453518
transform 1 0 176 0 1 1570
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1713453518
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1713453518
transform 1 0 3440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1713453518
transform 1 0 3432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1713453518
transform 1 0 3424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1713453518
transform 1 0 3368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1713453518
transform 1 0 3360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1713453518
transform 1 0 3352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1713453518
transform 1 0 3304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3399
timestamp 1713453518
transform 1 0 3296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1713453518
transform 1 0 3288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1713453518
transform 1 0 3280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1713453518
transform 1 0 3232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1713453518
transform 1 0 3224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1713453518
transform 1 0 3216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1713453518
transform 1 0 3208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1713453518
transform 1 0 3200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1713453518
transform 1 0 3168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1713453518
transform 1 0 3160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1713453518
transform 1 0 3152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1713453518
transform 1 0 3120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1713453518
transform 1 0 3112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1713453518
transform 1 0 3104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1713453518
transform 1 0 3064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1713453518
transform 1 0 3056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1713453518
transform 1 0 3048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1713453518
transform 1 0 3040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1713453518
transform 1 0 3000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1713453518
transform 1 0 2992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1713453518
transform 1 0 2984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1713453518
transform 1 0 2952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1713453518
transform 1 0 2944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1713453518
transform 1 0 2936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1713453518
transform 1 0 2928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1713453518
transform 1 0 2880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1713453518
transform 1 0 2872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1713453518
transform 1 0 2864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1713453518
transform 1 0 2856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1713453518
transform 1 0 2824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1713453518
transform 1 0 2816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1713453518
transform 1 0 2776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1713453518
transform 1 0 2768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1713453518
transform 1 0 2760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1713453518
transform 1 0 2752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1713453518
transform 1 0 2744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1713453518
transform 1 0 2704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1713453518
transform 1 0 2696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1713453518
transform 1 0 2664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1713453518
transform 1 0 2656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1713453518
transform 1 0 2648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1713453518
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1713453518
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1713453518
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1713453518
transform 1 0 2560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1713453518
transform 1 0 2552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1713453518
transform 1 0 2544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1713453518
transform 1 0 2536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1713453518
transform 1 0 2488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3448
timestamp 1713453518
transform 1 0 2480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1713453518
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1713453518
transform 1 0 2432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1713453518
transform 1 0 2424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1713453518
transform 1 0 2416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1713453518
transform 1 0 2408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1713453518
transform 1 0 2400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1713453518
transform 1 0 2352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1713453518
transform 1 0 2344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1713453518
transform 1 0 2336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3458
timestamp 1713453518
transform 1 0 2328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1713453518
transform 1 0 2296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1713453518
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1713453518
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1713453518
transform 1 0 2232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1713453518
transform 1 0 2224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3464
timestamp 1713453518
transform 1 0 2216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1713453518
transform 1 0 2208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1713453518
transform 1 0 2200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1713453518
transform 1 0 2192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1713453518
transform 1 0 2152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3469
timestamp 1713453518
transform 1 0 2144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1713453518
transform 1 0 2112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1713453518
transform 1 0 2104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1713453518
transform 1 0 2096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1713453518
transform 1 0 2064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1713453518
transform 1 0 2056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1713453518
transform 1 0 2048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1713453518
transform 1 0 2040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1713453518
transform 1 0 2032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1713453518
transform 1 0 1984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1713453518
transform 1 0 1976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1713453518
transform 1 0 1968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1713453518
transform 1 0 1960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1713453518
transform 1 0 1928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3483
timestamp 1713453518
transform 1 0 1920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1713453518
transform 1 0 1912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1713453518
transform 1 0 1872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1713453518
transform 1 0 1864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1713453518
transform 1 0 1856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1713453518
transform 1 0 1848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1713453518
transform 1 0 1840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1713453518
transform 1 0 1800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1713453518
transform 1 0 1792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1713453518
transform 1 0 1784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1713453518
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1713453518
transform 1 0 1736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3495
timestamp 1713453518
transform 1 0 1728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1713453518
transform 1 0 1720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1713453518
transform 1 0 1712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1713453518
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1713453518
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1713453518
transform 1 0 1640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1713453518
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1713453518
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1713453518
transform 1 0 1616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1713453518
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1713453518
transform 1 0 1576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1713453518
transform 1 0 1568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1713453518
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3508
timestamp 1713453518
transform 1 0 1552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1713453518
transform 1 0 1512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1713453518
transform 1 0 1504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1713453518
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1713453518
transform 1 0 1464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1713453518
transform 1 0 1456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1713453518
transform 1 0 1448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1713453518
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1713453518
transform 1 0 1408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1713453518
transform 1 0 1400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1713453518
transform 1 0 1392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1713453518
transform 1 0 1352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1713453518
transform 1 0 1344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1713453518
transform 1 0 1336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1713453518
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1713453518
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1713453518
transform 1 0 1288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3525
timestamp 1713453518
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1713453518
transform 1 0 1240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1713453518
transform 1 0 1232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1713453518
transform 1 0 1224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1713453518
transform 1 0 1216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1713453518
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1713453518
transform 1 0 1168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1713453518
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1713453518
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1713453518
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1713453518
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1713453518
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1713453518
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1713453518
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1713453518
transform 1 0 1008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1713453518
transform 1 0 1000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1713453518
transform 1 0 992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1713453518
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1713453518
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3544
timestamp 1713453518
transform 1 0 800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1713453518
transform 1 0 792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1713453518
transform 1 0 784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1713453518
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1713453518
transform 1 0 728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1713453518
transform 1 0 688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1713453518
transform 1 0 680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1713453518
transform 1 0 672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1713453518
transform 1 0 664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1713453518
transform 1 0 656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1713453518
transform 1 0 592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1713453518
transform 1 0 584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1713453518
transform 1 0 544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1713453518
transform 1 0 536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1713453518
transform 1 0 528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1713453518
transform 1 0 472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1713453518
transform 1 0 464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1713453518
transform 1 0 424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1713453518
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1713453518
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1713453518
transform 1 0 360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1713453518
transform 1 0 352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1713453518
transform 1 0 248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3567
timestamp 1713453518
transform 1 0 240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1713453518
transform 1 0 232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1713453518
transform 1 0 224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1713453518
transform 1 0 216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1713453518
transform 1 0 184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1713453518
transform 1 0 176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1713453518
transform 1 0 120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1713453518
transform 1 0 112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3575
timestamp 1713453518
transform 1 0 104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1713453518
transform 1 0 96 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1713453518
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1713453518
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1713453518
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1713453518
transform 1 0 3440 0 1 1370
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1713453518
transform 1 0 3432 0 1 1370
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1713453518
transform 1 0 3424 0 1 1370
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1713453518
transform 1 0 3360 0 1 1370
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1713453518
transform 1 0 3352 0 1 1370
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1713453518
transform 1 0 3320 0 1 1370
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1713453518
transform 1 0 3312 0 1 1370
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1713453518
transform 1 0 3304 0 1 1370
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1713453518
transform 1 0 3248 0 1 1370
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1713453518
transform 1 0 3240 0 1 1370
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1713453518
transform 1 0 3232 0 1 1370
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1713453518
transform 1 0 3224 0 1 1370
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1713453518
transform 1 0 3216 0 1 1370
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1713453518
transform 1 0 3208 0 1 1370
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1713453518
transform 1 0 3168 0 1 1370
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1713453518
transform 1 0 3160 0 1 1370
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1713453518
transform 1 0 3120 0 1 1370
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1713453518
transform 1 0 3112 0 1 1370
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1713453518
transform 1 0 3104 0 1 1370
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1713453518
transform 1 0 3096 0 1 1370
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1713453518
transform 1 0 3088 0 1 1370
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1713453518
transform 1 0 3048 0 1 1370
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1713453518
transform 1 0 3040 0 1 1370
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1713453518
transform 1 0 3016 0 1 1370
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1713453518
transform 1 0 3008 0 1 1370
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1713453518
transform 1 0 3000 0 1 1370
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1713453518
transform 1 0 2992 0 1 1370
box -8 -3 16 105
use FILL  FILL_3607
timestamp 1713453518
transform 1 0 2984 0 1 1370
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1713453518
transform 1 0 2936 0 1 1370
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1713453518
transform 1 0 2928 0 1 1370
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1713453518
transform 1 0 2920 0 1 1370
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1713453518
transform 1 0 2912 0 1 1370
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1713453518
transform 1 0 2904 0 1 1370
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1713453518
transform 1 0 2856 0 1 1370
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1713453518
transform 1 0 2848 0 1 1370
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1713453518
transform 1 0 2840 0 1 1370
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1713453518
transform 1 0 2808 0 1 1370
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1713453518
transform 1 0 2800 0 1 1370
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1713453518
transform 1 0 2792 0 1 1370
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1713453518
transform 1 0 2784 0 1 1370
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1713453518
transform 1 0 2776 0 1 1370
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1713453518
transform 1 0 2768 0 1 1370
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1713453518
transform 1 0 2720 0 1 1370
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1713453518
transform 1 0 2712 0 1 1370
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1713453518
transform 1 0 2704 0 1 1370
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1713453518
transform 1 0 2696 0 1 1370
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1713453518
transform 1 0 2688 0 1 1370
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1713453518
transform 1 0 2648 0 1 1370
box -8 -3 16 105
use FILL  FILL_3628
timestamp 1713453518
transform 1 0 2640 0 1 1370
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1713453518
transform 1 0 2632 0 1 1370
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1713453518
transform 1 0 2592 0 1 1370
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1713453518
transform 1 0 2584 0 1 1370
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1713453518
transform 1 0 2576 0 1 1370
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1713453518
transform 1 0 2568 0 1 1370
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1713453518
transform 1 0 2528 0 1 1370
box -8 -3 16 105
use FILL  FILL_3635
timestamp 1713453518
transform 1 0 2520 0 1 1370
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1713453518
transform 1 0 2512 0 1 1370
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1713453518
transform 1 0 2504 0 1 1370
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1713453518
transform 1 0 2464 0 1 1370
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1713453518
transform 1 0 2456 0 1 1370
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1713453518
transform 1 0 2448 0 1 1370
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1713453518
transform 1 0 2440 0 1 1370
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1713453518
transform 1 0 2432 0 1 1370
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1713453518
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1713453518
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_3645
timestamp 1713453518
transform 1 0 2360 0 1 1370
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1713453518
transform 1 0 2352 0 1 1370
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1713453518
transform 1 0 2344 0 1 1370
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1713453518
transform 1 0 2336 0 1 1370
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1713453518
transform 1 0 2288 0 1 1370
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1713453518
transform 1 0 2280 0 1 1370
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1713453518
transform 1 0 2272 0 1 1370
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1713453518
transform 1 0 2264 0 1 1370
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1713453518
transform 1 0 2232 0 1 1370
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1713453518
transform 1 0 2224 0 1 1370
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1713453518
transform 1 0 2216 0 1 1370
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1713453518
transform 1 0 2208 0 1 1370
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1713453518
transform 1 0 2200 0 1 1370
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1713453518
transform 1 0 2152 0 1 1370
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1713453518
transform 1 0 2144 0 1 1370
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1713453518
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1713453518
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1713453518
transform 1 0 2088 0 1 1370
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1713453518
transform 1 0 2080 0 1 1370
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1713453518
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_3665
timestamp 1713453518
transform 1 0 2024 0 1 1370
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1713453518
transform 1 0 2016 0 1 1370
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1713453518
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1713453518
transform 1 0 2000 0 1 1370
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1713453518
transform 1 0 1992 0 1 1370
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1713453518
transform 1 0 1960 0 1 1370
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1713453518
transform 1 0 1952 0 1 1370
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1713453518
transform 1 0 1944 0 1 1370
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1713453518
transform 1 0 1936 0 1 1370
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1713453518
transform 1 0 1888 0 1 1370
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1713453518
transform 1 0 1880 0 1 1370
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1713453518
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use FILL  FILL_3677
timestamp 1713453518
transform 1 0 1864 0 1 1370
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1713453518
transform 1 0 1856 0 1 1370
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1713453518
transform 1 0 1848 0 1 1370
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1713453518
transform 1 0 1808 0 1 1370
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1713453518
transform 1 0 1800 0 1 1370
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1713453518
transform 1 0 1792 0 1 1370
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1713453518
transform 1 0 1784 0 1 1370
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1713453518
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1713453518
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1713453518
transform 1 0 1728 0 1 1370
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1713453518
transform 1 0 1720 0 1 1370
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1713453518
transform 1 0 1712 0 1 1370
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1713453518
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1713453518
transform 1 0 1648 0 1 1370
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1713453518
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1713453518
transform 1 0 1632 0 1 1370
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1713453518
transform 1 0 1624 0 1 1370
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1713453518
transform 1 0 1616 0 1 1370
box -8 -3 16 105
use FILL  FILL_3695
timestamp 1713453518
transform 1 0 1608 0 1 1370
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1713453518
transform 1 0 1536 0 1 1370
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1713453518
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1713453518
transform 1 0 1520 0 1 1370
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1713453518
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1713453518
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1713453518
transform 1 0 1496 0 1 1370
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1713453518
transform 1 0 1464 0 1 1370
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1713453518
transform 1 0 1424 0 1 1370
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1713453518
transform 1 0 1416 0 1 1370
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1713453518
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1713453518
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1713453518
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1713453518
transform 1 0 1360 0 1 1370
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1713453518
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1713453518
transform 1 0 1344 0 1 1370
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1713453518
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1713453518
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1713453518
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1713453518
transform 1 0 1272 0 1 1370
box -8 -3 16 105
use FILL  FILL_3715
timestamp 1713453518
transform 1 0 1264 0 1 1370
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1713453518
transform 1 0 1200 0 1 1370
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1713453518
transform 1 0 1192 0 1 1370
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1713453518
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1713453518
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_3720
timestamp 1713453518
transform 1 0 1168 0 1 1370
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1713453518
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1713453518
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1713453518
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1713453518
transform 1 0 1072 0 1 1370
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1713453518
transform 1 0 1064 0 1 1370
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1713453518
transform 1 0 1056 0 1 1370
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1713453518
transform 1 0 1048 0 1 1370
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1713453518
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1713453518
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_3730
timestamp 1713453518
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1713453518
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1713453518
transform 1 0 848 0 1 1370
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1713453518
transform 1 0 840 0 1 1370
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1713453518
transform 1 0 832 0 1 1370
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1713453518
transform 1 0 824 0 1 1370
box -8 -3 16 105
use FILL  FILL_3736
timestamp 1713453518
transform 1 0 752 0 1 1370
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1713453518
transform 1 0 744 0 1 1370
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1713453518
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1713453518
transform 1 0 688 0 1 1370
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1713453518
transform 1 0 680 0 1 1370
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1713453518
transform 1 0 624 0 1 1370
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1713453518
transform 1 0 616 0 1 1370
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1713453518
transform 1 0 608 0 1 1370
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1713453518
transform 1 0 520 0 1 1370
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1713453518
transform 1 0 512 0 1 1370
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1713453518
transform 1 0 504 0 1 1370
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1713453518
transform 1 0 496 0 1 1370
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1713453518
transform 1 0 400 0 1 1370
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1713453518
transform 1 0 392 0 1 1370
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1713453518
transform 1 0 288 0 1 1370
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1713453518
transform 1 0 280 0 1 1370
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1713453518
transform 1 0 272 0 1 1370
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1713453518
transform 1 0 264 0 1 1370
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1713453518
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1713453518
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1713453518
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_3757
timestamp 1713453518
transform 1 0 3440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1713453518
transform 1 0 3432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1713453518
transform 1 0 3424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1713453518
transform 1 0 3376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1713453518
transform 1 0 3368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1713453518
transform 1 0 3360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1713453518
transform 1 0 3352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1713453518
transform 1 0 3320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1713453518
transform 1 0 3312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1713453518
transform 1 0 3304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1713453518
transform 1 0 3296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3768
timestamp 1713453518
transform 1 0 3288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1713453518
transform 1 0 3240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1713453518
transform 1 0 3232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1713453518
transform 1 0 3224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1713453518
transform 1 0 3216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1713453518
transform 1 0 3208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1713453518
transform 1 0 3200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1713453518
transform 1 0 3192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1713453518
transform 1 0 3184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1713453518
transform 1 0 3136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1713453518
transform 1 0 3128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1713453518
transform 1 0 3120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3780
timestamp 1713453518
transform 1 0 3112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1713453518
transform 1 0 3104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1713453518
transform 1 0 3072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1713453518
transform 1 0 3064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1713453518
transform 1 0 3056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3785
timestamp 1713453518
transform 1 0 3048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1713453518
transform 1 0 3040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1713453518
transform 1 0 3000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1713453518
transform 1 0 2992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3789
timestamp 1713453518
transform 1 0 2984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1713453518
transform 1 0 2976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1713453518
transform 1 0 2968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1713453518
transform 1 0 2960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1713453518
transform 1 0 2912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1713453518
transform 1 0 2904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1713453518
transform 1 0 2896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1713453518
transform 1 0 2888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1713453518
transform 1 0 2856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1713453518
transform 1 0 2848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1713453518
transform 1 0 2840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1713453518
transform 1 0 2832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1713453518
transform 1 0 2824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1713453518
transform 1 0 2776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1713453518
transform 1 0 2768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1713453518
transform 1 0 2760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1713453518
transform 1 0 2752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3806
timestamp 1713453518
transform 1 0 2712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1713453518
transform 1 0 2704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1713453518
transform 1 0 2696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1713453518
transform 1 0 2656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1713453518
transform 1 0 2648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1713453518
transform 1 0 2640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1713453518
transform 1 0 2632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1713453518
transform 1 0 2624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1713453518
transform 1 0 2600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1713453518
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1713453518
transform 1 0 2552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3817
timestamp 1713453518
transform 1 0 2544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1713453518
transform 1 0 2536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1713453518
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1713453518
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1713453518
transform 1 0 2480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1713453518
transform 1 0 2448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1713453518
transform 1 0 2440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1713453518
transform 1 0 2432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3825
timestamp 1713453518
transform 1 0 2384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1713453518
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1713453518
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1713453518
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1713453518
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1713453518
transform 1 0 2344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1713453518
transform 1 0 2296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1713453518
transform 1 0 2288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1713453518
transform 1 0 2280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1713453518
transform 1 0 2272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1713453518
transform 1 0 2224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1713453518
transform 1 0 2216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1713453518
transform 1 0 2208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1713453518
transform 1 0 2200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1713453518
transform 1 0 2160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1713453518
transform 1 0 2152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3841
timestamp 1713453518
transform 1 0 2144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1713453518
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1713453518
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1713453518
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1713453518
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1713453518
transform 1 0 2040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1713453518
transform 1 0 2032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1713453518
transform 1 0 2024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1713453518
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1713453518
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1713453518
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1713453518
transform 1 0 1952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1713453518
transform 1 0 1944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1713453518
transform 1 0 1936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1713453518
transform 1 0 1896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1713453518
transform 1 0 1864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3857
timestamp 1713453518
transform 1 0 1856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1713453518
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1713453518
transform 1 0 1800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1713453518
transform 1 0 1792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1713453518
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1713453518
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1713453518
transform 1 0 1768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1713453518
transform 1 0 1760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1713453518
transform 1 0 1720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1713453518
transform 1 0 1712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1713453518
transform 1 0 1704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1713453518
transform 1 0 1696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1713453518
transform 1 0 1648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1713453518
transform 1 0 1640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1713453518
transform 1 0 1632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1713453518
transform 1 0 1624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1713453518
transform 1 0 1592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1713453518
transform 1 0 1568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1713453518
transform 1 0 1560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1713453518
transform 1 0 1552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1713453518
transform 1 0 1544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1713453518
transform 1 0 1504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1713453518
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3880
timestamp 1713453518
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1713453518
transform 1 0 1424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1713453518
transform 1 0 1416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1713453518
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1713453518
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1713453518
transform 1 0 1392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1713453518
transform 1 0 1344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1713453518
transform 1 0 1336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1713453518
transform 1 0 1328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1713453518
transform 1 0 1320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1713453518
transform 1 0 1272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1713453518
transform 1 0 1264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1713453518
transform 1 0 1256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1713453518
transform 1 0 1248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1713453518
transform 1 0 1240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1713453518
transform 1 0 1232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1713453518
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1713453518
transform 1 0 1176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1713453518
transform 1 0 1168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1713453518
transform 1 0 1128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1713453518
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1713453518
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1713453518
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1713453518
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1713453518
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1713453518
transform 1 0 1016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1713453518
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1713453518
transform 1 0 904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1713453518
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1713453518
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1713453518
transform 1 0 816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1713453518
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1713453518
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1713453518
transform 1 0 704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1713453518
transform 1 0 680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1713453518
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1713453518
transform 1 0 600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1713453518
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1713453518
transform 1 0 584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1713453518
transform 1 0 496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1713453518
transform 1 0 488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1713453518
transform 1 0 480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1713453518
transform 1 0 392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1713453518
transform 1 0 384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1713453518
transform 1 0 376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1713453518
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3926
timestamp 1713453518
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1713453518
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1713453518
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1713453518
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1713453518
transform 1 0 3440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1713453518
transform 1 0 3432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1713453518
transform 1 0 3424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1713453518
transform 1 0 3416 0 1 1170
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1713453518
transform 1 0 3376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1713453518
transform 1 0 3368 0 1 1170
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1713453518
transform 1 0 3360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1713453518
transform 1 0 3352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1713453518
transform 1 0 3312 0 1 1170
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1713453518
transform 1 0 3304 0 1 1170
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1713453518
transform 1 0 3296 0 1 1170
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1713453518
transform 1 0 3264 0 1 1170
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1713453518
transform 1 0 3256 0 1 1170
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1713453518
transform 1 0 3248 0 1 1170
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1713453518
transform 1 0 3240 0 1 1170
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1713453518
transform 1 0 3232 0 1 1170
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1713453518
transform 1 0 3200 0 1 1170
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1713453518
transform 1 0 3192 0 1 1170
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1713453518
transform 1 0 3184 0 1 1170
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1713453518
transform 1 0 3176 0 1 1170
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1713453518
transform 1 0 3168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1713453518
transform 1 0 3128 0 1 1170
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1713453518
transform 1 0 3120 0 1 1170
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1713453518
transform 1 0 3112 0 1 1170
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1713453518
transform 1 0 3104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1713453518
transform 1 0 3080 0 1 1170
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1713453518
transform 1 0 3072 0 1 1170
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1713453518
transform 1 0 3064 0 1 1170
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1713453518
transform 1 0 3032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1713453518
transform 1 0 3024 0 1 1170
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1713453518
transform 1 0 3016 0 1 1170
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1713453518
transform 1 0 3008 0 1 1170
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1713453518
transform 1 0 2968 0 1 1170
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1713453518
transform 1 0 2960 0 1 1170
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1713453518
transform 1 0 2952 0 1 1170
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1713453518
transform 1 0 2944 0 1 1170
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1713453518
transform 1 0 2936 0 1 1170
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1713453518
transform 1 0 2904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1713453518
transform 1 0 2896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1713453518
transform 1 0 2888 0 1 1170
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1713453518
transform 1 0 2880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1713453518
transform 1 0 2848 0 1 1170
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1713453518
transform 1 0 2840 0 1 1170
box -8 -3 16 105
use FILL  FILL_3973
timestamp 1713453518
transform 1 0 2832 0 1 1170
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1713453518
transform 1 0 2808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1713453518
transform 1 0 2800 0 1 1170
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1713453518
transform 1 0 2792 0 1 1170
box -8 -3 16 105
use FILL  FILL_3977
timestamp 1713453518
transform 1 0 2744 0 1 1170
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1713453518
transform 1 0 2736 0 1 1170
box -8 -3 16 105
use FILL  FILL_3979
timestamp 1713453518
transform 1 0 2728 0 1 1170
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1713453518
transform 1 0 2720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1713453518
transform 1 0 2712 0 1 1170
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1713453518
transform 1 0 2704 0 1 1170
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1713453518
transform 1 0 2696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1713453518
transform 1 0 2632 0 1 1170
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1713453518
transform 1 0 2624 0 1 1170
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1713453518
transform 1 0 2616 0 1 1170
box -8 -3 16 105
use FILL  FILL_3987
timestamp 1713453518
transform 1 0 2608 0 1 1170
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1713453518
transform 1 0 2600 0 1 1170
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1713453518
transform 1 0 2560 0 1 1170
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1713453518
transform 1 0 2552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1713453518
transform 1 0 2544 0 1 1170
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1713453518
transform 1 0 2504 0 1 1170
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1713453518
transform 1 0 2496 0 1 1170
box -8 -3 16 105
use FILL  FILL_3994
timestamp 1713453518
transform 1 0 2488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1713453518
transform 1 0 2480 0 1 1170
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1713453518
transform 1 0 2440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3997
timestamp 1713453518
transform 1 0 2432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1713453518
transform 1 0 2424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1713453518
transform 1 0 2384 0 1 1170
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1713453518
transform 1 0 2376 0 1 1170
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1713453518
transform 1 0 2368 0 1 1170
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1713453518
transform 1 0 2360 0 1 1170
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1713453518
transform 1 0 2352 0 1 1170
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1713453518
transform 1 0 2304 0 1 1170
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1713453518
transform 1 0 2296 0 1 1170
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1713453518
transform 1 0 2288 0 1 1170
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1713453518
transform 1 0 2280 0 1 1170
box -8 -3 16 105
use FILL  FILL_4008
timestamp 1713453518
transform 1 0 2248 0 1 1170
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1713453518
transform 1 0 2240 0 1 1170
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1713453518
transform 1 0 2232 0 1 1170
box -8 -3 16 105
use FILL  FILL_4011
timestamp 1713453518
transform 1 0 2192 0 1 1170
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1713453518
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1713453518
transform 1 0 2176 0 1 1170
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1713453518
transform 1 0 2152 0 1 1170
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1713453518
transform 1 0 2144 0 1 1170
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1713453518
transform 1 0 2136 0 1 1170
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1713453518
transform 1 0 2128 0 1 1170
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1713453518
transform 1 0 2080 0 1 1170
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1713453518
transform 1 0 2072 0 1 1170
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1713453518
transform 1 0 2064 0 1 1170
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1713453518
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1713453518
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1713453518
transform 1 0 2008 0 1 1170
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1713453518
transform 1 0 2000 0 1 1170
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1713453518
transform 1 0 1992 0 1 1170
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1713453518
transform 1 0 1984 0 1 1170
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1713453518
transform 1 0 1976 0 1 1170
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1713453518
transform 1 0 1928 0 1 1170
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1713453518
transform 1 0 1920 0 1 1170
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1713453518
transform 1 0 1912 0 1 1170
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1713453518
transform 1 0 1872 0 1 1170
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1713453518
transform 1 0 1864 0 1 1170
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1713453518
transform 1 0 1856 0 1 1170
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1713453518
transform 1 0 1848 0 1 1170
box -8 -3 16 105
use FILL  FILL_4035
timestamp 1713453518
transform 1 0 1816 0 1 1170
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1713453518
transform 1 0 1808 0 1 1170
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1713453518
transform 1 0 1800 0 1 1170
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1713453518
transform 1 0 1760 0 1 1170
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1713453518
transform 1 0 1752 0 1 1170
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1713453518
transform 1 0 1744 0 1 1170
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1713453518
transform 1 0 1736 0 1 1170
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1713453518
transform 1 0 1728 0 1 1170
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1713453518
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1713453518
transform 1 0 1688 0 1 1170
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1713453518
transform 1 0 1680 0 1 1170
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1713453518
transform 1 0 1672 0 1 1170
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1713453518
transform 1 0 1632 0 1 1170
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1713453518
transform 1 0 1624 0 1 1170
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1713453518
transform 1 0 1616 0 1 1170
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1713453518
transform 1 0 1608 0 1 1170
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1713453518
transform 1 0 1600 0 1 1170
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1713453518
transform 1 0 1544 0 1 1170
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1713453518
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1713453518
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1713453518
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1713453518
transform 1 0 1480 0 1 1170
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1713453518
transform 1 0 1472 0 1 1170
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1713453518
transform 1 0 1464 0 1 1170
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1713453518
transform 1 0 1432 0 1 1170
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1713453518
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1713453518
transform 1 0 1416 0 1 1170
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1713453518
transform 1 0 1408 0 1 1170
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1713453518
transform 1 0 1376 0 1 1170
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1713453518
transform 1 0 1352 0 1 1170
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1713453518
transform 1 0 1344 0 1 1170
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1713453518
transform 1 0 1336 0 1 1170
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1713453518
transform 1 0 1328 0 1 1170
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1713453518
transform 1 0 1280 0 1 1170
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1713453518
transform 1 0 1272 0 1 1170
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1713453518
transform 1 0 1264 0 1 1170
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1713453518
transform 1 0 1256 0 1 1170
box -8 -3 16 105
use FILL  FILL_4072
timestamp 1713453518
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1713453518
transform 1 0 1208 0 1 1170
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1713453518
transform 1 0 1200 0 1 1170
box -8 -3 16 105
use FILL  FILL_4075
timestamp 1713453518
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1713453518
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1713453518
transform 1 0 1136 0 1 1170
box -8 -3 16 105
use FILL  FILL_4078
timestamp 1713453518
transform 1 0 1128 0 1 1170
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1713453518
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1713453518
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1713453518
transform 1 0 1104 0 1 1170
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1713453518
transform 1 0 1048 0 1 1170
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1713453518
transform 1 0 1040 0 1 1170
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1713453518
transform 1 0 1032 0 1 1170
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1713453518
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1713453518
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1713453518
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1713453518
transform 1 0 808 0 1 1170
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1713453518
transform 1 0 800 0 1 1170
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1713453518
transform 1 0 792 0 1 1170
box -8 -3 16 105
use FILL  FILL_4091
timestamp 1713453518
transform 1 0 696 0 1 1170
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1713453518
transform 1 0 688 0 1 1170
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1713453518
transform 1 0 680 0 1 1170
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1713453518
transform 1 0 672 0 1 1170
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1713453518
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1713453518
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1713453518
transform 1 0 592 0 1 1170
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1713453518
transform 1 0 584 0 1 1170
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1713453518
transform 1 0 576 0 1 1170
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1713453518
transform 1 0 528 0 1 1170
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1713453518
transform 1 0 520 0 1 1170
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1713453518
transform 1 0 512 0 1 1170
box -8 -3 16 105
use FILL  FILL_4103
timestamp 1713453518
transform 1 0 504 0 1 1170
box -8 -3 16 105
use FILL  FILL_4104
timestamp 1713453518
transform 1 0 440 0 1 1170
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1713453518
transform 1 0 432 0 1 1170
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1713453518
transform 1 0 424 0 1 1170
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1713453518
transform 1 0 416 0 1 1170
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1713453518
transform 1 0 312 0 1 1170
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1713453518
transform 1 0 304 0 1 1170
box -8 -3 16 105
use FILL  FILL_4110
timestamp 1713453518
transform 1 0 296 0 1 1170
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1713453518
transform 1 0 288 0 1 1170
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1713453518
transform 1 0 208 0 1 1170
box -8 -3 16 105
use FILL  FILL_4113
timestamp 1713453518
transform 1 0 200 0 1 1170
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1713453518
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1713453518
transform 1 0 184 0 1 1170
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1713453518
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1713453518
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1713453518
transform 1 0 3440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1713453518
transform 1 0 3432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1713453518
transform 1 0 3424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1713453518
transform 1 0 3376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4122
timestamp 1713453518
transform 1 0 3368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1713453518
transform 1 0 3360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1713453518
transform 1 0 3352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1713453518
transform 1 0 3344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1713453518
transform 1 0 3312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1713453518
transform 1 0 3304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1713453518
transform 1 0 3264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1713453518
transform 1 0 3256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1713453518
transform 1 0 3248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1713453518
transform 1 0 3240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1713453518
transform 1 0 3232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1713453518
transform 1 0 3224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1713453518
transform 1 0 3216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1713453518
transform 1 0 3176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1713453518
transform 1 0 3168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1713453518
transform 1 0 3160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4138
timestamp 1713453518
transform 1 0 3128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1713453518
transform 1 0 3120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1713453518
transform 1 0 3112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1713453518
transform 1 0 3104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1713453518
transform 1 0 3096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1713453518
transform 1 0 3088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1713453518
transform 1 0 3040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1713453518
transform 1 0 3032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1713453518
transform 1 0 3024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1713453518
transform 1 0 3016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1713453518
transform 1 0 3008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1713453518
transform 1 0 2960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1713453518
transform 1 0 2952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1713453518
transform 1 0 2944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1713453518
transform 1 0 2936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1713453518
transform 1 0 2928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4154
timestamp 1713453518
transform 1 0 2904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1713453518
transform 1 0 2856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1713453518
transform 1 0 2848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1713453518
transform 1 0 2840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1713453518
transform 1 0 2832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1713453518
transform 1 0 2824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1713453518
transform 1 0 2792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1713453518
transform 1 0 2760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1713453518
transform 1 0 2752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1713453518
transform 1 0 2744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1713453518
transform 1 0 2736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4165
timestamp 1713453518
transform 1 0 2728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1713453518
transform 1 0 2680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1713453518
transform 1 0 2672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1713453518
transform 1 0 2664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1713453518
transform 1 0 2640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1713453518
transform 1 0 2632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1713453518
transform 1 0 2608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1713453518
transform 1 0 2600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1713453518
transform 1 0 2552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1713453518
transform 1 0 2544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1713453518
transform 1 0 2536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1713453518
transform 1 0 2528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4177
timestamp 1713453518
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1713453518
transform 1 0 2472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1713453518
transform 1 0 2464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1713453518
transform 1 0 2456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1713453518
transform 1 0 2416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1713453518
transform 1 0 2408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1713453518
transform 1 0 2376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1713453518
transform 1 0 2368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1713453518
transform 1 0 2320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4186
timestamp 1713453518
transform 1 0 2312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1713453518
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1713453518
transform 1 0 2296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1713453518
transform 1 0 2288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1713453518
transform 1 0 2224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1713453518
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4192
timestamp 1713453518
transform 1 0 2208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1713453518
transform 1 0 2200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1713453518
transform 1 0 2152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1713453518
transform 1 0 2144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1713453518
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1713453518
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1713453518
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4199
timestamp 1713453518
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1713453518
transform 1 0 2056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1713453518
transform 1 0 2048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1713453518
transform 1 0 2008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1713453518
transform 1 0 2000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1713453518
transform 1 0 1992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1713453518
transform 1 0 1952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1713453518
transform 1 0 1912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1713453518
transform 1 0 1904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1713453518
transform 1 0 1896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1713453518
transform 1 0 1848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1713453518
transform 1 0 1840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4211
timestamp 1713453518
transform 1 0 1832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1713453518
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1713453518
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1713453518
transform 1 0 1776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1713453518
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1713453518
transform 1 0 1712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1713453518
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1713453518
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1713453518
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1713453518
transform 1 0 1632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4221
timestamp 1713453518
transform 1 0 1624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1713453518
transform 1 0 1616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1713453518
transform 1 0 1592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1713453518
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1713453518
transform 1 0 1544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4226
timestamp 1713453518
transform 1 0 1536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1713453518
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1713453518
transform 1 0 1480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1713453518
transform 1 0 1472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1713453518
transform 1 0 1424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1713453518
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4232
timestamp 1713453518
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1713453518
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1713453518
transform 1 0 1392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1713453518
transform 1 0 1336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1713453518
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1713453518
transform 1 0 1320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1713453518
transform 1 0 1312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1713453518
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1713453518
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1713453518
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1713453518
transform 1 0 1224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1713453518
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4244
timestamp 1713453518
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1713453518
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1713453518
transform 1 0 1144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1713453518
transform 1 0 1136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1713453518
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1713453518
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1713453518
transform 1 0 1048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1713453518
transform 1 0 1040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1713453518
transform 1 0 1032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1713453518
transform 1 0 1024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1713453518
transform 1 0 952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1713453518
transform 1 0 944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1713453518
transform 1 0 936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1713453518
transform 1 0 832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1713453518
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1713453518
transform 1 0 816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4260
timestamp 1713453518
transform 1 0 688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4261
timestamp 1713453518
transform 1 0 680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1713453518
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4263
timestamp 1713453518
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4264
timestamp 1713453518
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1713453518
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4266
timestamp 1713453518
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4267
timestamp 1713453518
transform 1 0 512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1713453518
transform 1 0 440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1713453518
transform 1 0 432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1713453518
transform 1 0 424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4271
timestamp 1713453518
transform 1 0 376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4272
timestamp 1713453518
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4273
timestamp 1713453518
transform 1 0 304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1713453518
transform 1 0 296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1713453518
transform 1 0 192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1713453518
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4277
timestamp 1713453518
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1713453518
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1713453518
transform 1 0 3440 0 1 970
box -8 -3 16 105
use FILL  FILL_4280
timestamp 1713453518
transform 1 0 3432 0 1 970
box -8 -3 16 105
use FILL  FILL_4281
timestamp 1713453518
transform 1 0 3424 0 1 970
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1713453518
transform 1 0 3360 0 1 970
box -8 -3 16 105
use FILL  FILL_4283
timestamp 1713453518
transform 1 0 3352 0 1 970
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1713453518
transform 1 0 3344 0 1 970
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1713453518
transform 1 0 3336 0 1 970
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1713453518
transform 1 0 3296 0 1 970
box -8 -3 16 105
use FILL  FILL_4287
timestamp 1713453518
transform 1 0 3256 0 1 970
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1713453518
transform 1 0 3248 0 1 970
box -8 -3 16 105
use FILL  FILL_4289
timestamp 1713453518
transform 1 0 3240 0 1 970
box -8 -3 16 105
use FILL  FILL_4290
timestamp 1713453518
transform 1 0 3232 0 1 970
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1713453518
transform 1 0 3224 0 1 970
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1713453518
transform 1 0 3216 0 1 970
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1713453518
transform 1 0 3176 0 1 970
box -8 -3 16 105
use FILL  FILL_4294
timestamp 1713453518
transform 1 0 3168 0 1 970
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1713453518
transform 1 0 3136 0 1 970
box -8 -3 16 105
use FILL  FILL_4296
timestamp 1713453518
transform 1 0 3128 0 1 970
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1713453518
transform 1 0 3120 0 1 970
box -8 -3 16 105
use FILL  FILL_4298
timestamp 1713453518
transform 1 0 3112 0 1 970
box -8 -3 16 105
use FILL  FILL_4299
timestamp 1713453518
transform 1 0 3104 0 1 970
box -8 -3 16 105
use FILL  FILL_4300
timestamp 1713453518
transform 1 0 3096 0 1 970
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1713453518
transform 1 0 3056 0 1 970
box -8 -3 16 105
use FILL  FILL_4302
timestamp 1713453518
transform 1 0 3048 0 1 970
box -8 -3 16 105
use FILL  FILL_4303
timestamp 1713453518
transform 1 0 3016 0 1 970
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1713453518
transform 1 0 3008 0 1 970
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1713453518
transform 1 0 3000 0 1 970
box -8 -3 16 105
use FILL  FILL_4306
timestamp 1713453518
transform 1 0 2992 0 1 970
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1713453518
transform 1 0 2984 0 1 970
box -8 -3 16 105
use FILL  FILL_4308
timestamp 1713453518
transform 1 0 2976 0 1 970
box -8 -3 16 105
use FILL  FILL_4309
timestamp 1713453518
transform 1 0 2912 0 1 970
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1713453518
transform 1 0 2904 0 1 970
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1713453518
transform 1 0 2896 0 1 970
box -8 -3 16 105
use FILL  FILL_4312
timestamp 1713453518
transform 1 0 2888 0 1 970
box -8 -3 16 105
use FILL  FILL_4313
timestamp 1713453518
transform 1 0 2880 0 1 970
box -8 -3 16 105
use FILL  FILL_4314
timestamp 1713453518
transform 1 0 2872 0 1 970
box -8 -3 16 105
use FILL  FILL_4315
timestamp 1713453518
transform 1 0 2832 0 1 970
box -8 -3 16 105
use FILL  FILL_4316
timestamp 1713453518
transform 1 0 2800 0 1 970
box -8 -3 16 105
use FILL  FILL_4317
timestamp 1713453518
transform 1 0 2792 0 1 970
box -8 -3 16 105
use FILL  FILL_4318
timestamp 1713453518
transform 1 0 2768 0 1 970
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1713453518
transform 1 0 2760 0 1 970
box -8 -3 16 105
use FILL  FILL_4320
timestamp 1713453518
transform 1 0 2752 0 1 970
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1713453518
transform 1 0 2688 0 1 970
box -8 -3 16 105
use FILL  FILL_4322
timestamp 1713453518
transform 1 0 2680 0 1 970
box -8 -3 16 105
use FILL  FILL_4323
timestamp 1713453518
transform 1 0 2672 0 1 970
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1713453518
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_4325
timestamp 1713453518
transform 1 0 2656 0 1 970
box -8 -3 16 105
use FILL  FILL_4326
timestamp 1713453518
transform 1 0 2584 0 1 970
box -8 -3 16 105
use FILL  FILL_4327
timestamp 1713453518
transform 1 0 2576 0 1 970
box -8 -3 16 105
use FILL  FILL_4328
timestamp 1713453518
transform 1 0 2568 0 1 970
box -8 -3 16 105
use FILL  FILL_4329
timestamp 1713453518
transform 1 0 2560 0 1 970
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1713453518
transform 1 0 2552 0 1 970
box -8 -3 16 105
use FILL  FILL_4331
timestamp 1713453518
transform 1 0 2472 0 1 970
box -8 -3 16 105
use FILL  FILL_4332
timestamp 1713453518
transform 1 0 2464 0 1 970
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1713453518
transform 1 0 2456 0 1 970
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1713453518
transform 1 0 2448 0 1 970
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1713453518
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_4336
timestamp 1713453518
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_4337
timestamp 1713453518
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_4338
timestamp 1713453518
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_4339
timestamp 1713453518
transform 1 0 2328 0 1 970
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1713453518
transform 1 0 2320 0 1 970
box -8 -3 16 105
use FILL  FILL_4341
timestamp 1713453518
transform 1 0 2248 0 1 970
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1713453518
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1713453518
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1713453518
transform 1 0 2224 0 1 970
box -8 -3 16 105
use FILL  FILL_4345
timestamp 1713453518
transform 1 0 2216 0 1 970
box -8 -3 16 105
use FILL  FILL_4346
timestamp 1713453518
transform 1 0 2152 0 1 970
box -8 -3 16 105
use FILL  FILL_4347
timestamp 1713453518
transform 1 0 2144 0 1 970
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1713453518
transform 1 0 2136 0 1 970
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1713453518
transform 1 0 2128 0 1 970
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1713453518
transform 1 0 2120 0 1 970
box -8 -3 16 105
use FILL  FILL_4351
timestamp 1713453518
transform 1 0 2056 0 1 970
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1713453518
transform 1 0 2048 0 1 970
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1713453518
transform 1 0 2040 0 1 970
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1713453518
transform 1 0 2032 0 1 970
box -8 -3 16 105
use FILL  FILL_4355
timestamp 1713453518
transform 1 0 1968 0 1 970
box -8 -3 16 105
use FILL  FILL_4356
timestamp 1713453518
transform 1 0 1960 0 1 970
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1713453518
transform 1 0 1952 0 1 970
box -8 -3 16 105
use FILL  FILL_4358
timestamp 1713453518
transform 1 0 1944 0 1 970
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1713453518
transform 1 0 1904 0 1 970
box -8 -3 16 105
use FILL  FILL_4360
timestamp 1713453518
transform 1 0 1864 0 1 970
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1713453518
transform 1 0 1856 0 1 970
box -8 -3 16 105
use FILL  FILL_4362
timestamp 1713453518
transform 1 0 1848 0 1 970
box -8 -3 16 105
use FILL  FILL_4363
timestamp 1713453518
transform 1 0 1840 0 1 970
box -8 -3 16 105
use FILL  FILL_4364
timestamp 1713453518
transform 1 0 1832 0 1 970
box -8 -3 16 105
use FILL  FILL_4365
timestamp 1713453518
transform 1 0 1760 0 1 970
box -8 -3 16 105
use FILL  FILL_4366
timestamp 1713453518
transform 1 0 1752 0 1 970
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1713453518
transform 1 0 1744 0 1 970
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1713453518
transform 1 0 1704 0 1 970
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1713453518
transform 1 0 1696 0 1 970
box -8 -3 16 105
use FILL  FILL_4370
timestamp 1713453518
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_4371
timestamp 1713453518
transform 1 0 1632 0 1 970
box -8 -3 16 105
use FILL  FILL_4372
timestamp 1713453518
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1713453518
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1713453518
transform 1 0 1608 0 1 970
box -8 -3 16 105
use FILL  FILL_4375
timestamp 1713453518
transform 1 0 1600 0 1 970
box -8 -3 16 105
use FILL  FILL_4376
timestamp 1713453518
transform 1 0 1536 0 1 970
box -8 -3 16 105
use FILL  FILL_4377
timestamp 1713453518
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_4378
timestamp 1713453518
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_4379
timestamp 1713453518
transform 1 0 1512 0 1 970
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1713453518
transform 1 0 1504 0 1 970
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1713453518
transform 1 0 1424 0 1 970
box -8 -3 16 105
use FILL  FILL_4382
timestamp 1713453518
transform 1 0 1416 0 1 970
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1713453518
transform 1 0 1408 0 1 970
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1713453518
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_4385
timestamp 1713453518
transform 1 0 1392 0 1 970
box -8 -3 16 105
use FILL  FILL_4386
timestamp 1713453518
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1713453518
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1713453518
transform 1 0 1304 0 1 970
box -8 -3 16 105
use FILL  FILL_4389
timestamp 1713453518
transform 1 0 1296 0 1 970
box -8 -3 16 105
use FILL  FILL_4390
timestamp 1713453518
transform 1 0 1256 0 1 970
box -8 -3 16 105
use FILL  FILL_4391
timestamp 1713453518
transform 1 0 1248 0 1 970
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1713453518
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_4393
timestamp 1713453518
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_4394
timestamp 1713453518
transform 1 0 1192 0 1 970
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1713453518
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_4396
timestamp 1713453518
transform 1 0 1120 0 1 970
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1713453518
transform 1 0 1112 0 1 970
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1713453518
transform 1 0 1088 0 1 970
box -8 -3 16 105
use FILL  FILL_4399
timestamp 1713453518
transform 1 0 1048 0 1 970
box -8 -3 16 105
use FILL  FILL_4400
timestamp 1713453518
transform 1 0 1040 0 1 970
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1713453518
transform 1 0 1032 0 1 970
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1713453518
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_4403
timestamp 1713453518
transform 1 0 952 0 1 970
box -8 -3 16 105
use FILL  FILL_4404
timestamp 1713453518
transform 1 0 944 0 1 970
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1713453518
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_4406
timestamp 1713453518
transform 1 0 832 0 1 970
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1713453518
transform 1 0 824 0 1 970
box -8 -3 16 105
use FILL  FILL_4408
timestamp 1713453518
transform 1 0 816 0 1 970
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1713453518
transform 1 0 808 0 1 970
box -8 -3 16 105
use FILL  FILL_4410
timestamp 1713453518
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_4411
timestamp 1713453518
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_4412
timestamp 1713453518
transform 1 0 712 0 1 970
box -8 -3 16 105
use FILL  FILL_4413
timestamp 1713453518
transform 1 0 704 0 1 970
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1713453518
transform 1 0 640 0 1 970
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1713453518
transform 1 0 632 0 1 970
box -8 -3 16 105
use FILL  FILL_4416
timestamp 1713453518
transform 1 0 624 0 1 970
box -8 -3 16 105
use FILL  FILL_4417
timestamp 1713453518
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1713453518
transform 1 0 568 0 1 970
box -8 -3 16 105
use FILL  FILL_4419
timestamp 1713453518
transform 1 0 512 0 1 970
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1713453518
transform 1 0 504 0 1 970
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1713453518
transform 1 0 496 0 1 970
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1713453518
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_4423
timestamp 1713453518
transform 1 0 408 0 1 970
box -8 -3 16 105
use FILL  FILL_4424
timestamp 1713453518
transform 1 0 400 0 1 970
box -8 -3 16 105
use FILL  FILL_4425
timestamp 1713453518
transform 1 0 392 0 1 970
box -8 -3 16 105
use FILL  FILL_4426
timestamp 1713453518
transform 1 0 384 0 1 970
box -8 -3 16 105
use FILL  FILL_4427
timestamp 1713453518
transform 1 0 296 0 1 970
box -8 -3 16 105
use FILL  FILL_4428
timestamp 1713453518
transform 1 0 288 0 1 970
box -8 -3 16 105
use FILL  FILL_4429
timestamp 1713453518
transform 1 0 280 0 1 970
box -8 -3 16 105
use FILL  FILL_4430
timestamp 1713453518
transform 1 0 200 0 1 970
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1713453518
transform 1 0 192 0 1 970
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1713453518
transform 1 0 184 0 1 970
box -8 -3 16 105
use FILL  FILL_4433
timestamp 1713453518
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1713453518
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_4435
timestamp 1713453518
transform 1 0 88 0 1 970
box -8 -3 16 105
use FILL  FILL_4436
timestamp 1713453518
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_4437
timestamp 1713453518
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1713453518
transform 1 0 3440 0 -1 970
box -8 -3 16 105
use FILL  FILL_4439
timestamp 1713453518
transform 1 0 3432 0 -1 970
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1713453518
transform 1 0 3392 0 -1 970
box -8 -3 16 105
use FILL  FILL_4441
timestamp 1713453518
transform 1 0 3384 0 -1 970
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1713453518
transform 1 0 3376 0 -1 970
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1713453518
transform 1 0 3328 0 -1 970
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1713453518
transform 1 0 3320 0 -1 970
box -8 -3 16 105
use FILL  FILL_4445
timestamp 1713453518
transform 1 0 3312 0 -1 970
box -8 -3 16 105
use FILL  FILL_4446
timestamp 1713453518
transform 1 0 3304 0 -1 970
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1713453518
transform 1 0 3248 0 -1 970
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1713453518
transform 1 0 3240 0 -1 970
box -8 -3 16 105
use FILL  FILL_4449
timestamp 1713453518
transform 1 0 3232 0 -1 970
box -8 -3 16 105
use FILL  FILL_4450
timestamp 1713453518
transform 1 0 3200 0 -1 970
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1713453518
transform 1 0 3192 0 -1 970
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1713453518
transform 1 0 3184 0 -1 970
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1713453518
transform 1 0 3152 0 -1 970
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1713453518
transform 1 0 3144 0 -1 970
box -8 -3 16 105
use FILL  FILL_4455
timestamp 1713453518
transform 1 0 3112 0 -1 970
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1713453518
transform 1 0 3104 0 -1 970
box -8 -3 16 105
use FILL  FILL_4457
timestamp 1713453518
transform 1 0 3096 0 -1 970
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1713453518
transform 1 0 3088 0 -1 970
box -8 -3 16 105
use FILL  FILL_4459
timestamp 1713453518
transform 1 0 3080 0 -1 970
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1713453518
transform 1 0 3072 0 -1 970
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1713453518
transform 1 0 3016 0 -1 970
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1713453518
transform 1 0 3008 0 -1 970
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1713453518
transform 1 0 2968 0 -1 970
box -8 -3 16 105
use FILL  FILL_4464
timestamp 1713453518
transform 1 0 2960 0 -1 970
box -8 -3 16 105
use FILL  FILL_4465
timestamp 1713453518
transform 1 0 2952 0 -1 970
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1713453518
transform 1 0 2944 0 -1 970
box -8 -3 16 105
use FILL  FILL_4467
timestamp 1713453518
transform 1 0 2936 0 -1 970
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1713453518
transform 1 0 2872 0 -1 970
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1713453518
transform 1 0 2864 0 -1 970
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1713453518
transform 1 0 2856 0 -1 970
box -8 -3 16 105
use FILL  FILL_4471
timestamp 1713453518
transform 1 0 2848 0 -1 970
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1713453518
transform 1 0 2840 0 -1 970
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1713453518
transform 1 0 2768 0 -1 970
box -8 -3 16 105
use FILL  FILL_4474
timestamp 1713453518
transform 1 0 2760 0 -1 970
box -8 -3 16 105
use FILL  FILL_4475
timestamp 1713453518
transform 1 0 2752 0 -1 970
box -8 -3 16 105
use FILL  FILL_4476
timestamp 1713453518
transform 1 0 2744 0 -1 970
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1713453518
transform 1 0 2736 0 -1 970
box -8 -3 16 105
use FILL  FILL_4478
timestamp 1713453518
transform 1 0 2728 0 -1 970
box -8 -3 16 105
use FILL  FILL_4479
timestamp 1713453518
transform 1 0 2664 0 -1 970
box -8 -3 16 105
use FILL  FILL_4480
timestamp 1713453518
transform 1 0 2656 0 -1 970
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1713453518
transform 1 0 2648 0 -1 970
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1713453518
transform 1 0 2608 0 -1 970
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1713453518
transform 1 0 2600 0 -1 970
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1713453518
transform 1 0 2528 0 -1 970
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1713453518
transform 1 0 2520 0 -1 970
box -8 -3 16 105
use FILL  FILL_4486
timestamp 1713453518
transform 1 0 2512 0 -1 970
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1713453518
transform 1 0 2504 0 -1 970
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1713453518
transform 1 0 2496 0 -1 970
box -8 -3 16 105
use FILL  FILL_4489
timestamp 1713453518
transform 1 0 2432 0 -1 970
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1713453518
transform 1 0 2384 0 -1 970
box -8 -3 16 105
use FILL  FILL_4491
timestamp 1713453518
transform 1 0 2376 0 -1 970
box -8 -3 16 105
use FILL  FILL_4492
timestamp 1713453518
transform 1 0 2368 0 -1 970
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1713453518
transform 1 0 2360 0 -1 970
box -8 -3 16 105
use FILL  FILL_4494
timestamp 1713453518
transform 1 0 2288 0 -1 970
box -8 -3 16 105
use FILL  FILL_4495
timestamp 1713453518
transform 1 0 2280 0 -1 970
box -8 -3 16 105
use FILL  FILL_4496
timestamp 1713453518
transform 1 0 2256 0 -1 970
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1713453518
transform 1 0 2248 0 -1 970
box -8 -3 16 105
use FILL  FILL_4498
timestamp 1713453518
transform 1 0 2200 0 -1 970
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1713453518
transform 1 0 2144 0 -1 970
box -8 -3 16 105
use FILL  FILL_4500
timestamp 1713453518
transform 1 0 2136 0 -1 970
box -8 -3 16 105
use FILL  FILL_4501
timestamp 1713453518
transform 1 0 2096 0 -1 970
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1713453518
transform 1 0 2088 0 -1 970
box -8 -3 16 105
use FILL  FILL_4503
timestamp 1713453518
transform 1 0 2040 0 -1 970
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1713453518
transform 1 0 2008 0 -1 970
box -8 -3 16 105
use FILL  FILL_4505
timestamp 1713453518
transform 1 0 2000 0 -1 970
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1713453518
transform 1 0 1992 0 -1 970
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1713453518
transform 1 0 1936 0 -1 970
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1713453518
transform 1 0 1928 0 -1 970
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1713453518
transform 1 0 1920 0 -1 970
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1713453518
transform 1 0 1856 0 -1 970
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1713453518
transform 1 0 1848 0 -1 970
box -8 -3 16 105
use FILL  FILL_4512
timestamp 1713453518
transform 1 0 1808 0 -1 970
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1713453518
transform 1 0 1800 0 -1 970
box -8 -3 16 105
use FILL  FILL_4514
timestamp 1713453518
transform 1 0 1752 0 -1 970
box -8 -3 16 105
use FILL  FILL_4515
timestamp 1713453518
transform 1 0 1744 0 -1 970
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1713453518
transform 1 0 1736 0 -1 970
box -8 -3 16 105
use FILL  FILL_4517
timestamp 1713453518
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_4518
timestamp 1713453518
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_4519
timestamp 1713453518
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1713453518
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1713453518
transform 1 0 1616 0 -1 970
box -8 -3 16 105
use FILL  FILL_4522
timestamp 1713453518
transform 1 0 1592 0 -1 970
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1713453518
transform 1 0 1584 0 -1 970
box -8 -3 16 105
use FILL  FILL_4524
timestamp 1713453518
transform 1 0 1576 0 -1 970
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1713453518
transform 1 0 1528 0 -1 970
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1713453518
transform 1 0 1488 0 -1 970
box -8 -3 16 105
use FILL  FILL_4527
timestamp 1713453518
transform 1 0 1480 0 -1 970
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1713453518
transform 1 0 1472 0 -1 970
box -8 -3 16 105
use FILL  FILL_4529
timestamp 1713453518
transform 1 0 1400 0 -1 970
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1713453518
transform 1 0 1392 0 -1 970
box -8 -3 16 105
use FILL  FILL_4531
timestamp 1713453518
transform 1 0 1368 0 -1 970
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1713453518
transform 1 0 1360 0 -1 970
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1713453518
transform 1 0 1328 0 -1 970
box -8 -3 16 105
use FILL  FILL_4534
timestamp 1713453518
transform 1 0 1296 0 -1 970
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1713453518
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use FILL  FILL_4536
timestamp 1713453518
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use FILL  FILL_4537
timestamp 1713453518
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use FILL  FILL_4538
timestamp 1713453518
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1713453518
transform 1 0 1184 0 -1 970
box -8 -3 16 105
use FILL  FILL_4540
timestamp 1713453518
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1713453518
transform 1 0 1168 0 -1 970
box -8 -3 16 105
use FILL  FILL_4542
timestamp 1713453518
transform 1 0 1088 0 -1 970
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1713453518
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1713453518
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1713453518
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1713453518
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1713453518
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1713453518
transform 1 0 976 0 -1 970
box -8 -3 16 105
use FILL  FILL_4549
timestamp 1713453518
transform 1 0 968 0 -1 970
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1713453518
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_4551
timestamp 1713453518
transform 1 0 952 0 -1 970
box -8 -3 16 105
use FILL  FILL_4552
timestamp 1713453518
transform 1 0 928 0 -1 970
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1713453518
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1713453518
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_4555
timestamp 1713453518
transform 1 0 848 0 -1 970
box -8 -3 16 105
use FILL  FILL_4556
timestamp 1713453518
transform 1 0 840 0 -1 970
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1713453518
transform 1 0 832 0 -1 970
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1713453518
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_4559
timestamp 1713453518
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_4560
timestamp 1713453518
transform 1 0 808 0 -1 970
box -8 -3 16 105
use FILL  FILL_4561
timestamp 1713453518
transform 1 0 744 0 -1 970
box -8 -3 16 105
use FILL  FILL_4562
timestamp 1713453518
transform 1 0 720 0 -1 970
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1713453518
transform 1 0 712 0 -1 970
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1713453518
transform 1 0 704 0 -1 970
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1713453518
transform 1 0 696 0 -1 970
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1713453518
transform 1 0 688 0 -1 970
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1713453518
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1713453518
transform 1 0 616 0 -1 970
box -8 -3 16 105
use FILL  FILL_4569
timestamp 1713453518
transform 1 0 608 0 -1 970
box -8 -3 16 105
use FILL  FILL_4570
timestamp 1713453518
transform 1 0 600 0 -1 970
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1713453518
transform 1 0 592 0 -1 970
box -8 -3 16 105
use FILL  FILL_4572
timestamp 1713453518
transform 1 0 520 0 -1 970
box -8 -3 16 105
use FILL  FILL_4573
timestamp 1713453518
transform 1 0 512 0 -1 970
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1713453518
transform 1 0 504 0 -1 970
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1713453518
transform 1 0 496 0 -1 970
box -8 -3 16 105
use FILL  FILL_4576
timestamp 1713453518
transform 1 0 456 0 -1 970
box -8 -3 16 105
use FILL  FILL_4577
timestamp 1713453518
transform 1 0 448 0 -1 970
box -8 -3 16 105
use FILL  FILL_4578
timestamp 1713453518
transform 1 0 408 0 -1 970
box -8 -3 16 105
use FILL  FILL_4579
timestamp 1713453518
transform 1 0 400 0 -1 970
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1713453518
transform 1 0 392 0 -1 970
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1713453518
transform 1 0 384 0 -1 970
box -8 -3 16 105
use FILL  FILL_4582
timestamp 1713453518
transform 1 0 320 0 -1 970
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1713453518
transform 1 0 312 0 -1 970
box -8 -3 16 105
use FILL  FILL_4584
timestamp 1713453518
transform 1 0 304 0 -1 970
box -8 -3 16 105
use FILL  FILL_4585
timestamp 1713453518
transform 1 0 296 0 -1 970
box -8 -3 16 105
use FILL  FILL_4586
timestamp 1713453518
transform 1 0 192 0 -1 970
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1713453518
transform 1 0 184 0 -1 970
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1713453518
transform 1 0 176 0 -1 970
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1713453518
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_4590
timestamp 1713453518
transform 1 0 3440 0 1 770
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1713453518
transform 1 0 3432 0 1 770
box -8 -3 16 105
use FILL  FILL_4592
timestamp 1713453518
transform 1 0 3376 0 1 770
box -8 -3 16 105
use FILL  FILL_4593
timestamp 1713453518
transform 1 0 3368 0 1 770
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1713453518
transform 1 0 3360 0 1 770
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1713453518
transform 1 0 3352 0 1 770
box -8 -3 16 105
use FILL  FILL_4596
timestamp 1713453518
transform 1 0 3344 0 1 770
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1713453518
transform 1 0 3272 0 1 770
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1713453518
transform 1 0 3264 0 1 770
box -8 -3 16 105
use FILL  FILL_4599
timestamp 1713453518
transform 1 0 3256 0 1 770
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1713453518
transform 1 0 3248 0 1 770
box -8 -3 16 105
use FILL  FILL_4601
timestamp 1713453518
transform 1 0 3240 0 1 770
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1713453518
transform 1 0 3184 0 1 770
box -8 -3 16 105
use FILL  FILL_4603
timestamp 1713453518
transform 1 0 3176 0 1 770
box -8 -3 16 105
use FILL  FILL_4604
timestamp 1713453518
transform 1 0 3168 0 1 770
box -8 -3 16 105
use FILL  FILL_4605
timestamp 1713453518
transform 1 0 3160 0 1 770
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1713453518
transform 1 0 3152 0 1 770
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1713453518
transform 1 0 3144 0 1 770
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1713453518
transform 1 0 3136 0 1 770
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1713453518
transform 1 0 3080 0 1 770
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1713453518
transform 1 0 3072 0 1 770
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1713453518
transform 1 0 3064 0 1 770
box -8 -3 16 105
use FILL  FILL_4612
timestamp 1713453518
transform 1 0 3056 0 1 770
box -8 -3 16 105
use FILL  FILL_4613
timestamp 1713453518
transform 1 0 3048 0 1 770
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1713453518
transform 1 0 3040 0 1 770
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1713453518
transform 1 0 2984 0 1 770
box -8 -3 16 105
use FILL  FILL_4616
timestamp 1713453518
transform 1 0 2976 0 1 770
box -8 -3 16 105
use FILL  FILL_4617
timestamp 1713453518
transform 1 0 2968 0 1 770
box -8 -3 16 105
use FILL  FILL_4618
timestamp 1713453518
transform 1 0 2944 0 1 770
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1713453518
transform 1 0 2936 0 1 770
box -8 -3 16 105
use FILL  FILL_4620
timestamp 1713453518
transform 1 0 2888 0 1 770
box -8 -3 16 105
use FILL  FILL_4621
timestamp 1713453518
transform 1 0 2880 0 1 770
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1713453518
transform 1 0 2872 0 1 770
box -8 -3 16 105
use FILL  FILL_4623
timestamp 1713453518
transform 1 0 2832 0 1 770
box -8 -3 16 105
use FILL  FILL_4624
timestamp 1713453518
transform 1 0 2824 0 1 770
box -8 -3 16 105
use FILL  FILL_4625
timestamp 1713453518
transform 1 0 2816 0 1 770
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1713453518
transform 1 0 2808 0 1 770
box -8 -3 16 105
use FILL  FILL_4627
timestamp 1713453518
transform 1 0 2760 0 1 770
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1713453518
transform 1 0 2736 0 1 770
box -8 -3 16 105
use FILL  FILL_4629
timestamp 1713453518
transform 1 0 2696 0 1 770
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1713453518
transform 1 0 2688 0 1 770
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1713453518
transform 1 0 2680 0 1 770
box -8 -3 16 105
use FILL  FILL_4632
timestamp 1713453518
transform 1 0 2616 0 1 770
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1713453518
transform 1 0 2608 0 1 770
box -8 -3 16 105
use FILL  FILL_4634
timestamp 1713453518
transform 1 0 2600 0 1 770
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1713453518
transform 1 0 2592 0 1 770
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1713453518
transform 1 0 2504 0 1 770
box -8 -3 16 105
use FILL  FILL_4637
timestamp 1713453518
transform 1 0 2496 0 1 770
box -8 -3 16 105
use FILL  FILL_4638
timestamp 1713453518
transform 1 0 2488 0 1 770
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1713453518
transform 1 0 2448 0 1 770
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1713453518
transform 1 0 2400 0 1 770
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1713453518
transform 1 0 2392 0 1 770
box -8 -3 16 105
use FILL  FILL_4642
timestamp 1713453518
transform 1 0 2384 0 1 770
box -8 -3 16 105
use FILL  FILL_4643
timestamp 1713453518
transform 1 0 2312 0 1 770
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1713453518
transform 1 0 2264 0 1 770
box -8 -3 16 105
use FILL  FILL_4645
timestamp 1713453518
transform 1 0 2256 0 1 770
box -8 -3 16 105
use FILL  FILL_4646
timestamp 1713453518
transform 1 0 2248 0 1 770
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1713453518
transform 1 0 2184 0 1 770
box -8 -3 16 105
use FILL  FILL_4648
timestamp 1713453518
transform 1 0 2176 0 1 770
box -8 -3 16 105
use FILL  FILL_4649
timestamp 1713453518
transform 1 0 2168 0 1 770
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1713453518
transform 1 0 2104 0 1 770
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1713453518
transform 1 0 2096 0 1 770
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1713453518
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_4653
timestamp 1713453518
transform 1 0 2008 0 1 770
box -8 -3 16 105
use FILL  FILL_4654
timestamp 1713453518
transform 1 0 2000 0 1 770
box -8 -3 16 105
use FILL  FILL_4655
timestamp 1713453518
transform 1 0 1992 0 1 770
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1713453518
transform 1 0 1984 0 1 770
box -8 -3 16 105
use FILL  FILL_4657
timestamp 1713453518
transform 1 0 1920 0 1 770
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1713453518
transform 1 0 1880 0 1 770
box -8 -3 16 105
use FILL  FILL_4659
timestamp 1713453518
transform 1 0 1872 0 1 770
box -8 -3 16 105
use FILL  FILL_4660
timestamp 1713453518
transform 1 0 1864 0 1 770
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1713453518
transform 1 0 1792 0 1 770
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1713453518
transform 1 0 1784 0 1 770
box -8 -3 16 105
use FILL  FILL_4663
timestamp 1713453518
transform 1 0 1776 0 1 770
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1713453518
transform 1 0 1768 0 1 770
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1713453518
transform 1 0 1688 0 1 770
box -8 -3 16 105
use FILL  FILL_4666
timestamp 1713453518
transform 1 0 1680 0 1 770
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1713453518
transform 1 0 1672 0 1 770
box -8 -3 16 105
use FILL  FILL_4668
timestamp 1713453518
transform 1 0 1664 0 1 770
box -8 -3 16 105
use FILL  FILL_4669
timestamp 1713453518
transform 1 0 1592 0 1 770
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1713453518
transform 1 0 1584 0 1 770
box -8 -3 16 105
use FILL  FILL_4671
timestamp 1713453518
transform 1 0 1576 0 1 770
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1713453518
transform 1 0 1536 0 1 770
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1713453518
transform 1 0 1488 0 1 770
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1713453518
transform 1 0 1480 0 1 770
box -8 -3 16 105
use FILL  FILL_4675
timestamp 1713453518
transform 1 0 1432 0 1 770
box -8 -3 16 105
use FILL  FILL_4676
timestamp 1713453518
transform 1 0 1424 0 1 770
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1713453518
transform 1 0 1376 0 1 770
box -8 -3 16 105
use FILL  FILL_4678
timestamp 1713453518
transform 1 0 1368 0 1 770
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1713453518
transform 1 0 1312 0 1 770
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1713453518
transform 1 0 1304 0 1 770
box -8 -3 16 105
use FILL  FILL_4681
timestamp 1713453518
transform 1 0 1296 0 1 770
box -8 -3 16 105
use FILL  FILL_4682
timestamp 1713453518
transform 1 0 1264 0 1 770
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1713453518
transform 1 0 1256 0 1 770
box -8 -3 16 105
use FILL  FILL_4684
timestamp 1713453518
transform 1 0 1200 0 1 770
box -8 -3 16 105
use FILL  FILL_4685
timestamp 1713453518
transform 1 0 1192 0 1 770
box -8 -3 16 105
use FILL  FILL_4686
timestamp 1713453518
transform 1 0 1184 0 1 770
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1713453518
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_4688
timestamp 1713453518
transform 1 0 1104 0 1 770
box -8 -3 16 105
use FILL  FILL_4689
timestamp 1713453518
transform 1 0 1096 0 1 770
box -8 -3 16 105
use FILL  FILL_4690
timestamp 1713453518
transform 1 0 1072 0 1 770
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1713453518
transform 1 0 1064 0 1 770
box -8 -3 16 105
use FILL  FILL_4692
timestamp 1713453518
transform 1 0 1000 0 1 770
box -8 -3 16 105
use FILL  FILL_4693
timestamp 1713453518
transform 1 0 992 0 1 770
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1713453518
transform 1 0 888 0 1 770
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1713453518
transform 1 0 880 0 1 770
box -8 -3 16 105
use FILL  FILL_4696
timestamp 1713453518
transform 1 0 840 0 1 770
box -8 -3 16 105
use FILL  FILL_4697
timestamp 1713453518
transform 1 0 832 0 1 770
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1713453518
transform 1 0 728 0 1 770
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1713453518
transform 1 0 720 0 1 770
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1713453518
transform 1 0 616 0 1 770
box -8 -3 16 105
use FILL  FILL_4701
timestamp 1713453518
transform 1 0 608 0 1 770
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1713453518
transform 1 0 600 0 1 770
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1713453518
transform 1 0 512 0 1 770
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1713453518
transform 1 0 504 0 1 770
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1713453518
transform 1 0 496 0 1 770
box -8 -3 16 105
use FILL  FILL_4706
timestamp 1713453518
transform 1 0 392 0 1 770
box -8 -3 16 105
use FILL  FILL_4707
timestamp 1713453518
transform 1 0 384 0 1 770
box -8 -3 16 105
use FILL  FILL_4708
timestamp 1713453518
transform 1 0 376 0 1 770
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1713453518
transform 1 0 368 0 1 770
box -8 -3 16 105
use FILL  FILL_4710
timestamp 1713453518
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1713453518
transform 1 0 272 0 1 770
box -8 -3 16 105
use FILL  FILL_4712
timestamp 1713453518
transform 1 0 264 0 1 770
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1713453518
transform 1 0 256 0 1 770
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1713453518
transform 1 0 152 0 1 770
box -8 -3 16 105
use FILL  FILL_4715
timestamp 1713453518
transform 1 0 144 0 1 770
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1713453518
transform 1 0 136 0 1 770
box -8 -3 16 105
use FILL  FILL_4717
timestamp 1713453518
transform 1 0 128 0 1 770
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1713453518
transform 1 0 120 0 1 770
box -8 -3 16 105
use FILL  FILL_4719
timestamp 1713453518
transform 1 0 112 0 1 770
box -8 -3 16 105
use FILL  FILL_4720
timestamp 1713453518
transform 1 0 80 0 1 770
box -8 -3 16 105
use FILL  FILL_4721
timestamp 1713453518
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_4722
timestamp 1713453518
transform 1 0 3440 0 -1 770
box -8 -3 16 105
use FILL  FILL_4723
timestamp 1713453518
transform 1 0 3368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4724
timestamp 1713453518
transform 1 0 3360 0 -1 770
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1713453518
transform 1 0 3336 0 -1 770
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1713453518
transform 1 0 3264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1713453518
transform 1 0 3256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4728
timestamp 1713453518
transform 1 0 3248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4729
timestamp 1713453518
transform 1 0 3224 0 -1 770
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1713453518
transform 1 0 3216 0 -1 770
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1713453518
transform 1 0 3160 0 -1 770
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1713453518
transform 1 0 3152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4733
timestamp 1713453518
transform 1 0 3144 0 -1 770
box -8 -3 16 105
use FILL  FILL_4734
timestamp 1713453518
transform 1 0 3080 0 -1 770
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1713453518
transform 1 0 3072 0 -1 770
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1713453518
transform 1 0 3032 0 -1 770
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1713453518
transform 1 0 3008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4738
timestamp 1713453518
transform 1 0 3000 0 -1 770
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1713453518
transform 1 0 2952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4740
timestamp 1713453518
transform 1 0 2904 0 -1 770
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1713453518
transform 1 0 2896 0 -1 770
box -8 -3 16 105
use FILL  FILL_4742
timestamp 1713453518
transform 1 0 2888 0 -1 770
box -8 -3 16 105
use FILL  FILL_4743
timestamp 1713453518
transform 1 0 2800 0 -1 770
box -8 -3 16 105
use FILL  FILL_4744
timestamp 1713453518
transform 1 0 2792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1713453518
transform 1 0 2784 0 -1 770
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1713453518
transform 1 0 2728 0 -1 770
box -8 -3 16 105
use FILL  FILL_4747
timestamp 1713453518
transform 1 0 2720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1713453518
transform 1 0 2712 0 -1 770
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1713453518
transform 1 0 2704 0 -1 770
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1713453518
transform 1 0 2640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1713453518
transform 1 0 2632 0 -1 770
box -8 -3 16 105
use FILL  FILL_4752
timestamp 1713453518
transform 1 0 2624 0 -1 770
box -8 -3 16 105
use FILL  FILL_4753
timestamp 1713453518
transform 1 0 2616 0 -1 770
box -8 -3 16 105
use FILL  FILL_4754
timestamp 1713453518
transform 1 0 2544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1713453518
transform 1 0 2536 0 -1 770
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1713453518
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use FILL  FILL_4757
timestamp 1713453518
transform 1 0 2480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1713453518
transform 1 0 2448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1713453518
transform 1 0 2440 0 -1 770
box -8 -3 16 105
use FILL  FILL_4760
timestamp 1713453518
transform 1 0 2400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1713453518
transform 1 0 2392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4762
timestamp 1713453518
transform 1 0 2384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1713453518
transform 1 0 2336 0 -1 770
box -8 -3 16 105
use FILL  FILL_4764
timestamp 1713453518
transform 1 0 2328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4765
timestamp 1713453518
transform 1 0 2272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4766
timestamp 1713453518
transform 1 0 2264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4767
timestamp 1713453518
transform 1 0 2256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1713453518
transform 1 0 2248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1713453518
transform 1 0 2240 0 -1 770
box -8 -3 16 105
use FILL  FILL_4770
timestamp 1713453518
transform 1 0 2168 0 -1 770
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1713453518
transform 1 0 2160 0 -1 770
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1713453518
transform 1 0 2152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1713453518
transform 1 0 2104 0 -1 770
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1713453518
transform 1 0 2096 0 -1 770
box -8 -3 16 105
use FILL  FILL_4775
timestamp 1713453518
transform 1 0 2088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1713453518
transform 1 0 2016 0 -1 770
box -8 -3 16 105
use FILL  FILL_4777
timestamp 1713453518
transform 1 0 2008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4778
timestamp 1713453518
transform 1 0 2000 0 -1 770
box -8 -3 16 105
use FILL  FILL_4779
timestamp 1713453518
transform 1 0 1960 0 -1 770
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1713453518
transform 1 0 1952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4781
timestamp 1713453518
transform 1 0 1888 0 -1 770
box -8 -3 16 105
use FILL  FILL_4782
timestamp 1713453518
transform 1 0 1880 0 -1 770
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1713453518
transform 1 0 1872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4784
timestamp 1713453518
transform 1 0 1800 0 -1 770
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1713453518
transform 1 0 1792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4786
timestamp 1713453518
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1713453518
transform 1 0 1744 0 -1 770
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1713453518
transform 1 0 1704 0 -1 770
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1713453518
transform 1 0 1656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4790
timestamp 1713453518
transform 1 0 1648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1713453518
transform 1 0 1576 0 -1 770
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1713453518
transform 1 0 1568 0 -1 770
box -8 -3 16 105
use FILL  FILL_4793
timestamp 1713453518
transform 1 0 1560 0 -1 770
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1713453518
transform 1 0 1552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4795
timestamp 1713453518
transform 1 0 1480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4796
timestamp 1713453518
transform 1 0 1440 0 -1 770
box -8 -3 16 105
use FILL  FILL_4797
timestamp 1713453518
transform 1 0 1432 0 -1 770
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1713453518
transform 1 0 1392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1713453518
transform 1 0 1344 0 -1 770
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1713453518
transform 1 0 1336 0 -1 770
box -8 -3 16 105
use FILL  FILL_4801
timestamp 1713453518
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4802
timestamp 1713453518
transform 1 0 1264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4803
timestamp 1713453518
transform 1 0 1256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1713453518
transform 1 0 1248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4805
timestamp 1713453518
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_4806
timestamp 1713453518
transform 1 0 1176 0 -1 770
box -8 -3 16 105
use FILL  FILL_4807
timestamp 1713453518
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use FILL  FILL_4808
timestamp 1713453518
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4809
timestamp 1713453518
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1713453518
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1713453518
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1713453518
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_4813
timestamp 1713453518
transform 1 0 1000 0 -1 770
box -8 -3 16 105
use FILL  FILL_4814
timestamp 1713453518
transform 1 0 992 0 -1 770
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1713453518
transform 1 0 984 0 -1 770
box -8 -3 16 105
use FILL  FILL_4816
timestamp 1713453518
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_4817
timestamp 1713453518
transform 1 0 872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1713453518
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_4819
timestamp 1713453518
transform 1 0 760 0 -1 770
box -8 -3 16 105
use FILL  FILL_4820
timestamp 1713453518
transform 1 0 752 0 -1 770
box -8 -3 16 105
use FILL  FILL_4821
timestamp 1713453518
transform 1 0 744 0 -1 770
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1713453518
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1713453518
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4824
timestamp 1713453518
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4825
timestamp 1713453518
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4826
timestamp 1713453518
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_4827
timestamp 1713453518
transform 1 0 624 0 -1 770
box -8 -3 16 105
use FILL  FILL_4828
timestamp 1713453518
transform 1 0 616 0 -1 770
box -8 -3 16 105
use FILL  FILL_4829
timestamp 1713453518
transform 1 0 536 0 -1 770
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1713453518
transform 1 0 528 0 -1 770
box -8 -3 16 105
use FILL  FILL_4831
timestamp 1713453518
transform 1 0 520 0 -1 770
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1713453518
transform 1 0 512 0 -1 770
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1713453518
transform 1 0 504 0 -1 770
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1713453518
transform 1 0 424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1713453518
transform 1 0 416 0 -1 770
box -8 -3 16 105
use FILL  FILL_4836
timestamp 1713453518
transform 1 0 408 0 -1 770
box -8 -3 16 105
use FILL  FILL_4837
timestamp 1713453518
transform 1 0 400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4838
timestamp 1713453518
transform 1 0 296 0 -1 770
box -8 -3 16 105
use FILL  FILL_4839
timestamp 1713453518
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1713453518
transform 1 0 280 0 -1 770
box -8 -3 16 105
use FILL  FILL_4841
timestamp 1713453518
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1713453518
transform 1 0 264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4843
timestamp 1713453518
transform 1 0 200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4844
timestamp 1713453518
transform 1 0 192 0 -1 770
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1713453518
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_4846
timestamp 1713453518
transform 1 0 3440 0 1 570
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1713453518
transform 1 0 3432 0 1 570
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1713453518
transform 1 0 3352 0 1 570
box -8 -3 16 105
use FILL  FILL_4849
timestamp 1713453518
transform 1 0 3344 0 1 570
box -8 -3 16 105
use FILL  FILL_4850
timestamp 1713453518
transform 1 0 3336 0 1 570
box -8 -3 16 105
use FILL  FILL_4851
timestamp 1713453518
transform 1 0 3328 0 1 570
box -8 -3 16 105
use FILL  FILL_4852
timestamp 1713453518
transform 1 0 3240 0 1 570
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1713453518
transform 1 0 3232 0 1 570
box -8 -3 16 105
use FILL  FILL_4854
timestamp 1713453518
transform 1 0 3224 0 1 570
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1713453518
transform 1 0 3216 0 1 570
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1713453518
transform 1 0 3208 0 1 570
box -8 -3 16 105
use FILL  FILL_4857
timestamp 1713453518
transform 1 0 3152 0 1 570
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1713453518
transform 1 0 3144 0 1 570
box -8 -3 16 105
use FILL  FILL_4859
timestamp 1713453518
transform 1 0 3136 0 1 570
box -8 -3 16 105
use FILL  FILL_4860
timestamp 1713453518
transform 1 0 3128 0 1 570
box -8 -3 16 105
use FILL  FILL_4861
timestamp 1713453518
transform 1 0 3120 0 1 570
box -8 -3 16 105
use FILL  FILL_4862
timestamp 1713453518
transform 1 0 3064 0 1 570
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1713453518
transform 1 0 3056 0 1 570
box -8 -3 16 105
use FILL  FILL_4864
timestamp 1713453518
transform 1 0 3048 0 1 570
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1713453518
transform 1 0 3008 0 1 570
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1713453518
transform 1 0 3000 0 1 570
box -8 -3 16 105
use FILL  FILL_4867
timestamp 1713453518
transform 1 0 2968 0 1 570
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1713453518
transform 1 0 2960 0 1 570
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1713453518
transform 1 0 2952 0 1 570
box -8 -3 16 105
use FILL  FILL_4870
timestamp 1713453518
transform 1 0 2904 0 1 570
box -8 -3 16 105
use FILL  FILL_4871
timestamp 1713453518
transform 1 0 2896 0 1 570
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1713453518
transform 1 0 2888 0 1 570
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1713453518
transform 1 0 2856 0 1 570
box -8 -3 16 105
use FILL  FILL_4874
timestamp 1713453518
transform 1 0 2848 0 1 570
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1713453518
transform 1 0 2840 0 1 570
box -8 -3 16 105
use FILL  FILL_4876
timestamp 1713453518
transform 1 0 2792 0 1 570
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1713453518
transform 1 0 2784 0 1 570
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1713453518
transform 1 0 2776 0 1 570
box -8 -3 16 105
use FILL  FILL_4879
timestamp 1713453518
transform 1 0 2744 0 1 570
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1713453518
transform 1 0 2736 0 1 570
box -8 -3 16 105
use FILL  FILL_4881
timestamp 1713453518
transform 1 0 2696 0 1 570
box -8 -3 16 105
use FILL  FILL_4882
timestamp 1713453518
transform 1 0 2688 0 1 570
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1713453518
transform 1 0 2664 0 1 570
box -8 -3 16 105
use FILL  FILL_4884
timestamp 1713453518
transform 1 0 2624 0 1 570
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1713453518
transform 1 0 2616 0 1 570
box -8 -3 16 105
use FILL  FILL_4886
timestamp 1713453518
transform 1 0 2608 0 1 570
box -8 -3 16 105
use FILL  FILL_4887
timestamp 1713453518
transform 1 0 2600 0 1 570
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1713453518
transform 1 0 2560 0 1 570
box -8 -3 16 105
use FILL  FILL_4889
timestamp 1713453518
transform 1 0 2520 0 1 570
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1713453518
transform 1 0 2512 0 1 570
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1713453518
transform 1 0 2504 0 1 570
box -8 -3 16 105
use FILL  FILL_4892
timestamp 1713453518
transform 1 0 2496 0 1 570
box -8 -3 16 105
use FILL  FILL_4893
timestamp 1713453518
transform 1 0 2424 0 1 570
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1713453518
transform 1 0 2416 0 1 570
box -8 -3 16 105
use FILL  FILL_4895
timestamp 1713453518
transform 1 0 2368 0 1 570
box -8 -3 16 105
use FILL  FILL_4896
timestamp 1713453518
transform 1 0 2360 0 1 570
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1713453518
transform 1 0 2352 0 1 570
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1713453518
transform 1 0 2272 0 1 570
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1713453518
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_4900
timestamp 1713453518
transform 1 0 2256 0 1 570
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1713453518
transform 1 0 2248 0 1 570
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1713453518
transform 1 0 2240 0 1 570
box -8 -3 16 105
use FILL  FILL_4903
timestamp 1713453518
transform 1 0 2176 0 1 570
box -8 -3 16 105
use FILL  FILL_4904
timestamp 1713453518
transform 1 0 2168 0 1 570
box -8 -3 16 105
use FILL  FILL_4905
timestamp 1713453518
transform 1 0 2112 0 1 570
box -8 -3 16 105
use FILL  FILL_4906
timestamp 1713453518
transform 1 0 2104 0 1 570
box -8 -3 16 105
use FILL  FILL_4907
timestamp 1713453518
transform 1 0 2096 0 1 570
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1713453518
transform 1 0 2088 0 1 570
box -8 -3 16 105
use FILL  FILL_4909
timestamp 1713453518
transform 1 0 2016 0 1 570
box -8 -3 16 105
use FILL  FILL_4910
timestamp 1713453518
transform 1 0 2008 0 1 570
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1713453518
transform 1 0 1968 0 1 570
box -8 -3 16 105
use FILL  FILL_4912
timestamp 1713453518
transform 1 0 1920 0 1 570
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1713453518
transform 1 0 1912 0 1 570
box -8 -3 16 105
use FILL  FILL_4914
timestamp 1713453518
transform 1 0 1904 0 1 570
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1713453518
transform 1 0 1856 0 1 570
box -8 -3 16 105
use FILL  FILL_4916
timestamp 1713453518
transform 1 0 1792 0 1 570
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1713453518
transform 1 0 1784 0 1 570
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1713453518
transform 1 0 1776 0 1 570
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1713453518
transform 1 0 1768 0 1 570
box -8 -3 16 105
use FILL  FILL_4920
timestamp 1713453518
transform 1 0 1704 0 1 570
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1713453518
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1713453518
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_4923
timestamp 1713453518
transform 1 0 1656 0 1 570
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1713453518
transform 1 0 1584 0 1 570
box -8 -3 16 105
use FILL  FILL_4925
timestamp 1713453518
transform 1 0 1576 0 1 570
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1713453518
transform 1 0 1568 0 1 570
box -8 -3 16 105
use FILL  FILL_4927
timestamp 1713453518
transform 1 0 1560 0 1 570
box -8 -3 16 105
use FILL  FILL_4928
timestamp 1713453518
transform 1 0 1480 0 1 570
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1713453518
transform 1 0 1472 0 1 570
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1713453518
transform 1 0 1464 0 1 570
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1713453518
transform 1 0 1408 0 1 570
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1713453518
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_4933
timestamp 1713453518
transform 1 0 1320 0 1 570
box -8 -3 16 105
use FILL  FILL_4934
timestamp 1713453518
transform 1 0 1312 0 1 570
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1713453518
transform 1 0 1304 0 1 570
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1713453518
transform 1 0 1296 0 1 570
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1713453518
transform 1 0 1240 0 1 570
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1713453518
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_4939
timestamp 1713453518
transform 1 0 1200 0 1 570
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1713453518
transform 1 0 1192 0 1 570
box -8 -3 16 105
use FILL  FILL_4941
timestamp 1713453518
transform 1 0 1184 0 1 570
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1713453518
transform 1 0 1112 0 1 570
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1713453518
transform 1 0 1104 0 1 570
box -8 -3 16 105
use FILL  FILL_4944
timestamp 1713453518
transform 1 0 1096 0 1 570
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1713453518
transform 1 0 1088 0 1 570
box -8 -3 16 105
use FILL  FILL_4946
timestamp 1713453518
transform 1 0 1056 0 1 570
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1713453518
transform 1 0 1000 0 1 570
box -8 -3 16 105
use FILL  FILL_4948
timestamp 1713453518
transform 1 0 992 0 1 570
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1713453518
transform 1 0 888 0 1 570
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1713453518
transform 1 0 880 0 1 570
box -8 -3 16 105
use FILL  FILL_4951
timestamp 1713453518
transform 1 0 872 0 1 570
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1713453518
transform 1 0 824 0 1 570
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1713453518
transform 1 0 816 0 1 570
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1713453518
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_4955
timestamp 1713453518
transform 1 0 760 0 1 570
box -8 -3 16 105
use FILL  FILL_4956
timestamp 1713453518
transform 1 0 712 0 1 570
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1713453518
transform 1 0 704 0 1 570
box -8 -3 16 105
use FILL  FILL_4958
timestamp 1713453518
transform 1 0 696 0 1 570
box -8 -3 16 105
use FILL  FILL_4959
timestamp 1713453518
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_4960
timestamp 1713453518
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1713453518
transform 1 0 576 0 1 570
box -8 -3 16 105
use FILL  FILL_4962
timestamp 1713453518
transform 1 0 472 0 1 570
box -8 -3 16 105
use FILL  FILL_4963
timestamp 1713453518
transform 1 0 464 0 1 570
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1713453518
transform 1 0 456 0 1 570
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1713453518
transform 1 0 408 0 1 570
box -8 -3 16 105
use FILL  FILL_4966
timestamp 1713453518
transform 1 0 400 0 1 570
box -8 -3 16 105
use FILL  FILL_4967
timestamp 1713453518
transform 1 0 296 0 1 570
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1713453518
transform 1 0 288 0 1 570
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1713453518
transform 1 0 280 0 1 570
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1713453518
transform 1 0 272 0 1 570
box -8 -3 16 105
use FILL  FILL_4971
timestamp 1713453518
transform 1 0 264 0 1 570
box -8 -3 16 105
use FILL  FILL_4972
timestamp 1713453518
transform 1 0 208 0 1 570
box -8 -3 16 105
use FILL  FILL_4973
timestamp 1713453518
transform 1 0 200 0 1 570
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1713453518
transform 1 0 192 0 1 570
box -8 -3 16 105
use FILL  FILL_4975
timestamp 1713453518
transform 1 0 184 0 1 570
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1713453518
transform 1 0 176 0 1 570
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1713453518
transform 1 0 168 0 1 570
box -8 -3 16 105
use FILL  FILL_4978
timestamp 1713453518
transform 1 0 160 0 1 570
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1713453518
transform 1 0 96 0 1 570
box -8 -3 16 105
use FILL  FILL_4980
timestamp 1713453518
transform 1 0 88 0 1 570
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1713453518
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_4982
timestamp 1713453518
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1713453518
transform 1 0 3384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1713453518
transform 1 0 3376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1713453518
transform 1 0 3296 0 -1 570
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1713453518
transform 1 0 3288 0 -1 570
box -8 -3 16 105
use FILL  FILL_4987
timestamp 1713453518
transform 1 0 3280 0 -1 570
box -8 -3 16 105
use FILL  FILL_4988
timestamp 1713453518
transform 1 0 3272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1713453518
transform 1 0 3208 0 -1 570
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1713453518
transform 1 0 3200 0 -1 570
box -8 -3 16 105
use FILL  FILL_4991
timestamp 1713453518
transform 1 0 3192 0 -1 570
box -8 -3 16 105
use FILL  FILL_4992
timestamp 1713453518
transform 1 0 3184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1713453518
transform 1 0 3120 0 -1 570
box -8 -3 16 105
use FILL  FILL_4994
timestamp 1713453518
transform 1 0 3112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4995
timestamp 1713453518
transform 1 0 3104 0 -1 570
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1713453518
transform 1 0 3096 0 -1 570
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1713453518
transform 1 0 3056 0 -1 570
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1713453518
transform 1 0 3048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1713453518
transform 1 0 3040 0 -1 570
box -8 -3 16 105
use FILL  FILL_5000
timestamp 1713453518
transform 1 0 3032 0 -1 570
box -8 -3 16 105
use FILL  FILL_5001
timestamp 1713453518
transform 1 0 3024 0 -1 570
box -8 -3 16 105
use FILL  FILL_5002
timestamp 1713453518
transform 1 0 3016 0 -1 570
box -8 -3 16 105
use FILL  FILL_5003
timestamp 1713453518
transform 1 0 2912 0 -1 570
box -8 -3 16 105
use FILL  FILL_5004
timestamp 1713453518
transform 1 0 2904 0 -1 570
box -8 -3 16 105
use FILL  FILL_5005
timestamp 1713453518
transform 1 0 2896 0 -1 570
box -8 -3 16 105
use FILL  FILL_5006
timestamp 1713453518
transform 1 0 2888 0 -1 570
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1713453518
transform 1 0 2840 0 -1 570
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1713453518
transform 1 0 2832 0 -1 570
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1713453518
transform 1 0 2824 0 -1 570
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1713453518
transform 1 0 2800 0 -1 570
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1713453518
transform 1 0 2792 0 -1 570
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1713453518
transform 1 0 2744 0 -1 570
box -8 -3 16 105
use FILL  FILL_5013
timestamp 1713453518
transform 1 0 2736 0 -1 570
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1713453518
transform 1 0 2704 0 -1 570
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1713453518
transform 1 0 2696 0 -1 570
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1713453518
transform 1 0 2688 0 -1 570
box -8 -3 16 105
use FILL  FILL_5017
timestamp 1713453518
transform 1 0 2680 0 -1 570
box -8 -3 16 105
use FILL  FILL_5018
timestamp 1713453518
transform 1 0 2608 0 -1 570
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1713453518
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1713453518
transform 1 0 2592 0 -1 570
box -8 -3 16 105
use FILL  FILL_5021
timestamp 1713453518
transform 1 0 2528 0 -1 570
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1713453518
transform 1 0 2520 0 -1 570
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1713453518
transform 1 0 2512 0 -1 570
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1713453518
transform 1 0 2480 0 -1 570
box -8 -3 16 105
use FILL  FILL_5025
timestamp 1713453518
transform 1 0 2472 0 -1 570
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1713453518
transform 1 0 2416 0 -1 570
box -8 -3 16 105
use FILL  FILL_5027
timestamp 1713453518
transform 1 0 2408 0 -1 570
box -8 -3 16 105
use FILL  FILL_5028
timestamp 1713453518
transform 1 0 2400 0 -1 570
box -8 -3 16 105
use FILL  FILL_5029
timestamp 1713453518
transform 1 0 2360 0 -1 570
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1713453518
transform 1 0 2312 0 -1 570
box -8 -3 16 105
use FILL  FILL_5031
timestamp 1713453518
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use FILL  FILL_5032
timestamp 1713453518
transform 1 0 2296 0 -1 570
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1713453518
transform 1 0 2248 0 -1 570
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1713453518
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_5035
timestamp 1713453518
transform 1 0 2184 0 -1 570
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1713453518
transform 1 0 2176 0 -1 570
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1713453518
transform 1 0 2168 0 -1 570
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1713453518
transform 1 0 2096 0 -1 570
box -8 -3 16 105
use FILL  FILL_5039
timestamp 1713453518
transform 1 0 2088 0 -1 570
box -8 -3 16 105
use FILL  FILL_5040
timestamp 1713453518
transform 1 0 2080 0 -1 570
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1713453518
transform 1 0 2072 0 -1 570
box -8 -3 16 105
use FILL  FILL_5042
timestamp 1713453518
transform 1 0 2000 0 -1 570
box -8 -3 16 105
use FILL  FILL_5043
timestamp 1713453518
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1713453518
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1713453518
transform 1 0 1976 0 -1 570
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1713453518
transform 1 0 1896 0 -1 570
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1713453518
transform 1 0 1888 0 -1 570
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1713453518
transform 1 0 1880 0 -1 570
box -8 -3 16 105
use FILL  FILL_5049
timestamp 1713453518
transform 1 0 1872 0 -1 570
box -8 -3 16 105
use FILL  FILL_5050
timestamp 1713453518
transform 1 0 1800 0 -1 570
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1713453518
transform 1 0 1792 0 -1 570
box -8 -3 16 105
use FILL  FILL_5052
timestamp 1713453518
transform 1 0 1752 0 -1 570
box -8 -3 16 105
use FILL  FILL_5053
timestamp 1713453518
transform 1 0 1744 0 -1 570
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1713453518
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1713453518
transform 1 0 1672 0 -1 570
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1713453518
transform 1 0 1664 0 -1 570
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1713453518
transform 1 0 1656 0 -1 570
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1713453518
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1713453518
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1713453518
transform 1 0 1520 0 -1 570
box -8 -3 16 105
use FILL  FILL_5061
timestamp 1713453518
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_5062
timestamp 1713453518
transform 1 0 1504 0 -1 570
box -8 -3 16 105
use FILL  FILL_5063
timestamp 1713453518
transform 1 0 1496 0 -1 570
box -8 -3 16 105
use FILL  FILL_5064
timestamp 1713453518
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use FILL  FILL_5065
timestamp 1713453518
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1713453518
transform 1 0 1376 0 -1 570
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1713453518
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use FILL  FILL_5068
timestamp 1713453518
transform 1 0 1360 0 -1 570
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1713453518
transform 1 0 1280 0 -1 570
box -8 -3 16 105
use FILL  FILL_5070
timestamp 1713453518
transform 1 0 1272 0 -1 570
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1713453518
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1713453518
transform 1 0 1256 0 -1 570
box -8 -3 16 105
use FILL  FILL_5073
timestamp 1713453518
transform 1 0 1224 0 -1 570
box -8 -3 16 105
use FILL  FILL_5074
timestamp 1713453518
transform 1 0 1160 0 -1 570
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1713453518
transform 1 0 1152 0 -1 570
box -8 -3 16 105
use FILL  FILL_5076
timestamp 1713453518
transform 1 0 1144 0 -1 570
box -8 -3 16 105
use FILL  FILL_5077
timestamp 1713453518
transform 1 0 1104 0 -1 570
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1713453518
transform 1 0 1096 0 -1 570
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1713453518
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1713453518
transform 1 0 1016 0 -1 570
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1713453518
transform 1 0 1008 0 -1 570
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1713453518
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use FILL  FILL_5083
timestamp 1713453518
transform 1 0 896 0 -1 570
box -8 -3 16 105
use FILL  FILL_5084
timestamp 1713453518
transform 1 0 888 0 -1 570
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1713453518
transform 1 0 784 0 -1 570
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1713453518
transform 1 0 776 0 -1 570
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1713453518
transform 1 0 672 0 -1 570
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1713453518
transform 1 0 664 0 -1 570
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1713453518
transform 1 0 600 0 -1 570
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1713453518
transform 1 0 592 0 -1 570
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1713453518
transform 1 0 520 0 -1 570
box -8 -3 16 105
use FILL  FILL_5092
timestamp 1713453518
transform 1 0 512 0 -1 570
box -8 -3 16 105
use FILL  FILL_5093
timestamp 1713453518
transform 1 0 504 0 -1 570
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1713453518
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_5095
timestamp 1713453518
transform 1 0 368 0 -1 570
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1713453518
transform 1 0 360 0 -1 570
box -8 -3 16 105
use FILL  FILL_5097
timestamp 1713453518
transform 1 0 256 0 -1 570
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1713453518
transform 1 0 248 0 -1 570
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1713453518
transform 1 0 240 0 -1 570
box -8 -3 16 105
use FILL  FILL_5100
timestamp 1713453518
transform 1 0 192 0 -1 570
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1713453518
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_5102
timestamp 1713453518
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1713453518
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1713453518
transform 1 0 3440 0 1 370
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1713453518
transform 1 0 3328 0 1 370
box -8 -3 16 105
use FILL  FILL_5106
timestamp 1713453518
transform 1 0 3320 0 1 370
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1713453518
transform 1 0 3224 0 1 370
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1713453518
transform 1 0 3216 0 1 370
box -8 -3 16 105
use FILL  FILL_5109
timestamp 1713453518
transform 1 0 3208 0 1 370
box -8 -3 16 105
use FILL  FILL_5110
timestamp 1713453518
transform 1 0 3200 0 1 370
box -8 -3 16 105
use FILL  FILL_5111
timestamp 1713453518
transform 1 0 3192 0 1 370
box -8 -3 16 105
use FILL  FILL_5112
timestamp 1713453518
transform 1 0 3120 0 1 370
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1713453518
transform 1 0 3112 0 1 370
box -8 -3 16 105
use FILL  FILL_5114
timestamp 1713453518
transform 1 0 3104 0 1 370
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1713453518
transform 1 0 3096 0 1 370
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1713453518
transform 1 0 2992 0 1 370
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1713453518
transform 1 0 2984 0 1 370
box -8 -3 16 105
use FILL  FILL_5118
timestamp 1713453518
transform 1 0 2976 0 1 370
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1713453518
transform 1 0 2968 0 1 370
box -8 -3 16 105
use FILL  FILL_5120
timestamp 1713453518
transform 1 0 2888 0 1 370
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1713453518
transform 1 0 2880 0 1 370
box -8 -3 16 105
use FILL  FILL_5122
timestamp 1713453518
transform 1 0 2872 0 1 370
box -8 -3 16 105
use FILL  FILL_5123
timestamp 1713453518
transform 1 0 2864 0 1 370
box -8 -3 16 105
use FILL  FILL_5124
timestamp 1713453518
transform 1 0 2856 0 1 370
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1713453518
transform 1 0 2784 0 1 370
box -8 -3 16 105
use FILL  FILL_5126
timestamp 1713453518
transform 1 0 2776 0 1 370
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1713453518
transform 1 0 2768 0 1 370
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1713453518
transform 1 0 2664 0 1 370
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1713453518
transform 1 0 2656 0 1 370
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1713453518
transform 1 0 2648 0 1 370
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1713453518
transform 1 0 2560 0 1 370
box -8 -3 16 105
use FILL  FILL_5132
timestamp 1713453518
transform 1 0 2552 0 1 370
box -8 -3 16 105
use FILL  FILL_5133
timestamp 1713453518
transform 1 0 2544 0 1 370
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1713453518
transform 1 0 2536 0 1 370
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1713453518
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1713453518
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_5137
timestamp 1713453518
transform 1 0 2424 0 1 370
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1713453518
transform 1 0 2416 0 1 370
box -8 -3 16 105
use FILL  FILL_5139
timestamp 1713453518
transform 1 0 2368 0 1 370
box -8 -3 16 105
use FILL  FILL_5140
timestamp 1713453518
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1713453518
transform 1 0 2304 0 1 370
box -8 -3 16 105
use FILL  FILL_5142
timestamp 1713453518
transform 1 0 2296 0 1 370
box -8 -3 16 105
use FILL  FILL_5143
timestamp 1713453518
transform 1 0 2288 0 1 370
box -8 -3 16 105
use FILL  FILL_5144
timestamp 1713453518
transform 1 0 2280 0 1 370
box -8 -3 16 105
use FILL  FILL_5145
timestamp 1713453518
transform 1 0 2224 0 1 370
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1713453518
transform 1 0 2216 0 1 370
box -8 -3 16 105
use FILL  FILL_5147
timestamp 1713453518
transform 1 0 2208 0 1 370
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1713453518
transform 1 0 2184 0 1 370
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1713453518
transform 1 0 2176 0 1 370
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1713453518
transform 1 0 2168 0 1 370
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1713453518
transform 1 0 2104 0 1 370
box -8 -3 16 105
use FILL  FILL_5152
timestamp 1713453518
transform 1 0 2096 0 1 370
box -8 -3 16 105
use FILL  FILL_5153
timestamp 1713453518
transform 1 0 2088 0 1 370
box -8 -3 16 105
use FILL  FILL_5154
timestamp 1713453518
transform 1 0 2080 0 1 370
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1713453518
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1713453518
transform 1 0 2064 0 1 370
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1713453518
transform 1 0 1992 0 1 370
box -8 -3 16 105
use FILL  FILL_5158
timestamp 1713453518
transform 1 0 1984 0 1 370
box -8 -3 16 105
use FILL  FILL_5159
timestamp 1713453518
transform 1 0 1976 0 1 370
box -8 -3 16 105
use FILL  FILL_5160
timestamp 1713453518
transform 1 0 1968 0 1 370
box -8 -3 16 105
use FILL  FILL_5161
timestamp 1713453518
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_5162
timestamp 1713453518
transform 1 0 1952 0 1 370
box -8 -3 16 105
use FILL  FILL_5163
timestamp 1713453518
transform 1 0 1912 0 1 370
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1713453518
transform 1 0 1872 0 1 370
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1713453518
transform 1 0 1864 0 1 370
box -8 -3 16 105
use FILL  FILL_5166
timestamp 1713453518
transform 1 0 1856 0 1 370
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1713453518
transform 1 0 1848 0 1 370
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1713453518
transform 1 0 1840 0 1 370
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1713453518
transform 1 0 1832 0 1 370
box -8 -3 16 105
use FILL  FILL_5170
timestamp 1713453518
transform 1 0 1824 0 1 370
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1713453518
transform 1 0 1752 0 1 370
box -8 -3 16 105
use FILL  FILL_5172
timestamp 1713453518
transform 1 0 1744 0 1 370
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1713453518
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_5174
timestamp 1713453518
transform 1 0 1728 0 1 370
box -8 -3 16 105
use FILL  FILL_5175
timestamp 1713453518
transform 1 0 1720 0 1 370
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1713453518
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_5177
timestamp 1713453518
transform 1 0 1656 0 1 370
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1713453518
transform 1 0 1632 0 1 370
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1713453518
transform 1 0 1624 0 1 370
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1713453518
transform 1 0 1592 0 1 370
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1713453518
transform 1 0 1584 0 1 370
box -8 -3 16 105
use FILL  FILL_5182
timestamp 1713453518
transform 1 0 1576 0 1 370
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1713453518
transform 1 0 1520 0 1 370
box -8 -3 16 105
use FILL  FILL_5184
timestamp 1713453518
transform 1 0 1512 0 1 370
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1713453518
transform 1 0 1504 0 1 370
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1713453518
transform 1 0 1432 0 1 370
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1713453518
transform 1 0 1424 0 1 370
box -8 -3 16 105
use FILL  FILL_5188
timestamp 1713453518
transform 1 0 1416 0 1 370
box -8 -3 16 105
use FILL  FILL_5189
timestamp 1713453518
transform 1 0 1408 0 1 370
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1713453518
transform 1 0 1368 0 1 370
box -8 -3 16 105
use FILL  FILL_5191
timestamp 1713453518
transform 1 0 1320 0 1 370
box -8 -3 16 105
use FILL  FILL_5192
timestamp 1713453518
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_5193
timestamp 1713453518
transform 1 0 1304 0 1 370
box -8 -3 16 105
use FILL  FILL_5194
timestamp 1713453518
transform 1 0 1248 0 1 370
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1713453518
transform 1 0 1240 0 1 370
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1713453518
transform 1 0 1232 0 1 370
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1713453518
transform 1 0 1224 0 1 370
box -8 -3 16 105
use FILL  FILL_5198
timestamp 1713453518
transform 1 0 1152 0 1 370
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1713453518
transform 1 0 1144 0 1 370
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1713453518
transform 1 0 1136 0 1 370
box -8 -3 16 105
use FILL  FILL_5201
timestamp 1713453518
transform 1 0 1128 0 1 370
box -8 -3 16 105
use FILL  FILL_5202
timestamp 1713453518
transform 1 0 1048 0 1 370
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1713453518
transform 1 0 1040 0 1 370
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1713453518
transform 1 0 1032 0 1 370
box -8 -3 16 105
use FILL  FILL_5205
timestamp 1713453518
transform 1 0 928 0 1 370
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1713453518
transform 1 0 920 0 1 370
box -8 -3 16 105
use FILL  FILL_5207
timestamp 1713453518
transform 1 0 912 0 1 370
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1713453518
transform 1 0 904 0 1 370
box -8 -3 16 105
use FILL  FILL_5209
timestamp 1713453518
transform 1 0 872 0 1 370
box -8 -3 16 105
use FILL  FILL_5210
timestamp 1713453518
transform 1 0 864 0 1 370
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1713453518
transform 1 0 856 0 1 370
box -8 -3 16 105
use FILL  FILL_5212
timestamp 1713453518
transform 1 0 800 0 1 370
box -8 -3 16 105
use FILL  FILL_5213
timestamp 1713453518
transform 1 0 792 0 1 370
box -8 -3 16 105
use FILL  FILL_5214
timestamp 1713453518
transform 1 0 784 0 1 370
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1713453518
transform 1 0 776 0 1 370
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1713453518
transform 1 0 720 0 1 370
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1713453518
transform 1 0 712 0 1 370
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1713453518
transform 1 0 704 0 1 370
box -8 -3 16 105
use FILL  FILL_5219
timestamp 1713453518
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_5220
timestamp 1713453518
transform 1 0 632 0 1 370
box -8 -3 16 105
use FILL  FILL_5221
timestamp 1713453518
transform 1 0 624 0 1 370
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1713453518
transform 1 0 616 0 1 370
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1713453518
transform 1 0 608 0 1 370
box -8 -3 16 105
use FILL  FILL_5224
timestamp 1713453518
transform 1 0 600 0 1 370
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1713453518
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_5226
timestamp 1713453518
transform 1 0 528 0 1 370
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1713453518
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_5228
timestamp 1713453518
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_5229
timestamp 1713453518
transform 1 0 448 0 1 370
box -8 -3 16 105
use FILL  FILL_5230
timestamp 1713453518
transform 1 0 440 0 1 370
box -8 -3 16 105
use FILL  FILL_5231
timestamp 1713453518
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1713453518
transform 1 0 376 0 1 370
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1713453518
transform 1 0 368 0 1 370
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1713453518
transform 1 0 336 0 1 370
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1713453518
transform 1 0 328 0 1 370
box -8 -3 16 105
use FILL  FILL_5236
timestamp 1713453518
transform 1 0 272 0 1 370
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1713453518
transform 1 0 264 0 1 370
box -8 -3 16 105
use FILL  FILL_5238
timestamp 1713453518
transform 1 0 256 0 1 370
box -8 -3 16 105
use FILL  FILL_5239
timestamp 1713453518
transform 1 0 248 0 1 370
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1713453518
transform 1 0 144 0 1 370
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1713453518
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_5242
timestamp 1713453518
transform 1 0 128 0 1 370
box -8 -3 16 105
use FILL  FILL_5243
timestamp 1713453518
transform 1 0 120 0 1 370
box -8 -3 16 105
use FILL  FILL_5244
timestamp 1713453518
transform 1 0 3440 0 -1 370
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1713453518
transform 1 0 3432 0 -1 370
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1713453518
transform 1 0 3352 0 -1 370
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1713453518
transform 1 0 3344 0 -1 370
box -8 -3 16 105
use FILL  FILL_5248
timestamp 1713453518
transform 1 0 3336 0 -1 370
box -8 -3 16 105
use FILL  FILL_5249
timestamp 1713453518
transform 1 0 3272 0 -1 370
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1713453518
transform 1 0 3264 0 -1 370
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1713453518
transform 1 0 3256 0 -1 370
box -8 -3 16 105
use FILL  FILL_5252
timestamp 1713453518
transform 1 0 3248 0 -1 370
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1713453518
transform 1 0 3160 0 -1 370
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1713453518
transform 1 0 3152 0 -1 370
box -8 -3 16 105
use FILL  FILL_5255
timestamp 1713453518
transform 1 0 3144 0 -1 370
box -8 -3 16 105
use FILL  FILL_5256
timestamp 1713453518
transform 1 0 3136 0 -1 370
box -8 -3 16 105
use FILL  FILL_5257
timestamp 1713453518
transform 1 0 3032 0 -1 370
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1713453518
transform 1 0 3024 0 -1 370
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1713453518
transform 1 0 3016 0 -1 370
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1713453518
transform 1 0 3008 0 -1 370
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1713453518
transform 1 0 3000 0 -1 370
box -8 -3 16 105
use FILL  FILL_5262
timestamp 1713453518
transform 1 0 2992 0 -1 370
box -8 -3 16 105
use FILL  FILL_5263
timestamp 1713453518
transform 1 0 2936 0 -1 370
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1713453518
transform 1 0 2928 0 -1 370
box -8 -3 16 105
use FILL  FILL_5265
timestamp 1713453518
transform 1 0 2920 0 -1 370
box -8 -3 16 105
use FILL  FILL_5266
timestamp 1713453518
transform 1 0 2912 0 -1 370
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1713453518
transform 1 0 2904 0 -1 370
box -8 -3 16 105
use FILL  FILL_5268
timestamp 1713453518
transform 1 0 2800 0 -1 370
box -8 -3 16 105
use FILL  FILL_5269
timestamp 1713453518
transform 1 0 2792 0 -1 370
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1713453518
transform 1 0 2784 0 -1 370
box -8 -3 16 105
use FILL  FILL_5271
timestamp 1713453518
transform 1 0 2744 0 -1 370
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1713453518
transform 1 0 2736 0 -1 370
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1713453518
transform 1 0 2728 0 -1 370
box -8 -3 16 105
use FILL  FILL_5274
timestamp 1713453518
transform 1 0 2624 0 -1 370
box -8 -3 16 105
use FILL  FILL_5275
timestamp 1713453518
transform 1 0 2584 0 -1 370
box -8 -3 16 105
use FILL  FILL_5276
timestamp 1713453518
transform 1 0 2576 0 -1 370
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1713453518
transform 1 0 2472 0 -1 370
box -8 -3 16 105
use FILL  FILL_5278
timestamp 1713453518
transform 1 0 2464 0 -1 370
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1713453518
transform 1 0 2368 0 -1 370
box -8 -3 16 105
use FILL  FILL_5280
timestamp 1713453518
transform 1 0 2360 0 -1 370
box -8 -3 16 105
use FILL  FILL_5281
timestamp 1713453518
transform 1 0 2296 0 -1 370
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1713453518
transform 1 0 2288 0 -1 370
box -8 -3 16 105
use FILL  FILL_5283
timestamp 1713453518
transform 1 0 2208 0 -1 370
box -8 -3 16 105
use FILL  FILL_5284
timestamp 1713453518
transform 1 0 2104 0 -1 370
box -8 -3 16 105
use FILL  FILL_5285
timestamp 1713453518
transform 1 0 2096 0 -1 370
box -8 -3 16 105
use FILL  FILL_5286
timestamp 1713453518
transform 1 0 2024 0 -1 370
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1713453518
transform 1 0 2016 0 -1 370
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1713453518
transform 1 0 2008 0 -1 370
box -8 -3 16 105
use FILL  FILL_5289
timestamp 1713453518
transform 1 0 1904 0 -1 370
box -8 -3 16 105
use FILL  FILL_5290
timestamp 1713453518
transform 1 0 1896 0 -1 370
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1713453518
transform 1 0 1888 0 -1 370
box -8 -3 16 105
use FILL  FILL_5292
timestamp 1713453518
transform 1 0 1784 0 -1 370
box -8 -3 16 105
use FILL  FILL_5293
timestamp 1713453518
transform 1 0 1776 0 -1 370
box -8 -3 16 105
use FILL  FILL_5294
timestamp 1713453518
transform 1 0 1672 0 -1 370
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1713453518
transform 1 0 1664 0 -1 370
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1713453518
transform 1 0 1560 0 -1 370
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1713453518
transform 1 0 1552 0 -1 370
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1713453518
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_5299
timestamp 1713453518
transform 1 0 1536 0 -1 370
box -8 -3 16 105
use FILL  FILL_5300
timestamp 1713453518
transform 1 0 1440 0 -1 370
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1713453518
transform 1 0 1432 0 -1 370
box -8 -3 16 105
use FILL  FILL_5302
timestamp 1713453518
transform 1 0 1424 0 -1 370
box -8 -3 16 105
use FILL  FILL_5303
timestamp 1713453518
transform 1 0 1416 0 -1 370
box -8 -3 16 105
use FILL  FILL_5304
timestamp 1713453518
transform 1 0 1312 0 -1 370
box -8 -3 16 105
use FILL  FILL_5305
timestamp 1713453518
transform 1 0 1304 0 -1 370
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1713453518
transform 1 0 1296 0 -1 370
box -8 -3 16 105
use FILL  FILL_5307
timestamp 1713453518
transform 1 0 1288 0 -1 370
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1713453518
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_5309
timestamp 1713453518
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1713453518
transform 1 0 1160 0 -1 370
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1713453518
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1713453518
transform 1 0 1144 0 -1 370
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1713453518
transform 1 0 1040 0 -1 370
box -8 -3 16 105
use FILL  FILL_5314
timestamp 1713453518
transform 1 0 1032 0 -1 370
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1713453518
transform 1 0 1024 0 -1 370
box -8 -3 16 105
use FILL  FILL_5316
timestamp 1713453518
transform 1 0 1016 0 -1 370
box -8 -3 16 105
use FILL  FILL_5317
timestamp 1713453518
transform 1 0 952 0 -1 370
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1713453518
transform 1 0 944 0 -1 370
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1713453518
transform 1 0 936 0 -1 370
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1713453518
transform 1 0 928 0 -1 370
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1713453518
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1713453518
transform 1 0 840 0 -1 370
box -8 -3 16 105
use FILL  FILL_5323
timestamp 1713453518
transform 1 0 832 0 -1 370
box -8 -3 16 105
use FILL  FILL_5324
timestamp 1713453518
transform 1 0 824 0 -1 370
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1713453518
transform 1 0 776 0 -1 370
box -8 -3 16 105
use FILL  FILL_5326
timestamp 1713453518
transform 1 0 768 0 -1 370
box -8 -3 16 105
use FILL  FILL_5327
timestamp 1713453518
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_5328
timestamp 1713453518
transform 1 0 712 0 -1 370
box -8 -3 16 105
use FILL  FILL_5329
timestamp 1713453518
transform 1 0 704 0 -1 370
box -8 -3 16 105
use FILL  FILL_5330
timestamp 1713453518
transform 1 0 632 0 -1 370
box -8 -3 16 105
use FILL  FILL_5331
timestamp 1713453518
transform 1 0 624 0 -1 370
box -8 -3 16 105
use FILL  FILL_5332
timestamp 1713453518
transform 1 0 616 0 -1 370
box -8 -3 16 105
use FILL  FILL_5333
timestamp 1713453518
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_5334
timestamp 1713453518
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_5335
timestamp 1713453518
transform 1 0 528 0 -1 370
box -8 -3 16 105
use FILL  FILL_5336
timestamp 1713453518
transform 1 0 520 0 -1 370
box -8 -3 16 105
use FILL  FILL_5337
timestamp 1713453518
transform 1 0 512 0 -1 370
box -8 -3 16 105
use FILL  FILL_5338
timestamp 1713453518
transform 1 0 504 0 -1 370
box -8 -3 16 105
use FILL  FILL_5339
timestamp 1713453518
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_5340
timestamp 1713453518
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_5341
timestamp 1713453518
transform 1 0 456 0 -1 370
box -8 -3 16 105
use FILL  FILL_5342
timestamp 1713453518
transform 1 0 416 0 -1 370
box -8 -3 16 105
use FILL  FILL_5343
timestamp 1713453518
transform 1 0 408 0 -1 370
box -8 -3 16 105
use FILL  FILL_5344
timestamp 1713453518
transform 1 0 376 0 -1 370
box -8 -3 16 105
use FILL  FILL_5345
timestamp 1713453518
transform 1 0 368 0 -1 370
box -8 -3 16 105
use FILL  FILL_5346
timestamp 1713453518
transform 1 0 320 0 -1 370
box -8 -3 16 105
use FILL  FILL_5347
timestamp 1713453518
transform 1 0 312 0 -1 370
box -8 -3 16 105
use FILL  FILL_5348
timestamp 1713453518
transform 1 0 304 0 -1 370
box -8 -3 16 105
use FILL  FILL_5349
timestamp 1713453518
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_5350
timestamp 1713453518
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_5351
timestamp 1713453518
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_5352
timestamp 1713453518
transform 1 0 176 0 -1 370
box -8 -3 16 105
use FILL  FILL_5353
timestamp 1713453518
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_5354
timestamp 1713453518
transform 1 0 3440 0 1 170
box -8 -3 16 105
use FILL  FILL_5355
timestamp 1713453518
transform 1 0 3432 0 1 170
box -8 -3 16 105
use FILL  FILL_5356
timestamp 1713453518
transform 1 0 3424 0 1 170
box -8 -3 16 105
use FILL  FILL_5357
timestamp 1713453518
transform 1 0 3416 0 1 170
box -8 -3 16 105
use FILL  FILL_5358
timestamp 1713453518
transform 1 0 3408 0 1 170
box -8 -3 16 105
use FILL  FILL_5359
timestamp 1713453518
transform 1 0 3400 0 1 170
box -8 -3 16 105
use FILL  FILL_5360
timestamp 1713453518
transform 1 0 3392 0 1 170
box -8 -3 16 105
use FILL  FILL_5361
timestamp 1713453518
transform 1 0 3384 0 1 170
box -8 -3 16 105
use FILL  FILL_5362
timestamp 1713453518
transform 1 0 3376 0 1 170
box -8 -3 16 105
use FILL  FILL_5363
timestamp 1713453518
transform 1 0 3272 0 1 170
box -8 -3 16 105
use FILL  FILL_5364
timestamp 1713453518
transform 1 0 3264 0 1 170
box -8 -3 16 105
use FILL  FILL_5365
timestamp 1713453518
transform 1 0 3256 0 1 170
box -8 -3 16 105
use FILL  FILL_5366
timestamp 1713453518
transform 1 0 3248 0 1 170
box -8 -3 16 105
use FILL  FILL_5367
timestamp 1713453518
transform 1 0 3184 0 1 170
box -8 -3 16 105
use FILL  FILL_5368
timestamp 1713453518
transform 1 0 3176 0 1 170
box -8 -3 16 105
use FILL  FILL_5369
timestamp 1713453518
transform 1 0 3168 0 1 170
box -8 -3 16 105
use FILL  FILL_5370
timestamp 1713453518
transform 1 0 3160 0 1 170
box -8 -3 16 105
use FILL  FILL_5371
timestamp 1713453518
transform 1 0 3152 0 1 170
box -8 -3 16 105
use FILL  FILL_5372
timestamp 1713453518
transform 1 0 3144 0 1 170
box -8 -3 16 105
use FILL  FILL_5373
timestamp 1713453518
transform 1 0 3104 0 1 170
box -8 -3 16 105
use FILL  FILL_5374
timestamp 1713453518
transform 1 0 3096 0 1 170
box -8 -3 16 105
use FILL  FILL_5375
timestamp 1713453518
transform 1 0 3088 0 1 170
box -8 -3 16 105
use FILL  FILL_5376
timestamp 1713453518
transform 1 0 3080 0 1 170
box -8 -3 16 105
use FILL  FILL_5377
timestamp 1713453518
transform 1 0 3024 0 1 170
box -8 -3 16 105
use FILL  FILL_5378
timestamp 1713453518
transform 1 0 3016 0 1 170
box -8 -3 16 105
use FILL  FILL_5379
timestamp 1713453518
transform 1 0 3008 0 1 170
box -8 -3 16 105
use FILL  FILL_5380
timestamp 1713453518
transform 1 0 2968 0 1 170
box -8 -3 16 105
use FILL  FILL_5381
timestamp 1713453518
transform 1 0 2936 0 1 170
box -8 -3 16 105
use FILL  FILL_5382
timestamp 1713453518
transform 1 0 2928 0 1 170
box -8 -3 16 105
use FILL  FILL_5383
timestamp 1713453518
transform 1 0 2920 0 1 170
box -8 -3 16 105
use FILL  FILL_5384
timestamp 1713453518
transform 1 0 2872 0 1 170
box -8 -3 16 105
use FILL  FILL_5385
timestamp 1713453518
transform 1 0 2864 0 1 170
box -8 -3 16 105
use FILL  FILL_5386
timestamp 1713453518
transform 1 0 2856 0 1 170
box -8 -3 16 105
use FILL  FILL_5387
timestamp 1713453518
transform 1 0 2792 0 1 170
box -8 -3 16 105
use FILL  FILL_5388
timestamp 1713453518
transform 1 0 2784 0 1 170
box -8 -3 16 105
use FILL  FILL_5389
timestamp 1713453518
transform 1 0 2776 0 1 170
box -8 -3 16 105
use FILL  FILL_5390
timestamp 1713453518
transform 1 0 2768 0 1 170
box -8 -3 16 105
use FILL  FILL_5391
timestamp 1713453518
transform 1 0 2704 0 1 170
box -8 -3 16 105
use FILL  FILL_5392
timestamp 1713453518
transform 1 0 2696 0 1 170
box -8 -3 16 105
use FILL  FILL_5393
timestamp 1713453518
transform 1 0 2656 0 1 170
box -8 -3 16 105
use FILL  FILL_5394
timestamp 1713453518
transform 1 0 2648 0 1 170
box -8 -3 16 105
use FILL  FILL_5395
timestamp 1713453518
transform 1 0 2640 0 1 170
box -8 -3 16 105
use FILL  FILL_5396
timestamp 1713453518
transform 1 0 2632 0 1 170
box -8 -3 16 105
use FILL  FILL_5397
timestamp 1713453518
transform 1 0 2584 0 1 170
box -8 -3 16 105
use FILL  FILL_5398
timestamp 1713453518
transform 1 0 2560 0 1 170
box -8 -3 16 105
use FILL  FILL_5399
timestamp 1713453518
transform 1 0 2552 0 1 170
box -8 -3 16 105
use FILL  FILL_5400
timestamp 1713453518
transform 1 0 2544 0 1 170
box -8 -3 16 105
use FILL  FILL_5401
timestamp 1713453518
transform 1 0 2480 0 1 170
box -8 -3 16 105
use FILL  FILL_5402
timestamp 1713453518
transform 1 0 2472 0 1 170
box -8 -3 16 105
use FILL  FILL_5403
timestamp 1713453518
transform 1 0 2464 0 1 170
box -8 -3 16 105
use FILL  FILL_5404
timestamp 1713453518
transform 1 0 2408 0 1 170
box -8 -3 16 105
use FILL  FILL_5405
timestamp 1713453518
transform 1 0 2400 0 1 170
box -8 -3 16 105
use FILL  FILL_5406
timestamp 1713453518
transform 1 0 2392 0 1 170
box -8 -3 16 105
use FILL  FILL_5407
timestamp 1713453518
transform 1 0 2384 0 1 170
box -8 -3 16 105
use FILL  FILL_5408
timestamp 1713453518
transform 1 0 2344 0 1 170
box -8 -3 16 105
use FILL  FILL_5409
timestamp 1713453518
transform 1 0 2304 0 1 170
box -8 -3 16 105
use FILL  FILL_5410
timestamp 1713453518
transform 1 0 2296 0 1 170
box -8 -3 16 105
use FILL  FILL_5411
timestamp 1713453518
transform 1 0 2288 0 1 170
box -8 -3 16 105
use FILL  FILL_5412
timestamp 1713453518
transform 1 0 2280 0 1 170
box -8 -3 16 105
use FILL  FILL_5413
timestamp 1713453518
transform 1 0 2272 0 1 170
box -8 -3 16 105
use FILL  FILL_5414
timestamp 1713453518
transform 1 0 2208 0 1 170
box -8 -3 16 105
use FILL  FILL_5415
timestamp 1713453518
transform 1 0 2200 0 1 170
box -8 -3 16 105
use FILL  FILL_5416
timestamp 1713453518
transform 1 0 2192 0 1 170
box -8 -3 16 105
use FILL  FILL_5417
timestamp 1713453518
transform 1 0 2184 0 1 170
box -8 -3 16 105
use FILL  FILL_5418
timestamp 1713453518
transform 1 0 2176 0 1 170
box -8 -3 16 105
use FILL  FILL_5419
timestamp 1713453518
transform 1 0 2112 0 1 170
box -8 -3 16 105
use FILL  FILL_5420
timestamp 1713453518
transform 1 0 2104 0 1 170
box -8 -3 16 105
use FILL  FILL_5421
timestamp 1713453518
transform 1 0 2096 0 1 170
box -8 -3 16 105
use FILL  FILL_5422
timestamp 1713453518
transform 1 0 2088 0 1 170
box -8 -3 16 105
use FILL  FILL_5423
timestamp 1713453518
transform 1 0 2080 0 1 170
box -8 -3 16 105
use FILL  FILL_5424
timestamp 1713453518
transform 1 0 2024 0 1 170
box -8 -3 16 105
use FILL  FILL_5425
timestamp 1713453518
transform 1 0 1992 0 1 170
box -8 -3 16 105
use FILL  FILL_5426
timestamp 1713453518
transform 1 0 1984 0 1 170
box -8 -3 16 105
use FILL  FILL_5427
timestamp 1713453518
transform 1 0 1976 0 1 170
box -8 -3 16 105
use FILL  FILL_5428
timestamp 1713453518
transform 1 0 1928 0 1 170
box -8 -3 16 105
use FILL  FILL_5429
timestamp 1713453518
transform 1 0 1920 0 1 170
box -8 -3 16 105
use FILL  FILL_5430
timestamp 1713453518
transform 1 0 1912 0 1 170
box -8 -3 16 105
use FILL  FILL_5431
timestamp 1713453518
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_5432
timestamp 1713453518
transform 1 0 1856 0 1 170
box -8 -3 16 105
use FILL  FILL_5433
timestamp 1713453518
transform 1 0 1848 0 1 170
box -8 -3 16 105
use FILL  FILL_5434
timestamp 1713453518
transform 1 0 1840 0 1 170
box -8 -3 16 105
use FILL  FILL_5435
timestamp 1713453518
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_5436
timestamp 1713453518
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_5437
timestamp 1713453518
transform 1 0 1816 0 1 170
box -8 -3 16 105
use FILL  FILL_5438
timestamp 1713453518
transform 1 0 1808 0 1 170
box -8 -3 16 105
use FILL  FILL_5439
timestamp 1713453518
transform 1 0 1800 0 1 170
box -8 -3 16 105
use FILL  FILL_5440
timestamp 1713453518
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_5441
timestamp 1713453518
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_5442
timestamp 1713453518
transform 1 0 1680 0 1 170
box -8 -3 16 105
use FILL  FILL_5443
timestamp 1713453518
transform 1 0 1672 0 1 170
box -8 -3 16 105
use FILL  FILL_5444
timestamp 1713453518
transform 1 0 1664 0 1 170
box -8 -3 16 105
use FILL  FILL_5445
timestamp 1713453518
transform 1 0 1656 0 1 170
box -8 -3 16 105
use FILL  FILL_5446
timestamp 1713453518
transform 1 0 1600 0 1 170
box -8 -3 16 105
use FILL  FILL_5447
timestamp 1713453518
transform 1 0 1592 0 1 170
box -8 -3 16 105
use FILL  FILL_5448
timestamp 1713453518
transform 1 0 1584 0 1 170
box -8 -3 16 105
use FILL  FILL_5449
timestamp 1713453518
transform 1 0 1560 0 1 170
box -8 -3 16 105
use FILL  FILL_5450
timestamp 1713453518
transform 1 0 1552 0 1 170
box -8 -3 16 105
use FILL  FILL_5451
timestamp 1713453518
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_5452
timestamp 1713453518
transform 1 0 1480 0 1 170
box -8 -3 16 105
use FILL  FILL_5453
timestamp 1713453518
transform 1 0 1472 0 1 170
box -8 -3 16 105
use FILL  FILL_5454
timestamp 1713453518
transform 1 0 1464 0 1 170
box -8 -3 16 105
use FILL  FILL_5455
timestamp 1713453518
transform 1 0 1456 0 1 170
box -8 -3 16 105
use FILL  FILL_5456
timestamp 1713453518
transform 1 0 1448 0 1 170
box -8 -3 16 105
use FILL  FILL_5457
timestamp 1713453518
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_5458
timestamp 1713453518
transform 1 0 1376 0 1 170
box -8 -3 16 105
use FILL  FILL_5459
timestamp 1713453518
transform 1 0 1344 0 1 170
box -8 -3 16 105
use FILL  FILL_5460
timestamp 1713453518
transform 1 0 1336 0 1 170
box -8 -3 16 105
use FILL  FILL_5461
timestamp 1713453518
transform 1 0 1328 0 1 170
box -8 -3 16 105
use FILL  FILL_5462
timestamp 1713453518
transform 1 0 1320 0 1 170
box -8 -3 16 105
use FILL  FILL_5463
timestamp 1713453518
transform 1 0 1280 0 1 170
box -8 -3 16 105
use FILL  FILL_5464
timestamp 1713453518
transform 1 0 1272 0 1 170
box -8 -3 16 105
use FILL  FILL_5465
timestamp 1713453518
transform 1 0 1224 0 1 170
box -8 -3 16 105
use FILL  FILL_5466
timestamp 1713453518
transform 1 0 1216 0 1 170
box -8 -3 16 105
use FILL  FILL_5467
timestamp 1713453518
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_5468
timestamp 1713453518
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_5469
timestamp 1713453518
transform 1 0 1096 0 1 170
box -8 -3 16 105
use FILL  FILL_5470
timestamp 1713453518
transform 1 0 1088 0 1 170
box -8 -3 16 105
use FILL  FILL_5471
timestamp 1713453518
transform 1 0 1048 0 1 170
box -8 -3 16 105
use FILL  FILL_5472
timestamp 1713453518
transform 1 0 1040 0 1 170
box -8 -3 16 105
use FILL  FILL_5473
timestamp 1713453518
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_5474
timestamp 1713453518
transform 1 0 928 0 1 170
box -8 -3 16 105
use FILL  FILL_5475
timestamp 1713453518
transform 1 0 920 0 1 170
box -8 -3 16 105
use FILL  FILL_5476
timestamp 1713453518
transform 1 0 912 0 1 170
box -8 -3 16 105
use FILL  FILL_5477
timestamp 1713453518
transform 1 0 840 0 1 170
box -8 -3 16 105
use FILL  FILL_5478
timestamp 1713453518
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_5479
timestamp 1713453518
transform 1 0 800 0 1 170
box -8 -3 16 105
use FILL  FILL_5480
timestamp 1713453518
transform 1 0 792 0 1 170
box -8 -3 16 105
use FILL  FILL_5481
timestamp 1713453518
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_5482
timestamp 1713453518
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_5483
timestamp 1713453518
transform 1 0 768 0 1 170
box -8 -3 16 105
use FILL  FILL_5484
timestamp 1713453518
transform 1 0 696 0 1 170
box -8 -3 16 105
use FILL  FILL_5485
timestamp 1713453518
transform 1 0 688 0 1 170
box -8 -3 16 105
use FILL  FILL_5486
timestamp 1713453518
transform 1 0 680 0 1 170
box -8 -3 16 105
use FILL  FILL_5487
timestamp 1713453518
transform 1 0 672 0 1 170
box -8 -3 16 105
use FILL  FILL_5488
timestamp 1713453518
transform 1 0 568 0 1 170
box -8 -3 16 105
use FILL  FILL_5489
timestamp 1713453518
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_5490
timestamp 1713453518
transform 1 0 552 0 1 170
box -8 -3 16 105
use FILL  FILL_5491
timestamp 1713453518
transform 1 0 448 0 1 170
box -8 -3 16 105
use FILL  FILL_5492
timestamp 1713453518
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_5493
timestamp 1713453518
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_5494
timestamp 1713453518
transform 1 0 424 0 1 170
box -8 -3 16 105
use FILL  FILL_5495
timestamp 1713453518
transform 1 0 360 0 1 170
box -8 -3 16 105
use FILL  FILL_5496
timestamp 1713453518
transform 1 0 352 0 1 170
box -8 -3 16 105
use FILL  FILL_5497
timestamp 1713453518
transform 1 0 344 0 1 170
box -8 -3 16 105
use FILL  FILL_5498
timestamp 1713453518
transform 1 0 240 0 1 170
box -8 -3 16 105
use FILL  FILL_5499
timestamp 1713453518
transform 1 0 232 0 1 170
box -8 -3 16 105
use FILL  FILL_5500
timestamp 1713453518
transform 1 0 224 0 1 170
box -8 -3 16 105
use FILL  FILL_5501
timestamp 1713453518
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_5502
timestamp 1713453518
transform 1 0 112 0 1 170
box -8 -3 16 105
use FILL  FILL_5503
timestamp 1713453518
transform 1 0 104 0 1 170
box -8 -3 16 105
use FILL  FILL_5504
timestamp 1713453518
transform 1 0 96 0 1 170
box -8 -3 16 105
use FILL  FILL_5505
timestamp 1713453518
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_5506
timestamp 1713453518
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_5507
timestamp 1713453518
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_5508
timestamp 1713453518
transform 1 0 3248 0 -1 170
box -8 -3 16 105
use FILL  FILL_5509
timestamp 1713453518
transform 1 0 3144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5510
timestamp 1713453518
transform 1 0 3136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5511
timestamp 1713453518
transform 1 0 3056 0 -1 170
box -8 -3 16 105
use FILL  FILL_5512
timestamp 1713453518
transform 1 0 3048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5513
timestamp 1713453518
transform 1 0 3000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5514
timestamp 1713453518
transform 1 0 2936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5515
timestamp 1713453518
transform 1 0 2872 0 -1 170
box -8 -3 16 105
use FILL  FILL_5516
timestamp 1713453518
transform 1 0 2784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5517
timestamp 1713453518
transform 1 0 2776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5518
timestamp 1713453518
transform 1 0 2768 0 -1 170
box -8 -3 16 105
use FILL  FILL_5519
timestamp 1713453518
transform 1 0 2688 0 -1 170
box -8 -3 16 105
use FILL  FILL_5520
timestamp 1713453518
transform 1 0 2680 0 -1 170
box -8 -3 16 105
use FILL  FILL_5521
timestamp 1713453518
transform 1 0 2656 0 -1 170
box -8 -3 16 105
use FILL  FILL_5522
timestamp 1713453518
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_5523
timestamp 1713453518
transform 1 0 2560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5524
timestamp 1713453518
transform 1 0 2552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5525
timestamp 1713453518
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5526
timestamp 1713453518
transform 1 0 2440 0 -1 170
box -8 -3 16 105
use FILL  FILL_5527
timestamp 1713453518
transform 1 0 2336 0 -1 170
box -8 -3 16 105
use FILL  FILL_5528
timestamp 1713453518
transform 1 0 2328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5529
timestamp 1713453518
transform 1 0 2224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5530
timestamp 1713453518
transform 1 0 2216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5531
timestamp 1713453518
transform 1 0 2192 0 -1 170
box -8 -3 16 105
use FILL  FILL_5532
timestamp 1713453518
transform 1 0 2112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5533
timestamp 1713453518
transform 1 0 2104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5534
timestamp 1713453518
transform 1 0 2064 0 -1 170
box -8 -3 16 105
use FILL  FILL_5535
timestamp 1713453518
transform 1 0 2000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5536
timestamp 1713453518
transform 1 0 1992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5537
timestamp 1713453518
transform 1 0 1944 0 -1 170
box -8 -3 16 105
use FILL  FILL_5538
timestamp 1713453518
transform 1 0 1840 0 -1 170
box -8 -3 16 105
use FILL  FILL_5539
timestamp 1713453518
transform 1 0 1832 0 -1 170
box -8 -3 16 105
use FILL  FILL_5540
timestamp 1713453518
transform 1 0 1744 0 -1 170
box -8 -3 16 105
use FILL  FILL_5541
timestamp 1713453518
transform 1 0 1736 0 -1 170
box -8 -3 16 105
use FILL  FILL_5542
timestamp 1713453518
transform 1 0 1672 0 -1 170
box -8 -3 16 105
use FILL  FILL_5543
timestamp 1713453518
transform 1 0 1568 0 -1 170
box -8 -3 16 105
use FILL  FILL_5544
timestamp 1713453518
transform 1 0 1560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5545
timestamp 1713453518
transform 1 0 1552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5546
timestamp 1713453518
transform 1 0 1544 0 -1 170
box -8 -3 16 105
use FILL  FILL_5547
timestamp 1713453518
transform 1 0 1456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5548
timestamp 1713453518
transform 1 0 1448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5549
timestamp 1713453518
transform 1 0 1440 0 -1 170
box -8 -3 16 105
use FILL  FILL_5550
timestamp 1713453518
transform 1 0 1432 0 -1 170
box -8 -3 16 105
use FILL  FILL_5551
timestamp 1713453518
transform 1 0 1376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5552
timestamp 1713453518
transform 1 0 1320 0 -1 170
box -8 -3 16 105
use FILL  FILL_5553
timestamp 1713453518
transform 1 0 1312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5554
timestamp 1713453518
transform 1 0 1304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5555
timestamp 1713453518
transform 1 0 1296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5556
timestamp 1713453518
transform 1 0 1208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5557
timestamp 1713453518
transform 1 0 1200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5558
timestamp 1713453518
transform 1 0 1192 0 -1 170
box -8 -3 16 105
use FILL  FILL_5559
timestamp 1713453518
transform 1 0 1088 0 -1 170
box -8 -3 16 105
use FILL  FILL_5560
timestamp 1713453518
transform 1 0 1048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5561
timestamp 1713453518
transform 1 0 944 0 -1 170
box -8 -3 16 105
use FILL  FILL_5562
timestamp 1713453518
transform 1 0 936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5563
timestamp 1713453518
transform 1 0 832 0 -1 170
box -8 -3 16 105
use FILL  FILL_5564
timestamp 1713453518
transform 1 0 728 0 -1 170
box -8 -3 16 105
use FILL  FILL_5565
timestamp 1713453518
transform 1 0 720 0 -1 170
box -8 -3 16 105
use FILL  FILL_5566
timestamp 1713453518
transform 1 0 616 0 -1 170
box -8 -3 16 105
use FILL  FILL_5567
timestamp 1713453518
transform 1 0 608 0 -1 170
box -8 -3 16 105
use FILL  FILL_5568
timestamp 1713453518
transform 1 0 504 0 -1 170
box -8 -3 16 105
use FILL  FILL_5569
timestamp 1713453518
transform 1 0 496 0 -1 170
box -8 -3 16 105
use FILL  FILL_5570
timestamp 1713453518
transform 1 0 488 0 -1 170
box -8 -3 16 105
use FILL  FILL_5571
timestamp 1713453518
transform 1 0 480 0 -1 170
box -8 -3 16 105
use FILL  FILL_5572
timestamp 1713453518
transform 1 0 368 0 -1 170
box -8 -3 16 105
use FILL  FILL_5573
timestamp 1713453518
transform 1 0 360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5574
timestamp 1713453518
transform 1 0 352 0 -1 170
box -8 -3 16 105
use FILL  FILL_5575
timestamp 1713453518
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_5576
timestamp 1713453518
transform 1 0 240 0 -1 170
box -8 -3 16 105
use FILL  FILL_5577
timestamp 1713453518
transform 1 0 232 0 -1 170
box -8 -3 16 105
use FILL  FILL_5578
timestamp 1713453518
transform 1 0 192 0 -1 170
box -8 -3 16 105
use FILL  FILL_5579
timestamp 1713453518
transform 1 0 184 0 -1 170
box -8 -3 16 105
use FILL  FILL_5580
timestamp 1713453518
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_5581
timestamp 1713453518
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1713453518
transform 1 0 2792 0 -1 170
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1713453518
transform 1 0 2576 0 -1 170
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1713453518
transform 1 0 2472 0 -1 170
box -5 -3 84 105
use INVX2  INVX2_0
timestamp 1713453518
transform 1 0 2376 0 1 370
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1713453518
transform 1 0 1840 0 1 570
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1713453518
transform 1 0 2192 0 1 370
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1713453518
transform 1 0 2424 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1713453518
transform 1 0 1560 0 1 370
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1713453518
transform 1 0 1336 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1713453518
transform 1 0 1240 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1713453518
transform 1 0 3336 0 1 370
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1713453518
transform 1 0 3304 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1713453518
transform 1 0 3416 0 1 570
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1713453518
transform 1 0 3128 0 1 370
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1713453518
transform 1 0 3392 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1713453518
transform 1 0 1152 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1713453518
transform 1 0 1112 0 1 370
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1713453518
transform 1 0 1288 0 1 370
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1713453518
transform 1 0 1112 0 1 770
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1713453518
transform 1 0 1312 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1713453518
transform 1 0 1600 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1713453518
transform 1 0 1528 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1713453518
transform 1 0 1464 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1713453518
transform 1 0 1184 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1713453518
transform 1 0 1576 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1713453518
transform 1 0 1448 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1713453518
transform 1 0 1200 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1713453518
transform 1 0 1088 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1713453518
transform 1 0 1168 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1713453518
transform 1 0 1552 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1713453518
transform 1 0 1600 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1713453518
transform 1 0 1152 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1713453518
transform 1 0 1120 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1713453518
transform 1 0 1168 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1713453518
transform 1 0 1424 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1713453518
transform 1 0 1312 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1713453518
transform 1 0 1376 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1713453518
transform 1 0 1200 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1713453518
transform 1 0 1672 0 1 370
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1713453518
transform 1 0 1152 0 1 570
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1713453518
transform 1 0 1376 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1713453518
transform 1 0 1584 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1713453518
transform 1 0 1600 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1713453518
transform 1 0 1096 0 1 970
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1713453518
transform 1 0 1168 0 1 570
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1713453518
transform 1 0 1136 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1713453518
transform 1 0 1344 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1713453518
transform 1 0 1440 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1713453518
transform 1 0 1432 0 1 970
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1713453518
transform 1 0 1640 0 1 370
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1713453518
transform 1 0 1168 0 1 770
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1713453518
transform 1 0 1368 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1713453518
transform 1 0 1472 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1713453518
transform 1 0 1512 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1713453518
transform 1 0 1360 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1713453518
transform 1 0 1600 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1713453518
transform 1 0 1184 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1713453518
transform 1 0 1448 0 1 570
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1713453518
transform 1 0 1192 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1713453518
transform 1 0 1472 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1713453518
transform 1 0 1360 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1713453518
transform 1 0 1448 0 1 970
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1713453518
transform 1 0 2448 0 1 170
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1713453518
transform 1 0 3080 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1713453518
transform 1 0 3064 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1713453518
transform 1 0 3312 0 1 570
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1713453518
transform 1 0 3296 0 1 570
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1713453518
transform 1 0 3328 0 1 770
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1713453518
transform 1 0 3008 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1713453518
transform 1 0 2728 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1713453518
transform 1 0 2768 0 1 770
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1713453518
transform 1 0 3416 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1713453518
transform 1 0 2992 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1713453518
transform 1 0 3288 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1713453518
transform 1 0 3384 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1713453518
transform 1 0 2744 0 1 770
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1713453518
transform 1 0 3248 0 1 570
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1713453518
transform 1 0 2632 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1713453518
transform 1 0 2912 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1713453518
transform 1 0 3168 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1713453518
transform 1 0 2952 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1713453518
transform 1 0 3000 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1713453518
transform 1 0 3344 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1713453518
transform 1 0 3280 0 1 770
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1713453518
transform 1 0 1792 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1713453518
transform 1 0 1792 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1713453518
transform 1 0 2776 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1713453518
transform 1 0 3248 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1713453518
transform 1 0 3208 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1713453518
transform 1 0 2752 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1713453518
transform 1 0 2584 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1713453518
transform 1 0 3336 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1713453518
transform 1 0 2264 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1713453518
transform 1 0 2216 0 1 770
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1713453518
transform 1 0 2560 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1713453518
transform 1 0 3400 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1713453518
transform 1 0 3176 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1713453518
transform 1 0 3256 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1713453518
transform 1 0 3312 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1713453518
transform 1 0 2688 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1713453518
transform 1 0 2688 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1713453518
transform 1 0 3232 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1713453518
transform 1 0 2528 0 1 570
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1713453518
transform 1 0 3232 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1713453518
transform 1 0 1864 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1713453518
transform 1 0 2936 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1713453518
transform 1 0 2608 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1713453518
transform 1 0 2648 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1713453518
transform 1 0 2952 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1713453518
transform 1 0 2952 0 1 770
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1713453518
transform 1 0 2920 0 1 970
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1713453518
transform 1 0 2816 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1713453518
transform 1 0 2232 0 1 770
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1713453518
transform 1 0 3016 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1713453518
transform 1 0 3416 0 1 770
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1713453518
transform 1 0 2448 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1713453518
transform 1 0 3272 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1713453518
transform 1 0 3024 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1713453518
transform 1 0 2616 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1713453518
transform 1 0 2784 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1713453518
transform 1 0 2232 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1713453518
transform 1 0 2544 0 1 570
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1713453518
transform 1 0 192 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1713453518
transform 1 0 136 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1713453518
transform 1 0 184 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1713453518
transform 1 0 232 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1713453518
transform 1 0 424 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1713453518
transform 1 0 608 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1713453518
transform 1 0 624 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1713453518
transform 1 0 208 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1713453518
transform 1 0 248 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1713453518
transform 1 0 248 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1713453518
transform 1 0 200 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1713453518
transform 1 0 184 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1713453518
transform 1 0 376 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1713453518
transform 1 0 208 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1713453518
transform 1 0 216 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1713453518
transform 1 0 216 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1713453518
transform 1 0 208 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1713453518
transform 1 0 208 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1713453518
transform 1 0 312 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1713453518
transform 1 0 328 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1713453518
transform 1 0 128 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1713453518
transform 1 0 192 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1713453518
transform 1 0 216 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1713453518
transform 1 0 192 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1713453518
transform 1 0 208 0 1 970
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1713453518
transform 1 0 80 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1713453518
transform 1 0 200 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1713453518
transform 1 0 96 0 1 970
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1713453518
transform 1 0 416 0 1 570
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1713453518
transform 1 0 280 0 1 370
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1713453518
transform 1 0 312 0 1 770
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1713453518
transform 1 0 760 0 1 370
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1713453518
transform 1 0 856 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1713453518
transform 1 0 840 0 1 370
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1713453518
transform 1 0 1328 0 1 370
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1713453518
transform 1 0 912 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1713453518
transform 1 0 2376 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1713453518
transform 1 0 2256 0 1 170
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1713453518
transform 1 0 2032 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1713453518
transform 1 0 3064 0 1 170
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1713453518
transform 1 0 2944 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1713453518
transform 1 0 2432 0 1 170
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1713453518
transform 1 0 1640 0 1 170
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1713453518
transform 1 0 1488 0 1 170
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1713453518
transform 1 0 2416 0 1 170
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1713453518
transform 1 0 2568 0 1 170
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1713453518
transform 1 0 352 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1713453518
transform 1 0 2648 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1713453518
transform 1 0 720 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1713453518
transform 1 0 2616 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1713453518
transform 1 0 2776 0 1 970
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1713453518
transform 1 0 3088 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1713453518
transform 1 0 632 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1713453518
transform 1 0 2480 0 1 970
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1713453518
transform 1 0 2912 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1713453518
transform 1 0 800 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1713453518
transform 1 0 2104 0 1 970
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1713453518
transform 1 0 2576 0 1 770
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1713453518
transform 1 0 744 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1713453518
transform 1 0 2112 0 1 770
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1713453518
transform 1 0 1904 0 1 770
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1713453518
transform 1 0 2520 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1713453518
transform 1 0 936 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1713453518
transform 1 0 2080 0 1 770
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1713453518
transform 1 0 792 0 1 970
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1713453518
transform 1 0 1536 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1713453518
transform 1 0 512 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1713453518
transform 1 0 736 0 1 970
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1713453518
transform 1 0 744 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1713453518
transform 1 0 1280 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1713453518
transform 1 0 1632 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1713453518
transform 1 0 1712 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1713453518
transform 1 0 680 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1713453518
transform 1 0 1408 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1713453518
transform 1 0 1592 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1713453518
transform 1 0 1856 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1713453518
transform 1 0 1704 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1713453518
transform 1 0 752 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1713453518
transform 1 0 848 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1713453518
transform 1 0 1376 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1713453518
transform 1 0 2152 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1713453518
transform 1 0 2048 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1713453518
transform 1 0 440 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1713453518
transform 1 0 2128 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1713453518
transform 1 0 2968 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1713453518
transform 1 0 936 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1713453518
transform 1 0 1144 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1713453518
transform 1 0 2968 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1713453518
transform 1 0 1024 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1713453518
transform 1 0 1192 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1713453518
transform 1 0 2928 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1713453518
transform 1 0 2864 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1713453518
transform 1 0 3272 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1713453518
transform 1 0 1128 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1713453518
transform 1 0 1312 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1713453518
transform 1 0 2672 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1713453518
transform 1 0 3416 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1713453518
transform 1 0 904 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1713453518
transform 1 0 488 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1713453518
transform 1 0 3384 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1713453518
transform 1 0 888 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1713453518
transform 1 0 2208 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1713453518
transform 1 0 2648 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1713453518
transform 1 0 3056 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_223
timestamp 1713453518
transform 1 0 3416 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1713453518
transform 1 0 864 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_225
timestamp 1713453518
transform 1 0 3056 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_226
timestamp 1713453518
transform 1 0 2304 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_227
timestamp 1713453518
transform 1 0 832 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_228
timestamp 1713453518
transform 1 0 1928 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_229
timestamp 1713453518
transform 1 0 456 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_230
timestamp 1713453518
transform 1 0 560 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1713453518
transform 1 0 632 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_232
timestamp 1713453518
transform 1 0 2312 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1713453518
transform 1 0 864 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_234
timestamp 1713453518
transform 1 0 2016 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_235
timestamp 1713453518
transform 1 0 896 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_236
timestamp 1713453518
transform 1 0 2552 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_237
timestamp 1713453518
transform 1 0 3368 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1713453518
transform 1 0 864 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_239
timestamp 1713453518
transform 1 0 2048 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1713453518
transform 1 0 3400 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_241
timestamp 1713453518
transform 1 0 808 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_242
timestamp 1713453518
transform 1 0 1880 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_243
timestamp 1713453518
transform 1 0 824 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_244
timestamp 1713453518
transform 1 0 2136 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_245
timestamp 1713453518
transform 1 0 2920 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1713453518
transform 1 0 2704 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_247
timestamp 1713453518
transform 1 0 2992 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_248
timestamp 1713453518
transform 1 0 624 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_249
timestamp 1713453518
transform 1 0 528 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_250
timestamp 1713453518
transform 1 0 600 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_251
timestamp 1713453518
transform 1 0 2152 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_252
timestamp 1713453518
transform 1 0 2888 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_253
timestamp 1713453518
transform 1 0 3416 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_254
timestamp 1713453518
transform 1 0 560 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_255
timestamp 1713453518
transform 1 0 3408 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_256
timestamp 1713453518
transform 1 0 2440 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_257
timestamp 1713453518
transform 1 0 1040 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_258
timestamp 1713453518
transform 1 0 1952 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_259
timestamp 1713453518
transform 1 0 2728 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_260
timestamp 1713453518
transform 1 0 2552 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_261
timestamp 1713453518
transform 1 0 3096 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_262
timestamp 1713453518
transform 1 0 1096 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_263
timestamp 1713453518
transform 1 0 2640 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_264
timestamp 1713453518
transform 1 0 3256 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_265
timestamp 1713453518
transform 1 0 1064 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_266
timestamp 1713453518
transform 1 0 2600 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_267
timestamp 1713453518
transform 1 0 3024 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_268
timestamp 1713453518
transform 1 0 984 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_269
timestamp 1713453518
transform 1 0 488 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_270
timestamp 1713453518
transform 1 0 528 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_271
timestamp 1713453518
transform 1 0 736 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_272
timestamp 1713453518
transform 1 0 2608 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_273
timestamp 1713453518
transform 1 0 2416 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_274
timestamp 1713453518
transform 1 0 688 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_275
timestamp 1713453518
transform 1 0 584 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_276
timestamp 1713453518
transform 1 0 592 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_277
timestamp 1713453518
transform 1 0 544 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_278
timestamp 1713453518
transform 1 0 672 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_279
timestamp 1713453518
transform 1 0 488 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_280
timestamp 1713453518
transform 1 0 728 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_281
timestamp 1713453518
transform 1 0 1936 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_282
timestamp 1713453518
transform 1 0 448 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_283
timestamp 1713453518
transform 1 0 536 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_284
timestamp 1713453518
transform 1 0 472 0 1 970
box -9 -3 26 105
use INVX2  INVX2_285
timestamp 1713453518
transform 1 0 1752 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_286
timestamp 1713453518
transform 1 0 1952 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_287
timestamp 1713453518
transform 1 0 1768 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_288
timestamp 1713453518
transform 1 0 2048 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_289
timestamp 1713453518
transform 1 0 1880 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_290
timestamp 1713453518
transform 1 0 2064 0 1 170
box -9 -3 26 105
use INVX2  INVX2_291
timestamp 1713453518
transform 1 0 1896 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_292
timestamp 1713453518
transform 1 0 2200 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_293
timestamp 1713453518
transform 1 0 1256 0 1 170
box -9 -3 26 105
use INVX2  INVX2_294
timestamp 1713453518
transform 1 0 1216 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_295
timestamp 1713453518
transform 1 0 576 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_296
timestamp 1713453518
transform 1 0 368 0 1 170
box -9 -3 26 105
use INVX2  INVX2_297
timestamp 1713453518
transform 1 0 200 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_298
timestamp 1713453518
transform 1 0 216 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_299
timestamp 1713453518
transform 1 0 480 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_300
timestamp 1713453518
transform 1 0 2152 0 1 570
box -9 -3 26 105
use INVX2  INVX2_301
timestamp 1713453518
transform 1 0 1072 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_302
timestamp 1713453518
transform 1 0 1120 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_303
timestamp 1713453518
transform 1 0 872 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_304
timestamp 1713453518
transform 1 0 1808 0 1 370
box -9 -3 26 105
use INVX2  INVX2_305
timestamp 1713453518
transform 1 0 576 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_306
timestamp 1713453518
transform 1 0 1576 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_307
timestamp 1713453518
transform 1 0 1328 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_308
timestamp 1713453518
transform 1 0 1192 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_309
timestamp 1713453518
transform 1 0 1080 0 1 770
box -9 -3 26 105
use INVX2  INVX2_310
timestamp 1713453518
transform 1 0 1200 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_311
timestamp 1713453518
transform 1 0 1184 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_312
timestamp 1713453518
transform 1 0 1272 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_313
timestamp 1713453518
transform 1 0 3064 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_314
timestamp 1713453518
transform 1 0 3264 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_315
timestamp 1713453518
transform 1 0 3344 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_316
timestamp 1713453518
transform 1 0 3288 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_317
timestamp 1713453518
transform 1 0 3408 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_318
timestamp 1713453518
transform 1 0 2808 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_319
timestamp 1713453518
transform 1 0 3320 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_320
timestamp 1713453518
transform 1 0 2736 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_321
timestamp 1713453518
transform 1 0 560 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_322
timestamp 1713453518
transform 1 0 2480 0 1 570
box -9 -3 26 105
use INVX2  INVX2_323
timestamp 1713453518
transform 1 0 1320 0 1 970
box -9 -3 26 105
use INVX2  INVX2_324
timestamp 1713453518
transform 1 0 1976 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_325
timestamp 1713453518
transform 1 0 1888 0 1 770
box -9 -3 26 105
use INVX2  INVX2_326
timestamp 1713453518
transform 1 0 2672 0 1 570
box -9 -3 26 105
use INVX2  INVX2_327
timestamp 1713453518
transform 1 0 2464 0 1 570
box -9 -3 26 105
use INVX2  INVX2_328
timestamp 1713453518
transform 1 0 2808 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_329
timestamp 1713453518
transform 1 0 904 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_330
timestamp 1713453518
transform 1 0 840 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_331
timestamp 1713453518
transform 1 0 896 0 1 170
box -9 -3 26 105
use INVX2  INVX2_332
timestamp 1713453518
transform 1 0 232 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_333
timestamp 1713453518
transform 1 0 2576 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_334
timestamp 1713453518
transform 1 0 2944 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_335
timestamp 1713453518
transform 1 0 520 0 1 770
box -9 -3 26 105
use INVX2  INVX2_336
timestamp 1713453518
transform 1 0 2224 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_337
timestamp 1713453518
transform 1 0 216 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_338
timestamp 1713453518
transform 1 0 1040 0 1 570
box -9 -3 26 105
use INVX2  INVX2_339
timestamp 1713453518
transform 1 0 3056 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_340
timestamp 1713453518
transform 1 0 2160 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_341
timestamp 1713453518
transform 1 0 2456 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_342
timestamp 1713453518
transform 1 0 1792 0 1 370
box -9 -3 26 105
use INVX2  INVX2_343
timestamp 1713453518
transform 1 0 1448 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_344
timestamp 1713453518
transform 1 0 1520 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_345
timestamp 1713453518
transform 1 0 2664 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_346
timestamp 1713453518
transform 1 0 248 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_347
timestamp 1713453518
transform 1 0 144 0 1 570
box -9 -3 26 105
use INVX2  INVX2_348
timestamp 1713453518
transform 1 0 392 0 1 370
box -9 -3 26 105
use INVX2  INVX2_349
timestamp 1713453518
transform 1 0 1568 0 1 170
box -9 -3 26 105
use INVX2  INVX2_350
timestamp 1713453518
transform 1 0 1432 0 1 170
box -9 -3 26 105
use INVX2  INVX2_351
timestamp 1713453518
transform 1 0 1496 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_352
timestamp 1713453518
transform 1 0 1416 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1713453518
transform 1 0 2548 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1713453518
transform 1 0 2508 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1713453518
transform 1 0 2772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1713453518
transform 1 0 2612 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1713453518
transform 1 0 2868 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1713453518
transform 1 0 2828 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1713453518
transform 1 0 1204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1713453518
transform 1 0 1140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1713453518
transform 1 0 1132 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1713453518
transform 1 0 1132 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1713453518
transform 1 0 1092 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1713453518
transform 1 0 1084 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1713453518
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1713453518
transform 1 0 1292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1713453518
transform 1 0 1220 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1713453518
transform 1 0 1212 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1713453518
transform 1 0 1180 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1713453518
transform 1 0 1180 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1713453518
transform 1 0 1668 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1713453518
transform 1 0 1252 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1713453518
transform 1 0 1228 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1713453518
transform 1 0 1148 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1713453518
transform 1 0 1116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1713453518
transform 1 0 1100 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1713453518
transform 1 0 1676 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1713453518
transform 1 0 1244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1713453518
transform 1 0 1220 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1713453518
transform 1 0 1156 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1713453518
transform 1 0 1796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1713453518
transform 1 0 1244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1713453518
transform 1 0 1228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1713453518
transform 1 0 1140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1713453518
transform 1 0 1124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1713453518
transform 1 0 1884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1713453518
transform 1 0 1668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1713453518
transform 1 0 1588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1713453518
transform 1 0 1548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1713453518
transform 1 0 1484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1713453518
transform 1 0 1460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1713453518
transform 1 0 1772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1713453518
transform 1 0 1564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1713453518
transform 1 0 1532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1713453518
transform 1 0 1364 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1713453518
transform 1 0 3132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1713453518
transform 1 0 3132 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1713453518
transform 1 0 3132 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1713453518
transform 1 0 3420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1713453518
transform 1 0 3412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1713453518
transform 1 0 3396 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1713453518
transform 1 0 3348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1713453518
transform 1 0 3276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1713453518
transform 1 0 3444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1713453518
transform 1 0 3444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1713453518
transform 1 0 3420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1713453518
transform 1 0 3308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1713453518
transform 1 0 3356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1713453518
transform 1 0 3340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1713453518
transform 1 0 3252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1713453518
transform 1 0 3220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1713453518
transform 1 0 2324 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1713453518
transform 1 0 2300 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1713453518
transform 1 0 2276 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1713453518
transform 1 0 2172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1713453518
transform 1 0 2140 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1713453518
transform 1 0 2436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1713453518
transform 1 0 2380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1713453518
transform 1 0 2252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1713453518
transform 1 0 2236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1713453518
transform 1 0 396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1713453518
transform 1 0 316 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1713453518
transform 1 0 724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1713453518
transform 1 0 668 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1713453518
transform 1 0 172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1713453518
transform 1 0 100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1713453518
transform 1 0 188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1713453518
transform 1 0 84 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1713453518
transform 1 0 292 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1713453518
transform 1 0 212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1713453518
transform 1 0 172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1713453518
transform 1 0 124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1713453518
transform 1 0 252 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1713453518
transform 1 0 204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1713453518
transform 1 0 260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1713453518
transform 1 0 236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1713453518
transform 1 0 172 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1713453518
transform 1 0 140 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1713453518
transform 1 0 660 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1713453518
transform 1 0 548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1713453518
transform 1 0 388 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1713453518
transform 1 0 932 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1713453518
transform 1 0 772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1713453518
transform 1 0 444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1713453518
transform 1 0 612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1713453518
transform 1 0 604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1713453518
transform 1 0 404 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1713453518
transform 1 0 420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1713453518
transform 1 0 356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1713453518
transform 1 0 308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1713453518
transform 1 0 476 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1713453518
transform 1 0 180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1713453518
transform 1 0 140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1713453518
transform 1 0 428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1713453518
transform 1 0 252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1713453518
transform 1 0 220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1713453518
transform 1 0 1348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1713453518
transform 1 0 1244 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1713453518
transform 1 0 1236 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1713453518
transform 1 0 1308 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1713453518
transform 1 0 1268 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1713453518
transform 1 0 1236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1713453518
transform 1 0 1220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1713453518
transform 1 0 828 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1713453518
transform 1 0 828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1713453518
transform 1 0 988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1713453518
transform 1 0 900 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1713453518
transform 1 0 1028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1713453518
transform 1 0 876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1713453518
transform 1 0 996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1713453518
transform 1 0 828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1713453518
transform 1 0 932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1713453518
transform 1 0 796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1713453518
transform 1 0 988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1713453518
transform 1 0 756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1713453518
transform 1 0 980 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1713453518
transform 1 0 772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1713453518
transform 1 0 932 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1713453518
transform 1 0 796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1713453518
transform 1 0 1004 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1713453518
transform 1 0 772 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1713453518
transform 1 0 908 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1713453518
transform 1 0 804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1713453518
transform 1 0 1028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1713453518
transform 1 0 908 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1713453518
transform 1 0 948 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1713453518
transform 1 0 796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1713453518
transform 1 0 988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1713453518
transform 1 0 980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1713453518
transform 1 0 1044 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1713453518
transform 1 0 908 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1713453518
transform 1 0 1044 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1713453518
transform 1 0 940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1713453518
transform 1 0 1004 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1713453518
transform 1 0 900 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1713453518
transform 1 0 988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1713453518
transform 1 0 820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1713453518
transform 1 0 972 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1713453518
transform 1 0 844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1713453518
transform 1 0 948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1713453518
transform 1 0 812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1713453518
transform 1 0 1004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1713453518
transform 1 0 868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1713453518
transform 1 0 1028 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1713453518
transform 1 0 868 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1713453518
transform 1 0 980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1713453518
transform 1 0 836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1713453518
transform 1 0 996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1713453518
transform 1 0 860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1713453518
transform 1 0 1044 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1713453518
transform 1 0 892 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1713453518
transform 1 0 1028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1713453518
transform 1 0 1028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1713453518
transform 1 0 1076 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1713453518
transform 1 0 932 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1713453518
transform 1 0 1100 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1713453518
transform 1 0 1020 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1713453518
transform 1 0 1004 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1713453518
transform 1 0 964 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1713453518
transform 1 0 972 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1713453518
transform 1 0 876 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1713453518
transform 1 0 876 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1713453518
transform 1 0 852 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1713453518
transform 1 0 828 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1713453518
transform 1 0 804 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1713453518
transform 1 0 884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1713453518
transform 1 0 740 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1713453518
transform 1 0 772 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1713453518
transform 1 0 524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1713453518
transform 1 0 868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1713453518
transform 1 0 860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1713453518
transform 1 0 836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1713453518
transform 1 0 524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1713453518
transform 1 0 764 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1713453518
transform 1 0 708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1713453518
transform 1 0 756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1713453518
transform 1 0 196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1713453518
transform 1 0 724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1713453518
transform 1 0 356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1713453518
transform 1 0 700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1713453518
transform 1 0 284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1713453518
transform 1 0 764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1713453518
transform 1 0 316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1713453518
transform 1 0 740 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1713453518
transform 1 0 396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1713453518
transform 1 0 756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1713453518
transform 1 0 452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1713453518
transform 1 0 852 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1713453518
transform 1 0 396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1713453518
transform 1 0 740 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1713453518
transform 1 0 380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1713453518
transform 1 0 924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1713453518
transform 1 0 868 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1713453518
transform 1 0 868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1713453518
transform 1 0 820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1713453518
transform 1 0 844 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1713453518
transform 1 0 404 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1713453518
transform 1 0 756 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1713453518
transform 1 0 436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1713453518
transform 1 0 804 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1713453518
transform 1 0 436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1713453518
transform 1 0 748 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1713453518
transform 1 0 436 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1713453518
transform 1 0 812 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1713453518
transform 1 0 564 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1713453518
transform 1 0 796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1713453518
transform 1 0 388 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1713453518
transform 1 0 788 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1713453518
transform 1 0 420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1713453518
transform 1 0 812 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1713453518
transform 1 0 476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1713453518
transform 1 0 836 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1713453518
transform 1 0 484 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1713453518
transform 1 0 924 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1713453518
transform 1 0 436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1713453518
transform 1 0 900 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1713453518
transform 1 0 804 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1713453518
transform 1 0 972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1713453518
transform 1 0 780 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1713453518
transform 1 0 884 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1713453518
transform 1 0 468 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1713453518
transform 1 0 812 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1713453518
transform 1 0 500 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1713453518
transform 1 0 812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1713453518
transform 1 0 364 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1713453518
transform 1 0 708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1713453518
transform 1 0 444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1713453518
transform 1 0 700 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1713453518
transform 1 0 380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1713453518
transform 1 0 2508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1713453518
transform 1 0 2484 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1713453518
transform 1 0 2388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1713453518
transform 1 0 2340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1713453518
transform 1 0 1868 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1713453518
transform 1 0 1108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1713453518
transform 1 0 2620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1713453518
transform 1 0 2524 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1713453518
transform 1 0 2492 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1713453518
transform 1 0 2476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1713453518
transform 1 0 2436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1713453518
transform 1 0 2036 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1713453518
transform 1 0 1900 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1713453518
transform 1 0 1900 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1713453518
transform 1 0 1804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1713453518
transform 1 0 1380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1713453518
transform 1 0 2652 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1713453518
transform 1 0 2556 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1713453518
transform 1 0 1708 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1713453518
transform 1 0 1636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1713453518
transform 1 0 2988 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1713453518
transform 1 0 2924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1713453518
transform 1 0 2924 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1713453518
transform 1 0 2804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1713453518
transform 1 0 2796 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1713453518
transform 1 0 2772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1713453518
transform 1 0 1628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1713453518
transform 1 0 3068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1713453518
transform 1 0 3068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1713453518
transform 1 0 2932 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1713453518
transform 1 0 1748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1713453518
transform 1 0 2252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1713453518
transform 1 0 2252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1713453518
transform 1 0 1892 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1713453518
transform 1 0 1852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1713453518
transform 1 0 2420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1713453518
transform 1 0 2364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1713453518
transform 1 0 2092 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1713453518
transform 1 0 2052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1713453518
transform 1 0 1740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1713453518
transform 1 0 2356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1713453518
transform 1 0 2220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1713453518
transform 1 0 2572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1713453518
transform 1 0 2500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1713453518
transform 1 0 2396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1713453518
transform 1 0 3332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1713453518
transform 1 0 2900 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1713453518
transform 1 0 2324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1713453518
transform 1 0 2764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1713453518
transform 1 0 2644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1713453518
transform 1 0 2596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1713453518
transform 1 0 3196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1713453518
transform 1 0 2724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1713453518
transform 1 0 2452 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1713453518
transform 1 0 3316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1713453518
transform 1 0 3012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1713453518
transform 1 0 2964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1713453518
transform 1 0 3140 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1713453518
transform 1 0 3092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1713453518
transform 1 0 3036 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1713453518
transform 1 0 356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1713453518
transform 1 0 348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1713453518
transform 1 0 348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1713453518
transform 1 0 204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1713453518
transform 1 0 900 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1713453518
transform 1 0 828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1713453518
transform 1 0 828 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1713453518
transform 1 0 780 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1713453518
transform 1 0 764 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1713453518
transform 1 0 740 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1713453518
transform 1 0 724 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1713453518
transform 1 0 660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1713453518
transform 1 0 556 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1713453518
transform 1 0 988 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1713453518
transform 1 0 908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1713453518
transform 1 0 836 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1713453518
transform 1 0 764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1713453518
transform 1 0 748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1713453518
transform 1 0 892 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1713453518
transform 1 0 876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1713453518
transform 1 0 772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1713453518
transform 1 0 764 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1713453518
transform 1 0 668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1713453518
transform 1 0 644 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1713453518
transform 1 0 2996 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1713453518
transform 1 0 2972 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1713453518
transform 1 0 2964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1713453518
transform 1 0 2852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1713453518
transform 1 0 2804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1713453518
transform 1 0 2748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1713453518
transform 1 0 2700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1713453518
transform 1 0 2540 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1713453518
transform 1 0 2516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1713453518
transform 1 0 3044 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1713453518
transform 1 0 2164 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1713453518
transform 1 0 2052 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1713453518
transform 1 0 2044 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1713453518
transform 1 0 1956 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1713453518
transform 1 0 1892 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1713453518
transform 1 0 2460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1713453518
transform 1 0 2452 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1713453518
transform 1 0 2420 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1713453518
transform 1 0 2388 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1713453518
transform 1 0 2364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1713453518
transform 1 0 2348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1713453518
transform 1 0 1852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1713453518
transform 1 0 1804 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1713453518
transform 1 0 2364 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1713453518
transform 1 0 2284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1713453518
transform 1 0 2252 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1713453518
transform 1 0 2236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1713453518
transform 1 0 2196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1713453518
transform 1 0 2148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1713453518
transform 1 0 2412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1713453518
transform 1 0 2412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1713453518
transform 1 0 2356 0 1 585
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1713453518
transform 1 0 2356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1713453518
transform 1 0 2348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1713453518
transform 1 0 2292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1713453518
transform 1 0 1564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1713453518
transform 1 0 1564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1713453518
transform 1 0 1532 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1713453518
transform 1 0 1644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1713453518
transform 1 0 1628 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1713453518
transform 1 0 1620 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1713453518
transform 1 0 1596 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1713453518
transform 1 0 1588 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1713453518
transform 1 0 1524 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1713453518
transform 1 0 1500 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1713453518
transform 1 0 1476 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1713453518
transform 1 0 1340 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1713453518
transform 1 0 1284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1713453518
transform 1 0 1268 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1713453518
transform 1 0 1260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1713453518
transform 1 0 1244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1713453518
transform 1 0 1236 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1713453518
transform 1 0 1148 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1713453518
transform 1 0 1132 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1713453518
transform 1 0 1116 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1713453518
transform 1 0 1116 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1713453518
transform 1 0 1396 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1713453518
transform 1 0 1348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1713453518
transform 1 0 1348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1713453518
transform 1 0 1364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1713453518
transform 1 0 1316 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1713453518
transform 1 0 1260 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1713453518
transform 1 0 1260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1713453518
transform 1 0 1540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1713453518
transform 1 0 1508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1713453518
transform 1 0 1508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1713453518
transform 1 0 1500 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1713453518
transform 1 0 1484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1713453518
transform 1 0 1460 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1713453518
transform 1 0 1420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1713453518
transform 1 0 1404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1713453518
transform 1 0 1380 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1713453518
transform 1 0 1372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1713453518
transform 1 0 1292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1713453518
transform 1 0 1276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1713453518
transform 1 0 1268 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1713453518
transform 1 0 1252 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1713453518
transform 1 0 1244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1713453518
transform 1 0 1236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1713453518
transform 1 0 1236 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1713453518
transform 1 0 1188 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1713453518
transform 1 0 3332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1713453518
transform 1 0 3332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1713453518
transform 1 0 3276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1713453518
transform 1 0 3268 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1713453518
transform 1 0 3220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1713453518
transform 1 0 3412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1713453518
transform 1 0 3396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1713453518
transform 1 0 3364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1713453518
transform 1 0 3164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1713453518
transform 1 0 3100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1713453518
transform 1 0 2596 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1713453518
transform 1 0 3388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1713453518
transform 1 0 3372 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1713453518
transform 1 0 3348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1713453518
transform 1 0 3284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1713453518
transform 1 0 1276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1713453518
transform 1 0 1236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1713453518
transform 1 0 1228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1713453518
transform 1 0 1196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1713453518
transform 1 0 1100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1713453518
transform 1 0 1084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1713453518
transform 1 0 1084 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1713453518
transform 1 0 1068 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1713453518
transform 1 0 1028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1713453518
transform 1 0 1028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1713453518
transform 1 0 1020 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1713453518
transform 1 0 1012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1713453518
transform 1 0 1004 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1713453518
transform 1 0 1148 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1713453518
transform 1 0 1132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1713453518
transform 1 0 1124 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1713453518
transform 1 0 2564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1713453518
transform 1 0 2508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1713453518
transform 1 0 2500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1713453518
transform 1 0 2492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1713453518
transform 1 0 2484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1713453518
transform 1 0 2484 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1713453518
transform 1 0 2460 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1713453518
transform 1 0 2452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1713453518
transform 1 0 2156 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1713453518
transform 1 0 1340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1713453518
transform 1 0 1164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1713453518
transform 1 0 1100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1713453518
transform 1 0 1084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1713453518
transform 1 0 1068 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1713453518
transform 1 0 1068 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1713453518
transform 1 0 1028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1713453518
transform 1 0 1028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1713453518
transform 1 0 1204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1713453518
transform 1 0 1180 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1713453518
transform 1 0 1172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1713453518
transform 1 0 1124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1713453518
transform 1 0 1124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1713453518
transform 1 0 1300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1713453518
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1713453518
transform 1 0 1156 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1713453518
transform 1 0 1100 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1713453518
transform 1 0 1092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1713453518
transform 1 0 1196 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1713453518
transform 1 0 1196 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1713453518
transform 1 0 1188 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1713453518
transform 1 0 1180 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1713453518
transform 1 0 1156 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1713453518
transform 1 0 1148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1713453518
transform 1 0 1132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1713453518
transform 1 0 1132 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1713453518
transform 1 0 1116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1713453518
transform 1 0 1076 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1713453518
transform 1 0 1332 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1713453518
transform 1 0 1332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1713453518
transform 1 0 1308 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1713453518
transform 1 0 1292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1713453518
transform 1 0 1244 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1713453518
transform 1 0 1636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1713453518
transform 1 0 1636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1713453518
transform 1 0 1612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1713453518
transform 1 0 1604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1713453518
transform 1 0 1564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1713453518
transform 1 0 1532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1713453518
transform 1 0 1532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1713453518
transform 1 0 1580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1713453518
transform 1 0 1572 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1713453518
transform 1 0 1548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1713453518
transform 1 0 1540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1713453518
transform 1 0 1532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1713453518
transform 1 0 1508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1713453518
transform 1 0 1500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1713453518
transform 1 0 1492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1713453518
transform 1 0 1484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1713453518
transform 1 0 1388 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1713453518
transform 1 0 1356 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1713453518
transform 1 0 1300 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1713453518
transform 1 0 1236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1713453518
transform 1 0 1188 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1713453518
transform 1 0 1172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1713453518
transform 1 0 1164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1713453518
transform 1 0 1148 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1713453518
transform 1 0 1116 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1713453518
transform 1 0 1108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1713453518
transform 1 0 1436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1713453518
transform 1 0 1212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1713453518
transform 1 0 1188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1713453518
transform 1 0 1156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1713453518
transform 1 0 1596 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1713453518
transform 1 0 1596 0 1 1755
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1713453518
transform 1 0 1572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1713453518
transform 1 0 1524 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1713453518
transform 1 0 1492 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1713453518
transform 1 0 1532 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1713453518
transform 1 0 1516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1713453518
transform 1 0 1484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1713453518
transform 1 0 1436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1713453518
transform 1 0 1340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1713453518
transform 1 0 1300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1713453518
transform 1 0 1300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1713453518
transform 1 0 1292 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1713453518
transform 1 0 1220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1713453518
transform 1 0 1404 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1713453518
transform 1 0 1380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1713453518
transform 1 0 1212 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1713453518
transform 1 0 1204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1713453518
transform 1 0 1196 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1713453518
transform 1 0 1148 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1713453518
transform 1 0 1148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1713453518
transform 1 0 1100 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1713453518
transform 1 0 1620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1713453518
transform 1 0 1524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1713453518
transform 1 0 1228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1713453518
transform 1 0 1140 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1713453518
transform 1 0 1140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1713453518
transform 1 0 1548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1713453518
transform 1 0 1548 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1713453518
transform 1 0 1524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1713453518
transform 1 0 1492 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1713453518
transform 1 0 1484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1713453518
transform 1 0 1644 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1713453518
transform 1 0 1636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1713453518
transform 1 0 1636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1713453518
transform 1 0 1628 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1713453518
transform 1 0 1612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1713453518
transform 1 0 1444 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1713453518
transform 1 0 1260 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1713453518
transform 1 0 1260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1713453518
transform 1 0 1236 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1713453518
transform 1 0 1212 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1713453518
transform 1 0 1204 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1713453518
transform 1 0 1172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1713453518
transform 1 0 1404 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1713453518
transform 1 0 1380 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1713453518
transform 1 0 1364 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1713453518
transform 1 0 1324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1713453518
transform 1 0 1260 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1713453518
transform 1 0 1228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1713453518
transform 1 0 1132 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1713453518
transform 1 0 1132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1713453518
transform 1 0 1108 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1713453518
transform 1 0 1436 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1713453518
transform 1 0 1388 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1713453518
transform 1 0 1388 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1713453518
transform 1 0 1332 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1713453518
transform 1 0 1276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1713453518
transform 1 0 1180 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1713453518
transform 1 0 1692 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1713453518
transform 1 0 1636 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1713453518
transform 1 0 1340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1713453518
transform 1 0 1324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1713453518
transform 1 0 1276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1713453518
transform 1 0 1212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1713453518
transform 1 0 1644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1713453518
transform 1 0 1596 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1713453518
transform 1 0 1468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1713453518
transform 1 0 1420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1713453518
transform 1 0 1412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1713453518
transform 1 0 1412 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1713453518
transform 1 0 1404 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1713453518
transform 1 0 1388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1713453518
transform 1 0 1244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1713453518
transform 1 0 1236 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1713453518
transform 1 0 1196 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1713453518
transform 1 0 1188 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1713453518
transform 1 0 1724 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1713453518
transform 1 0 1684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1713453518
transform 1 0 1420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1713453518
transform 1 0 1388 0 1 2055
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1713453518
transform 1 0 1388 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1713453518
transform 1 0 1348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1713453518
transform 1 0 1348 0 1 2055
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1713453518
transform 1 0 1348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1713453518
transform 1 0 1316 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1713453518
transform 1 0 1164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1713453518
transform 1 0 1156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1713453518
transform 1 0 1124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1713453518
transform 1 0 1116 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1713453518
transform 1 0 1380 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1713453518
transform 1 0 1284 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1713453518
transform 1 0 1172 0 1 2895
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1713453518
transform 1 0 1164 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1713453518
transform 1 0 1164 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1713453518
transform 1 0 1164 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1713453518
transform 1 0 1684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1713453518
transform 1 0 1628 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1713453518
transform 1 0 1628 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1713453518
transform 1 0 1572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1713453518
transform 1 0 1556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1713453518
transform 1 0 1460 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1713453518
transform 1 0 1636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1713453518
transform 1 0 1612 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1713453518
transform 1 0 1572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1713453518
transform 1 0 1524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1713453518
transform 1 0 1508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1713453518
transform 1 0 1436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1713453518
transform 1 0 1108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1713453518
transform 1 0 1092 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1713453518
transform 1 0 1060 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1713453518
transform 1 0 1028 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1713453518
transform 1 0 1028 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1713453518
transform 1 0 1228 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1713453518
transform 1 0 1212 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1713453518
transform 1 0 1212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1713453518
transform 1 0 1444 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1713453518
transform 1 0 1388 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1713453518
transform 1 0 1380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1713453518
transform 1 0 1372 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1713453518
transform 1 0 1356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1713453518
transform 1 0 1180 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1713453518
transform 1 0 1164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1713453518
transform 1 0 1156 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1713453518
transform 1 0 1148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1713453518
transform 1 0 1380 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1713453518
transform 1 0 1364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1713453518
transform 1 0 1204 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1713453518
transform 1 0 1172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1713453518
transform 1 0 1628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1713453518
transform 1 0 1492 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1713453518
transform 1 0 1492 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1713453518
transform 1 0 1492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1713453518
transform 1 0 1476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1713453518
transform 1 0 1452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1713453518
transform 1 0 1532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1713453518
transform 1 0 1484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1713453518
transform 1 0 1476 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1713453518
transform 1 0 1444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1713453518
transform 1 0 1396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1713453518
transform 1 0 1340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1713453518
transform 1 0 1324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1713453518
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1713453518
transform 1 0 1692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1713453518
transform 1 0 1668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1713453518
transform 1 0 1324 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1713453518
transform 1 0 1292 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1713453518
transform 1 0 1284 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1713453518
transform 1 0 1180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1713453518
transform 1 0 1140 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1713453518
transform 1 0 1100 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1713453518
transform 1 0 1444 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1713453518
transform 1 0 1420 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1713453518
transform 1 0 1404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1713453518
transform 1 0 1380 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1713453518
transform 1 0 1380 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1713453518
transform 1 0 1708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1713453518
transform 1 0 1684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1713453518
transform 1 0 1652 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1713453518
transform 1 0 1580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1713453518
transform 1 0 1500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1713453518
transform 1 0 1492 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1713453518
transform 1 0 1684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1713453518
transform 1 0 1628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1713453518
transform 1 0 1612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1713453518
transform 1 0 1524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1713453518
transform 1 0 1492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1713453518
transform 1 0 1460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1713453518
transform 1 0 1460 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1713453518
transform 1 0 1428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1713453518
transform 1 0 1396 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1713453518
transform 1 0 1388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1713453518
transform 1 0 1620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1713453518
transform 1 0 1620 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1713453518
transform 1 0 1492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1713453518
transform 1 0 1244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1713453518
transform 1 0 1204 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1713453518
transform 1 0 1676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1713453518
transform 1 0 1604 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1713453518
transform 1 0 1492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1713453518
transform 1 0 1324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1713453518
transform 1 0 1284 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1713453518
transform 1 0 1268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1713453518
transform 1 0 1252 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1713453518
transform 1 0 1252 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1713453518
transform 1 0 1212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1713453518
transform 1 0 1132 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1713453518
transform 1 0 1612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1713453518
transform 1 0 1532 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1713453518
transform 1 0 1452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1713453518
transform 1 0 1436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1713453518
transform 1 0 1540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1713453518
transform 1 0 1404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1713453518
transform 1 0 1372 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1713453518
transform 1 0 1340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1713453518
transform 1 0 1476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1713453518
transform 1 0 1476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1713453518
transform 1 0 2460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1713453518
transform 1 0 1692 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1713453518
transform 1 0 3092 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1713453518
transform 1 0 3084 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1713453518
transform 1 0 2996 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1713453518
transform 1 0 3124 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1713453518
transform 1 0 3060 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1713453518
transform 1 0 3060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1713453518
transform 1 0 3020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1713453518
transform 1 0 2908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1713453518
transform 1 0 3316 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1713453518
transform 1 0 3316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1713453518
transform 1 0 3308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1713453518
transform 1 0 3284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1713453518
transform 1 0 3276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1713453518
transform 1 0 3420 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1713453518
transform 1 0 3388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1713453518
transform 1 0 3308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1713453518
transform 1 0 3268 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1713453518
transform 1 0 3268 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1713453518
transform 1 0 2788 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1713453518
transform 1 0 3388 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1713453518
transform 1 0 3332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1713453518
transform 1 0 3268 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1713453518
transform 1 0 3196 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1713453518
transform 1 0 3076 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1713453518
transform 1 0 3388 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1713453518
transform 1 0 3388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1713453518
transform 1 0 3020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1713453518
transform 1 0 2820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1713453518
transform 1 0 2244 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1713453518
transform 1 0 2148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1713453518
transform 1 0 3412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1713453518
transform 1 0 2812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1713453518
transform 1 0 2740 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1713453518
transform 1 0 2716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1713453518
transform 1 0 2708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1713453518
transform 1 0 2708 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1713453518
transform 1 0 2692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1713453518
transform 1 0 2148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1713453518
transform 1 0 2900 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1713453518
transform 1 0 2796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1713453518
transform 1 0 2772 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1713453518
transform 1 0 2628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1713453518
transform 1 0 2124 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1713453518
transform 1 0 1900 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1713453518
transform 1 0 1796 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1713453518
transform 1 0 3428 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1713453518
transform 1 0 3428 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1713453518
transform 1 0 3292 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1713453518
transform 1 0 3260 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1713453518
transform 1 0 3244 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1713453518
transform 1 0 3220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1713453518
transform 1 0 3076 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1713453518
transform 1 0 3052 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1713453518
transform 1 0 2988 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1713453518
transform 1 0 2444 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1713453518
transform 1 0 1852 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1713453518
transform 1 0 1724 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1713453518
transform 1 0 3340 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1713453518
transform 1 0 3340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1713453518
transform 1 0 3316 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1713453518
transform 1 0 3100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1713453518
transform 1 0 2924 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1713453518
transform 1 0 2916 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1713453518
transform 1 0 3372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1713453518
transform 1 0 3348 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1713453518
transform 1 0 3348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1713453518
transform 1 0 3340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1713453518
transform 1 0 3044 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1713453518
transform 1 0 2980 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1713453518
transform 1 0 2980 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1713453518
transform 1 0 2756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1713453518
transform 1 0 2684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1713453518
transform 1 0 1980 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1713453518
transform 1 0 1964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1713453518
transform 1 0 1948 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1713453518
transform 1 0 3268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1713453518
transform 1 0 3260 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1713453518
transform 1 0 3228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1713453518
transform 1 0 3156 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1713453518
transform 1 0 3124 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1713453518
transform 1 0 3116 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1713453518
transform 1 0 2628 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1713453518
transform 1 0 2596 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1713453518
transform 1 0 2372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1713453518
transform 1 0 2092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1713453518
transform 1 0 1428 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1713453518
transform 1 0 2956 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1713453518
transform 1 0 2924 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1713453518
transform 1 0 2852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1713453518
transform 1 0 2548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1713453518
transform 1 0 1924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1713453518
transform 1 0 1836 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1713453518
transform 1 0 3180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1713453518
transform 1 0 3132 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1713453518
transform 1 0 3124 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1713453518
transform 1 0 3116 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1713453518
transform 1 0 3116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1713453518
transform 1 0 3020 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1713453518
transform 1 0 2964 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1713453518
transform 1 0 2964 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1713453518
transform 1 0 2860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1713453518
transform 1 0 2812 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1713453518
transform 1 0 3308 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1713453518
transform 1 0 3036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1713453518
transform 1 0 3028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1713453518
transform 1 0 2980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1713453518
transform 1 0 2876 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1713453518
transform 1 0 2300 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1713453518
transform 1 0 3396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1713453518
transform 1 0 3388 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1713453518
transform 1 0 3340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1713453518
transform 1 0 3300 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1713453518
transform 1 0 3292 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1713453518
transform 1 0 3372 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1713453518
transform 1 0 3340 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1713453518
transform 1 0 3292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1713453518
transform 1 0 3196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1713453518
transform 1 0 3308 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1713453518
transform 1 0 3308 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1713453518
transform 1 0 1804 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1713453518
transform 1 0 1804 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1713453518
transform 1 0 3372 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1713453518
transform 1 0 2972 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1713453518
transform 1 0 1916 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1713453518
transform 1 0 1828 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1713453518
transform 1 0 1764 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1713453518
transform 1 0 2884 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1713453518
transform 1 0 2788 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1713453518
transform 1 0 2788 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1713453518
transform 1 0 1980 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1713453518
transform 1 0 1508 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1713453518
transform 1 0 1460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1713453518
transform 1 0 1428 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1713453518
transform 1 0 3284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1713453518
transform 1 0 3284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1713453518
transform 1 0 3260 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1713453518
transform 1 0 3260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1713453518
transform 1 0 3236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1713453518
transform 1 0 3236 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1713453518
transform 1 0 3228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1713453518
transform 1 0 2748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1713453518
transform 1 0 2748 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1713453518
transform 1 0 2740 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1713453518
transform 1 0 2740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1713453518
transform 1 0 2364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1713453518
transform 1 0 1948 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1713453518
transform 1 0 2916 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1713453518
transform 1 0 2836 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1713453518
transform 1 0 2764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1713453518
transform 1 0 2620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1713453518
transform 1 0 2548 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1713453518
transform 1 0 3356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1713453518
transform 1 0 3340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1713453518
transform 1 0 3332 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1713453518
transform 1 0 3308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1713453518
transform 1 0 2796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1713453518
transform 1 0 2652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1713453518
transform 1 0 2212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1713453518
transform 1 0 2252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1713453518
transform 1 0 2036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1713453518
transform 1 0 1900 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1713453518
transform 1 0 2212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1713453518
transform 1 0 2084 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1713453518
transform 1 0 1748 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1713453518
transform 1 0 2884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1713453518
transform 1 0 2836 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1713453518
transform 1 0 2580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1713453518
transform 1 0 2580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1713453518
transform 1 0 1908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1713453518
transform 1 0 1908 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1713453518
transform 1 0 3404 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1713453518
transform 1 0 3380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1713453518
transform 1 0 3348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1713453518
transform 1 0 3212 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1713453518
transform 1 0 3212 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1713453518
transform 1 0 3164 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1713453518
transform 1 0 3148 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1713453518
transform 1 0 3044 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1713453518
transform 1 0 3036 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1713453518
transform 1 0 1812 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1713453518
transform 1 0 1684 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1713453518
transform 1 0 3300 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1713453518
transform 1 0 3300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1713453518
transform 1 0 3340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1713453518
transform 1 0 3332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1713453518
transform 1 0 3324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1713453518
transform 1 0 3324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1713453518
transform 1 0 3052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1713453518
transform 1 0 2820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1713453518
transform 1 0 2668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1713453518
transform 1 0 2140 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1713453518
transform 1 0 3180 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1713453518
transform 1 0 3036 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1713453518
transform 1 0 2692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1713453518
transform 1 0 2220 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1713453518
transform 1 0 3396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1713453518
transform 1 0 3348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1713453518
transform 1 0 3276 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1713453518
transform 1 0 3236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1713453518
transform 1 0 2412 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1713453518
transform 1 0 2340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1713453518
transform 1 0 3124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1713453518
transform 1 0 3124 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1713453518
transform 1 0 3108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1713453518
transform 1 0 2716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1713453518
transform 1 0 2508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1713453518
transform 1 0 2252 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1713453518
transform 1 0 1972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1713453518
transform 1 0 1948 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1713453518
transform 1 0 3244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1713453518
transform 1 0 3212 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1713453518
transform 1 0 3148 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1713453518
transform 1 0 3108 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1713453518
transform 1 0 3084 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1713453518
transform 1 0 2868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1713453518
transform 1 0 2868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1713453518
transform 1 0 2812 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1713453518
transform 1 0 2156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1713453518
transform 1 0 1980 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1713453518
transform 1 0 1900 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1713453518
transform 1 0 3028 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1713453518
transform 1 0 2932 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1713453518
transform 1 0 2916 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1713453518
transform 1 0 3148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1713453518
transform 1 0 2964 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1713453518
transform 1 0 2604 0 1 2095
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1713453518
transform 1 0 2380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1713453518
transform 1 0 1948 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1713453518
transform 1 0 2828 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1713453518
transform 1 0 2812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1713453518
transform 1 0 2628 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1713453518
transform 1 0 2428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1713453518
transform 1 0 1996 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1713453518
transform 1 0 3140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1713453518
transform 1 0 2964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1713453518
transform 1 0 2908 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1713453518
transform 1 0 2732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1713453518
transform 1 0 2716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1713453518
transform 1 0 2708 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1713453518
transform 1 0 2700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1713453518
transform 1 0 2300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1713453518
transform 1 0 3012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1713453518
transform 1 0 2940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1713453518
transform 1 0 2932 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1713453518
transform 1 0 2996 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1713453518
transform 1 0 2932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1713453518
transform 1 0 2900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1713453518
transform 1 0 2828 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1713453518
transform 1 0 2780 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1713453518
transform 1 0 2196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1713453518
transform 1 0 2188 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1713453518
transform 1 0 2236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1713453518
transform 1 0 2004 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1713453518
transform 1 0 1828 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1713453518
transform 1 0 3028 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1713453518
transform 1 0 3004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1713453518
transform 1 0 2988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1713453518
transform 1 0 2932 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1713453518
transform 1 0 2844 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1713453518
transform 1 0 2020 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1713453518
transform 1 0 3444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1713453518
transform 1 0 3404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1713453518
transform 1 0 3308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1713453518
transform 1 0 3156 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1713453518
transform 1 0 3108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1713453518
transform 1 0 2484 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1713453518
transform 1 0 2444 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1713453518
transform 1 0 2380 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1713453518
transform 1 0 2204 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1713453518
transform 1 0 2196 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1713453518
transform 1 0 3276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1713453518
transform 1 0 3260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1713453518
transform 1 0 3260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1713453518
transform 1 0 3244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1713453518
transform 1 0 3324 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1713453518
transform 1 0 3292 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1713453518
transform 1 0 3044 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1713453518
transform 1 0 2668 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1713453518
transform 1 0 2460 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1713453518
transform 1 0 2876 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1713453518
transform 1 0 2868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1713453518
transform 1 0 2860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1713453518
transform 1 0 2628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1713453518
transform 1 0 2620 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1713453518
transform 1 0 2804 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1713453518
transform 1 0 2788 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1713453518
transform 1 0 2724 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1713453518
transform 1 0 2196 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1713453518
transform 1 0 2500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1713453518
transform 1 0 2244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1713453518
transform 1 0 2004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1713453518
transform 1 0 3052 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1713453518
transform 1 0 2996 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1713453518
transform 1 0 2820 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1713453518
transform 1 0 2644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1713453518
transform 1 0 2564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1713453518
transform 1 0 1900 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1713453518
transform 1 0 1868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1713453518
transform 1 0 244 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1713453518
transform 1 0 220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1713453518
transform 1 0 220 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1713453518
transform 1 0 204 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1713453518
transform 1 0 236 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1713453518
transform 1 0 212 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1713453518
transform 1 0 284 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1713453518
transform 1 0 260 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1713453518
transform 1 0 468 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1713453518
transform 1 0 452 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1713453518
transform 1 0 660 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1713453518
transform 1 0 636 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1713453518
transform 1 0 644 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1713453518
transform 1 0 604 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1713453518
transform 1 0 260 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1713453518
transform 1 0 236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1713453518
transform 1 0 300 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1713453518
transform 1 0 276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1713453518
transform 1 0 300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1713453518
transform 1 0 284 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1713453518
transform 1 0 252 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1713453518
transform 1 0 212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1713453518
transform 1 0 196 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1713453518
transform 1 0 188 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1713453518
transform 1 0 428 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1713453518
transform 1 0 388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1713453518
transform 1 0 260 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1713453518
transform 1 0 220 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1713453518
transform 1 0 260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1713453518
transform 1 0 244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1713453518
transform 1 0 268 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1713453518
transform 1 0 244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1713453518
transform 1 0 260 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1713453518
transform 1 0 220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1713453518
transform 1 0 220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1713453518
transform 1 0 148 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1713453518
transform 1 0 324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1713453518
transform 1 0 284 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1713453518
transform 1 0 476 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1713453518
transform 1 0 356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1713453518
transform 1 0 180 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1713453518
transform 1 0 156 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1713453518
transform 1 0 236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1713453518
transform 1 0 220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1713453518
transform 1 0 268 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1713453518
transform 1 0 244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1713453518
transform 1 0 236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1713453518
transform 1 0 220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1713453518
transform 1 0 260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1713453518
transform 1 0 228 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1713453518
transform 1 0 196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1713453518
transform 1 0 92 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1713453518
transform 1 0 92 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1713453518
transform 1 0 220 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1713453518
transform 1 0 116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1713453518
transform 1 0 148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1713453518
transform 1 0 116 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1713453518
transform 1 0 436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1713453518
transform 1 0 436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1713453518
transform 1 0 380 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1713453518
transform 1 0 308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1713453518
transform 1 0 324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1713453518
transform 1 0 292 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1713453518
transform 1 0 988 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1713453518
transform 1 0 964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1713453518
transform 1 0 932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1713453518
transform 1 0 860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1713453518
transform 1 0 812 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1713453518
transform 1 0 676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1713453518
transform 1 0 588 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1713453518
transform 1 0 468 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1713453518
transform 1 0 1372 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1713453518
transform 1 0 1292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1713453518
transform 1 0 996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1713453518
transform 1 0 884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1713453518
transform 1 0 820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1713453518
transform 1 0 740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1713453518
transform 1 0 740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1713453518
transform 1 0 700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1713453518
transform 1 0 636 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1713453518
transform 1 0 580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1713453518
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1713453518
transform 1 0 852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1713453518
transform 1 0 820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1713453518
transform 1 0 812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1713453518
transform 1 0 2396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1713453518
transform 1 0 1308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1713453518
transform 1 0 1044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1713453518
transform 1 0 1036 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1713453518
transform 1 0 980 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1713453518
transform 1 0 924 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1713453518
transform 1 0 892 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1713453518
transform 1 0 692 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1713453518
transform 1 0 692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1713453518
transform 1 0 572 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1713453518
transform 1 0 548 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1713453518
transform 1 0 2428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1713453518
transform 1 0 2364 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1713453518
transform 1 0 2364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1713453518
transform 1 0 2260 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1713453518
transform 1 0 2260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1713453518
transform 1 0 2212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1713453518
transform 1 0 2076 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1713453518
transform 1 0 2132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1713453518
transform 1 0 2012 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1713453518
transform 1 0 2004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1713453518
transform 1 0 3100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1713453518
transform 1 0 2940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1713453518
transform 1 0 2972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1713453518
transform 1 0 2956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1713453518
transform 1 0 2908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1713453518
transform 1 0 2860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1713453518
transform 1 0 2748 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1713453518
transform 1 0 2636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1713453518
transform 1 0 2436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1713453518
transform 1 0 2012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1713453518
transform 1 0 1948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1713453518
transform 1 0 2276 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1713453518
transform 1 0 1676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1713453518
transform 1 0 1652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1713453518
transform 1 0 1540 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1713453518
transform 1 0 1356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1713453518
transform 1 0 1460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1713453518
transform 1 0 1396 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1713453518
transform 1 0 3108 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1713453518
transform 1 0 3052 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1713453518
transform 1 0 2868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1713453518
transform 1 0 2412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1713453518
transform 1 0 1956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1713453518
transform 1 0 412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1713453518
transform 1 0 380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1713453518
transform 1 0 3324 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1713453518
transform 1 0 2692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1713453518
transform 1 0 3148 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1713453518
transform 1 0 2652 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1713453518
transform 1 0 2652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1713453518
transform 1 0 2748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1713453518
transform 1 0 2508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1713453518
transform 1 0 3164 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1713453518
transform 1 0 3124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1713453518
transform 1 0 2700 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1713453518
transform 1 0 2620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1713453518
transform 1 0 2500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1713453518
transform 1 0 3012 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1713453518
transform 1 0 2964 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1713453518
transform 1 0 2116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1713453518
transform 1 0 2076 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1713453518
transform 1 0 2588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1713453518
transform 1 0 2588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1713453518
transform 1 0 2132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1713453518
transform 1 0 2124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1713453518
transform 1 0 1916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1713453518
transform 1 0 1916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1713453518
transform 1 0 2596 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1713453518
transform 1 0 2556 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1713453518
transform 1 0 2100 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1713453518
transform 1 0 2100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1713453518
transform 1 0 1348 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1713453518
transform 1 0 1348 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1713453518
transform 1 0 1324 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1713453518
transform 1 0 1300 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1713453518
transform 1 0 1700 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1713453518
transform 1 0 1684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1713453518
transform 1 0 1628 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1713453518
transform 1 0 1620 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1713453518
transform 1 0 2076 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1713453518
transform 1 0 1908 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1713453518
transform 1 0 1764 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1713453518
transform 1 0 1452 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1713453518
transform 1 0 1396 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1713453518
transform 1 0 1372 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1713453518
transform 1 0 1740 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1713453518
transform 1 0 1604 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1713453518
transform 1 0 1572 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1713453518
transform 1 0 1516 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1713453518
transform 1 0 2260 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1713453518
transform 1 0 1868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1713453518
transform 1 0 2020 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1713453518
transform 1 0 1900 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1713453518
transform 1 0 1724 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1713453518
transform 1 0 1404 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1713453518
transform 1 0 1404 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1713453518
transform 1 0 2220 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1713453518
transform 1 0 2204 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1713453518
transform 1 0 2172 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1713453518
transform 1 0 2172 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1713453518
transform 1 0 2260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1713453518
transform 1 0 2260 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1713453518
transform 1 0 2100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1713453518
transform 1 0 3044 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1713453518
transform 1 0 3004 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1713453518
transform 1 0 1364 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1713453518
transform 1 0 1196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1713453518
transform 1 0 3012 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1713453518
transform 1 0 3012 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1713453518
transform 1 0 2436 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1713453518
transform 1 0 1244 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1713453518
transform 1 0 3060 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1713453518
transform 1 0 2908 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1713453518
transform 1 0 2900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1713453518
transform 1 0 2868 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1713453518
transform 1 0 2868 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1713453518
transform 1 0 3284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1713453518
transform 1 0 3276 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1713453518
transform 1 0 2276 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1713453518
transform 1 0 1308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1713453518
transform 1 0 2668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1713453518
transform 1 0 2668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1713453518
transform 1 0 3412 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1713453518
transform 1 0 3388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1713453518
transform 1 0 548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1713453518
transform 1 0 508 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1713453518
transform 1 0 3396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1713453518
transform 1 0 3380 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1713453518
transform 1 0 2244 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1713453518
transform 1 0 2244 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1713453518
transform 1 0 2772 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1713453518
transform 1 0 2684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1713453518
transform 1 0 2612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1713453518
transform 1 0 3076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1713453518
transform 1 0 3052 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1713453518
transform 1 0 3412 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1713453518
transform 1 0 3388 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1713453518
transform 1 0 3092 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1713453518
transform 1 0 3092 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1713453518
transform 1 0 2388 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1713453518
transform 1 0 2340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1713453518
transform 1 0 524 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1713453518
transform 1 0 460 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1713453518
transform 1 0 420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1713453518
transform 1 0 580 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1713453518
transform 1 0 580 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1713453518
transform 1 0 572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1713453518
transform 1 0 764 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1713453518
transform 1 0 764 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1713453518
transform 1 0 724 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1713453518
transform 1 0 676 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1713453518
transform 1 0 644 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1713453518
transform 1 0 2340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1713453518
transform 1 0 2340 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1713453518
transform 1 0 2788 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1713453518
transform 1 0 2644 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1713453518
transform 1 0 2596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1713453518
transform 1 0 3412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1713453518
transform 1 0 3364 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1713453518
transform 1 0 1892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1713453518
transform 1 0 1892 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1713453518
transform 1 0 2836 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1713453518
transform 1 0 2772 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1713453518
transform 1 0 2380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1713453518
transform 1 0 2156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1713453518
transform 1 0 3036 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1713453518
transform 1 0 2996 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1713453518
transform 1 0 2956 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1713453518
transform 1 0 2716 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1713453518
transform 1 0 2660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1713453518
transform 1 0 3012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1713453518
transform 1 0 2900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1713453518
transform 1 0 636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1713453518
transform 1 0 636 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1713453518
transform 1 0 548 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1713453518
transform 1 0 548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1713453518
transform 1 0 524 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1713453518
transform 1 0 508 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1713453518
transform 1 0 508 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1713453518
transform 1 0 700 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1713453518
transform 1 0 700 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1713453518
transform 1 0 636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1713453518
transform 1 0 636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1713453518
transform 1 0 604 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1713453518
transform 1 0 580 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1713453518
transform 1 0 2188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1713453518
transform 1 0 2060 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1713453518
transform 1 0 2996 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1713453518
transform 1 0 2956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1713453518
transform 1 0 3404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1713453518
transform 1 0 3404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1713453518
transform 1 0 3412 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1713453518
transform 1 0 3380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1713453518
transform 1 0 2524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1713453518
transform 1 0 2492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1713453518
transform 1 0 3132 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1713453518
transform 1 0 2780 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1713453518
transform 1 0 2756 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1713453518
transform 1 0 2556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1713453518
transform 1 0 2556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1713453518
transform 1 0 3076 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1713453518
transform 1 0 2932 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1713453518
transform 1 0 2804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1713453518
transform 1 0 2660 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1713453518
transform 1 0 2724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1713453518
transform 1 0 2660 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1713453518
transform 1 0 2660 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1713453518
transform 1 0 2636 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1713453518
transform 1 0 2620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1713453518
transform 1 0 3164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1713453518
transform 1 0 3052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1713453518
transform 1 0 532 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1713453518
transform 1 0 500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1713453518
transform 1 0 500 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1713453518
transform 1 0 644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1713453518
transform 1 0 596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1713453518
transform 1 0 556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1713453518
transform 1 0 556 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1713453518
transform 1 0 3292 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1713453518
transform 1 0 2724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1713453518
transform 1 0 2628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1713453518
transform 1 0 2428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1713453518
transform 1 0 2412 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1713453518
transform 1 0 732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1713453518
transform 1 0 700 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1713453518
transform 1 0 692 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1713453518
transform 1 0 676 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1713453518
transform 1 0 676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1713453518
transform 1 0 612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1713453518
transform 1 0 604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1713453518
transform 1 0 548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1713453518
transform 1 0 492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1713453518
transform 1 0 692 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1713453518
transform 1 0 652 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1713453518
transform 1 0 484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1713453518
transform 1 0 476 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1713453518
transform 1 0 468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1713453518
transform 1 0 580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1713453518
transform 1 0 532 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1713453518
transform 1 0 460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1713453518
transform 1 0 452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1713453518
transform 1 0 564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1713453518
transform 1 0 548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1713453518
transform 1 0 484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1713453518
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1713453518
transform 1 0 388 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1713453518
transform 1 0 364 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1713453518
transform 1 0 1828 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1713453518
transform 1 0 1804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1713453518
transform 1 0 1772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1713453518
transform 1 0 2132 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1713453518
transform 1 0 1988 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1713453518
transform 1 0 1956 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1713453518
transform 1 0 1940 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1713453518
transform 1 0 1916 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1713453518
transform 1 0 1860 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1713453518
transform 1 0 1788 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1713453518
transform 1 0 1756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1713453518
transform 1 0 2052 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1713453518
transform 1 0 2012 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1713453518
transform 1 0 1916 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1713453518
transform 1 0 1884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1713453518
transform 1 0 1860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1713453518
transform 1 0 2148 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1713453518
transform 1 0 2068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1713453518
transform 1 0 2052 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1713453518
transform 1 0 2348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1713453518
transform 1 0 2220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1713453518
transform 1 0 2220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1713453518
transform 1 0 1300 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1713453518
transform 1 0 1276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1713453518
transform 1 0 1228 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1713453518
transform 1 0 1012 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1713453518
transform 1 0 596 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1713453518
transform 1 0 588 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1713453518
transform 1 0 588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1713453518
transform 1 0 556 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1713453518
transform 1 0 548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1713453518
transform 1 0 540 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1713453518
transform 1 0 1068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1713453518
transform 1 0 1068 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1713453518
transform 1 0 900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1713453518
transform 1 0 876 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1713453518
transform 1 0 716 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1713453518
transform 1 0 668 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1713453518
transform 1 0 556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1713453518
transform 1 0 540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1713453518
transform 1 0 436 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1713453518
transform 1 0 412 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1713453518
transform 1 0 396 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1713453518
transform 1 0 348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1713453518
transform 1 0 316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1713453518
transform 1 0 188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1713453518
transform 1 0 148 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1713453518
transform 1 0 220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1713453518
transform 1 0 188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1713453518
transform 1 0 532 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1713453518
transform 1 0 484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1713453518
transform 1 0 468 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1713453518
transform 1 0 452 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1713453518
transform 1 0 396 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1713453518
transform 1 0 268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1713453518
transform 1 0 140 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1713453518
transform 1 0 100 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1713453518
transform 1 0 964 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1713453518
transform 1 0 956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1713453518
transform 1 0 852 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1713453518
transform 1 0 636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1713453518
transform 1 0 524 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1713453518
transform 1 0 468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1713453518
transform 1 0 404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1713453518
transform 1 0 316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1713453518
transform 1 0 316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1713453518
transform 1 0 212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1713453518
transform 1 0 164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1713453518
transform 1 0 108 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1713453518
transform 1 0 100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1713453518
transform 1 0 92 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1713453518
transform 1 0 340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1713453518
transform 1 0 268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1713453518
transform 1 0 220 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1713453518
transform 1 0 204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1713453518
transform 1 0 100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1713453518
transform 1 0 100 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1713453518
transform 1 0 100 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1713453518
transform 1 0 100 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1713453518
transform 1 0 92 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1713453518
transform 1 0 92 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1713453518
transform 1 0 92 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1713453518
transform 1 0 92 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1713453518
transform 1 0 92 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1713453518
transform 1 0 92 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1713453518
transform 1 0 1076 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1713453518
transform 1 0 1060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1713453518
transform 1 0 524 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1713453518
transform 1 0 516 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1713453518
transform 1 0 492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1713453518
transform 1 0 308 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1713453518
transform 1 0 180 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1713453518
transform 1 0 116 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1713453518
transform 1 0 100 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1713453518
transform 1 0 92 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1713453518
transform 1 0 92 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1713453518
transform 1 0 92 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1713453518
transform 1 0 92 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1713453518
transform 1 0 84 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1713453518
transform 1 0 3364 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1713453518
transform 1 0 3292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1713453518
transform 1 0 3268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1713453518
transform 1 0 3164 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1713453518
transform 1 0 3052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1713453518
transform 1 0 2356 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1713453518
transform 1 0 2244 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1713453518
transform 1 0 1804 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1713453518
transform 1 0 1716 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1713453518
transform 1 0 1692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1713453518
transform 1 0 1588 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1713453518
transform 1 0 1580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1713453518
transform 1 0 1332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1713453518
transform 1 0 1316 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1713453518
transform 1 0 260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1713453518
transform 1 0 220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1713453518
transform 1 0 116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1713453518
transform 1 0 92 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1713453518
transform 1 0 1116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1713453518
transform 1 0 1108 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1713453518
transform 1 0 788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1713453518
transform 1 0 748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1713453518
transform 1 0 740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1713453518
transform 1 0 636 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1713453518
transform 1 0 612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1713453518
transform 1 0 588 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1713453518
transform 1 0 420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1713453518
transform 1 0 412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1713453518
transform 1 0 276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1713453518
transform 1 0 212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1713453518
transform 1 0 172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1713453518
transform 1 0 100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1713453518
transform 1 0 788 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1713453518
transform 1 0 788 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1713453518
transform 1 0 748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1713453518
transform 1 0 732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1713453518
transform 1 0 484 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1713453518
transform 1 0 332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1713453518
transform 1 0 332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1713453518
transform 1 0 324 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1713453518
transform 1 0 324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1713453518
transform 1 0 316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1713453518
transform 1 0 308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1713453518
transform 1 0 292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1713453518
transform 1 0 268 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1713453518
transform 1 0 260 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1713453518
transform 1 0 804 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1713453518
transform 1 0 724 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1713453518
transform 1 0 700 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1713453518
transform 1 0 700 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1713453518
transform 1 0 692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1713453518
transform 1 0 396 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1713453518
transform 1 0 380 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1713453518
transform 1 0 380 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1713453518
transform 1 0 372 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1713453518
transform 1 0 324 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1713453518
transform 1 0 324 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1713453518
transform 1 0 308 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1713453518
transform 1 0 292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1713453518
transform 1 0 284 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1713453518
transform 1 0 948 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1713453518
transform 1 0 948 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1713453518
transform 1 0 924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1713453518
transform 1 0 916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1713453518
transform 1 0 908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1713453518
transform 1 0 908 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1713453518
transform 1 0 908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1713453518
transform 1 0 900 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1713453518
transform 1 0 868 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1713453518
transform 1 0 852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1713453518
transform 1 0 852 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1713453518
transform 1 0 836 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1713453518
transform 1 0 828 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1713453518
transform 1 0 748 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1713453518
transform 1 0 996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1713453518
transform 1 0 956 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1713453518
transform 1 0 956 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1713453518
transform 1 0 956 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1713453518
transform 1 0 948 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1713453518
transform 1 0 948 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1713453518
transform 1 0 924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1713453518
transform 1 0 924 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1713453518
transform 1 0 916 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1713453518
transform 1 0 916 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1713453518
transform 1 0 908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1713453518
transform 1 0 900 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1713453518
transform 1 0 892 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1713453518
transform 1 0 868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1713453518
transform 1 0 3012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1713453518
transform 1 0 2932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1713453518
transform 1 0 2820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1713453518
transform 1 0 2684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1713453518
transform 1 0 2644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1713453518
transform 1 0 2492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1713453518
transform 1 0 2124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1713453518
transform 1 0 1020 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1713453518
transform 1 0 924 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1713453518
transform 1 0 892 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1713453518
transform 1 0 828 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1713453518
transform 1 0 804 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1713453518
transform 1 0 796 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1713453518
transform 1 0 748 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1713453518
transform 1 0 100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1713453518
transform 1 0 92 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1713453518
transform 1 0 732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1713453518
transform 1 0 724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1713453518
transform 1 0 716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1713453518
transform 1 0 708 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1713453518
transform 1 0 900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1713453518
transform 1 0 804 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1713453518
transform 1 0 804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1713453518
transform 1 0 732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1713453518
transform 1 0 796 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1713453518
transform 1 0 764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1713453518
transform 1 0 748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1713453518
transform 1 0 772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1713453518
transform 1 0 772 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1713453518
transform 1 0 764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1713453518
transform 1 0 756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1713453518
transform 1 0 732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1713453518
transform 1 0 716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1713453518
transform 1 0 708 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1713453518
transform 1 0 708 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1713453518
transform 1 0 708 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1713453518
transform 1 0 940 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1713453518
transform 1 0 932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1713453518
transform 1 0 908 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1713453518
transform 1 0 908 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1713453518
transform 1 0 876 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1713453518
transform 1 0 844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1713453518
transform 1 0 812 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1713453518
transform 1 0 796 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1713453518
transform 1 0 868 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1713453518
transform 1 0 852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1713453518
transform 1 0 852 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1713453518
transform 1 0 836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1713453518
transform 1 0 836 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1713453518
transform 1 0 836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1713453518
transform 1 0 804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1713453518
transform 1 0 804 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1713453518
transform 1 0 780 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1713453518
transform 1 0 836 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1713453518
transform 1 0 836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1713453518
transform 1 0 796 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1713453518
transform 1 0 796 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1713453518
transform 1 0 932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1713453518
transform 1 0 900 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1713453518
transform 1 0 900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1713453518
transform 1 0 876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1713453518
transform 1 0 860 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1713453518
transform 1 0 844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1713453518
transform 1 0 772 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1713453518
transform 1 0 772 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1713453518
transform 1 0 996 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1713453518
transform 1 0 948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1713453518
transform 1 0 948 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1713453518
transform 1 0 924 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1713453518
transform 1 0 924 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1713453518
transform 1 0 916 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1713453518
transform 1 0 916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1713453518
transform 1 0 908 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1713453518
transform 1 0 892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1713453518
transform 1 0 892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1713453518
transform 1 0 884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1713453518
transform 1 0 876 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1713453518
transform 1 0 868 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1713453518
transform 1 0 852 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1713453518
transform 1 0 852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1713453518
transform 1 0 852 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1713453518
transform 1 0 828 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1713453518
transform 1 0 820 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1713453518
transform 1 0 812 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1713453518
transform 1 0 796 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1713453518
transform 1 0 932 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1713453518
transform 1 0 892 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1713453518
transform 1 0 884 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1713453518
transform 1 0 860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1713453518
transform 1 0 836 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1713453518
transform 1 0 836 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1713453518
transform 1 0 796 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1713453518
transform 1 0 796 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1713453518
transform 1 0 796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1713453518
transform 1 0 796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1713453518
transform 1 0 788 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1713453518
transform 1 0 780 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1713453518
transform 1 0 780 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1713453518
transform 1 0 780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1713453518
transform 1 0 764 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1713453518
transform 1 0 748 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1713453518
transform 1 0 748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1713453518
transform 1 0 732 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1713453518
transform 1 0 724 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1713453518
transform 1 0 580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1713453518
transform 1 0 564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1713453518
transform 1 0 676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1713453518
transform 1 0 644 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1713453518
transform 1 0 628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1713453518
transform 1 0 572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1713453518
transform 1 0 444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1713453518
transform 1 0 396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1713453518
transform 1 0 324 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1713453518
transform 1 0 324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1713453518
transform 1 0 316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1713453518
transform 1 0 308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1713453518
transform 1 0 300 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1713453518
transform 1 0 292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1713453518
transform 1 0 284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1713453518
transform 1 0 284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1713453518
transform 1 0 284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1713453518
transform 1 0 276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1713453518
transform 1 0 276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1713453518
transform 1 0 268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1713453518
transform 1 0 244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1713453518
transform 1 0 204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1713453518
transform 1 0 132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1713453518
transform 1 0 124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1713453518
transform 1 0 524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1713453518
transform 1 0 508 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1713453518
transform 1 0 500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1713453518
transform 1 0 500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1713453518
transform 1 0 492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1713453518
transform 1 0 676 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1713453518
transform 1 0 676 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1713453518
transform 1 0 620 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1713453518
transform 1 0 612 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1713453518
transform 1 0 556 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1713453518
transform 1 0 556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1713453518
transform 1 0 532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1713453518
transform 1 0 524 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1713453518
transform 1 0 516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1713453518
transform 1 0 508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1713453518
transform 1 0 492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1713453518
transform 1 0 492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1713453518
transform 1 0 484 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1713453518
transform 1 0 484 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1713453518
transform 1 0 476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1713453518
transform 1 0 476 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1713453518
transform 1 0 476 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1713453518
transform 1 0 468 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1713453518
transform 1 0 460 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1713453518
transform 1 0 460 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1713453518
transform 1 0 452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1713453518
transform 1 0 452 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1713453518
transform 1 0 444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1713453518
transform 1 0 444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1713453518
transform 1 0 436 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1713453518
transform 1 0 420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1713453518
transform 1 0 404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1713453518
transform 1 0 404 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1713453518
transform 1 0 236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1713453518
transform 1 0 220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1713453518
transform 1 0 404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1713453518
transform 1 0 396 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1713453518
transform 1 0 348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1713453518
transform 1 0 332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1713453518
transform 1 0 332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1713453518
transform 1 0 252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1713453518
transform 1 0 236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1713453518
transform 1 0 236 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1713453518
transform 1 0 236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1713453518
transform 1 0 228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1713453518
transform 1 0 228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1713453518
transform 1 0 228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1713453518
transform 1 0 212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1713453518
transform 1 0 212 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1713453518
transform 1 0 212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1713453518
transform 1 0 212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1713453518
transform 1 0 204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1713453518
transform 1 0 148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1713453518
transform 1 0 140 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1713453518
transform 1 0 2212 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1713453518
transform 1 0 2188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1713453518
transform 1 0 2228 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1713453518
transform 1 0 2172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1713453518
transform 1 0 1932 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1713453518
transform 1 0 1652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1713453518
transform 1 0 1612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1713453518
transform 1 0 1548 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1713453518
transform 1 0 1508 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1713453518
transform 1 0 2388 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1713453518
transform 1 0 2340 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1713453518
transform 1 0 2332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1713453518
transform 1 0 2308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1713453518
transform 1 0 2276 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1713453518
transform 1 0 2204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1713453518
transform 1 0 2196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1713453518
transform 1 0 3380 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1713453518
transform 1 0 3380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1713453518
transform 1 0 3316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1713453518
transform 1 0 3236 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1713453518
transform 1 0 3196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1713453518
transform 1 0 3188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1713453518
transform 1 0 3124 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1713453518
transform 1 0 3108 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1713453518
transform 1 0 3092 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1713453518
transform 1 0 3092 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1713453518
transform 1 0 3084 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1713453518
transform 1 0 3084 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1713453518
transform 1 0 3076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1713453518
transform 1 0 3068 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1713453518
transform 1 0 2892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1713453518
transform 1 0 2884 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1713453518
transform 1 0 2884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1713453518
transform 1 0 2812 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1713453518
transform 1 0 2796 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1713453518
transform 1 0 2780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1713453518
transform 1 0 2756 0 1 1095
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1713453518
transform 1 0 2748 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1713453518
transform 1 0 2732 0 1 1095
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1713453518
transform 1 0 2732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1713453518
transform 1 0 2732 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1713453518
transform 1 0 2708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1713453518
transform 1 0 2684 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1713453518
transform 1 0 2668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1713453518
transform 1 0 2660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1713453518
transform 1 0 2644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1713453518
transform 1 0 2260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1713453518
transform 1 0 2220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1713453518
transform 1 0 2948 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1713453518
transform 1 0 2844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1713453518
transform 1 0 2780 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1713453518
transform 1 0 2716 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1713453518
transform 1 0 2716 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1713453518
transform 1 0 2660 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1713453518
transform 1 0 2604 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1713453518
transform 1 0 2604 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1713453518
transform 1 0 2508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1713453518
transform 1 0 2500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1713453518
transform 1 0 2500 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1713453518
transform 1 0 2484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1713453518
transform 1 0 2476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1713453518
transform 1 0 2468 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1713453518
transform 1 0 2428 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1713453518
transform 1 0 2420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1713453518
transform 1 0 2412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1713453518
transform 1 0 2404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1713453518
transform 1 0 2404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1713453518
transform 1 0 2356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1713453518
transform 1 0 2348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1713453518
transform 1 0 2332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1713453518
transform 1 0 2332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1713453518
transform 1 0 2324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1713453518
transform 1 0 2324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1713453518
transform 1 0 2300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1713453518
transform 1 0 2292 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1713453518
transform 1 0 2292 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1713453518
transform 1 0 2292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1713453518
transform 1 0 2284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1713453518
transform 1 0 2284 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1713453518
transform 1 0 2284 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1713453518
transform 1 0 2284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1713453518
transform 1 0 3404 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1713453518
transform 1 0 3372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1713453518
transform 1 0 3300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1713453518
transform 1 0 3292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1713453518
transform 1 0 3084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1713453518
transform 1 0 2996 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1713453518
transform 1 0 2988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1713453518
transform 1 0 2988 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1713453518
transform 1 0 2988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1713453518
transform 1 0 2964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1713453518
transform 1 0 2948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1713453518
transform 1 0 2884 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1713453518
transform 1 0 2876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1713453518
transform 1 0 2860 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1713453518
transform 1 0 2820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1713453518
transform 1 0 3436 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1713453518
transform 1 0 3436 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1713453518
transform 1 0 3428 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1713453518
transform 1 0 3428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1713453518
transform 1 0 3404 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1713453518
transform 1 0 3380 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1713453518
transform 1 0 3356 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1713453518
transform 1 0 3332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1713453518
transform 1 0 3268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1713453518
transform 1 0 3164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1713453518
transform 1 0 3164 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1713453518
transform 1 0 3028 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1713453518
transform 1 0 3012 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1713453518
transform 1 0 3404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1713453518
transform 1 0 3396 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1713453518
transform 1 0 3388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1713453518
transform 1 0 3388 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1713453518
transform 1 0 3372 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1713453518
transform 1 0 3348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1713453518
transform 1 0 3340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1713453518
transform 1 0 3332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1713453518
transform 1 0 3316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1713453518
transform 1 0 3308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1713453518
transform 1 0 3300 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1713453518
transform 1 0 3244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1713453518
transform 1 0 3236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1713453518
transform 1 0 3100 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1713453518
transform 1 0 3084 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1713453518
transform 1 0 3084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1713453518
transform 1 0 3044 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1713453518
transform 1 0 2972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1713453518
transform 1 0 2972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1713453518
transform 1 0 2940 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1713453518
transform 1 0 2940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1713453518
transform 1 0 2932 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1713453518
transform 1 0 2924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1713453518
transform 1 0 2916 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1713453518
transform 1 0 2804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1713453518
transform 1 0 2804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1713453518
transform 1 0 2804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1713453518
transform 1 0 3260 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1713453518
transform 1 0 3236 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1713453518
transform 1 0 3236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1713453518
transform 1 0 3236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1713453518
transform 1 0 3204 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1713453518
transform 1 0 3196 0 1 1613
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1713453518
transform 1 0 3188 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1713453518
transform 1 0 3188 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1713453518
transform 1 0 3172 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1713453518
transform 1 0 3164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1713453518
transform 1 0 3164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1713453518
transform 1 0 3132 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1713453518
transform 1 0 3116 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1713453518
transform 1 0 3116 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1713453518
transform 1 0 3068 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1713453518
transform 1 0 3068 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1713453518
transform 1 0 3036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1713453518
transform 1 0 2988 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1713453518
transform 1 0 2980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1713453518
transform 1 0 2940 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1713453518
transform 1 0 2844 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1713453518
transform 1 0 2836 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1713453518
transform 1 0 2828 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1713453518
transform 1 0 2820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1713453518
transform 1 0 2788 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1713453518
transform 1 0 2788 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1713453518
transform 1 0 2740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1713453518
transform 1 0 2724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1713453518
transform 1 0 2716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1713453518
transform 1 0 2684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1713453518
transform 1 0 2676 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1713453518
transform 1 0 2652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1713453518
transform 1 0 2876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1713453518
transform 1 0 2780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1713453518
transform 1 0 2580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1713453518
transform 1 0 2556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1713453518
transform 1 0 2956 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1713453518
transform 1 0 2588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1713453518
transform 1 0 2452 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1713453518
transform 1 0 2276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1713453518
transform 1 0 2596 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1713453518
transform 1 0 2564 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1713453518
transform 1 0 2564 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1713453518
transform 1 0 2564 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1713453518
transform 1 0 2540 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1713453518
transform 1 0 2540 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1713453518
transform 1 0 2516 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1713453518
transform 1 0 2420 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1713453518
transform 1 0 2420 0 1 555
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1713453518
transform 1 0 2412 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1713453518
transform 1 0 2372 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1713453518
transform 1 0 2372 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1713453518
transform 1 0 2348 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1713453518
transform 1 0 2308 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1713453518
transform 1 0 2268 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1713453518
transform 1 0 2212 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1713453518
transform 1 0 2212 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1713453518
transform 1 0 2204 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1713453518
transform 1 0 2092 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1713453518
transform 1 0 2084 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1713453518
transform 1 0 2076 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1713453518
transform 1 0 2020 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1713453518
transform 1 0 2012 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1713453518
transform 1 0 1964 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1713453518
transform 1 0 1932 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1713453518
transform 1 0 1916 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1713453518
transform 1 0 1908 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1713453518
transform 1 0 1892 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1713453518
transform 1 0 1892 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1713453518
transform 1 0 1892 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1713453518
transform 1 0 1884 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1713453518
transform 1 0 1884 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1713453518
transform 1 0 1860 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1713453518
transform 1 0 1844 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1713453518
transform 1 0 1844 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1713453518
transform 1 0 1828 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1713453518
transform 1 0 1820 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1713453518
transform 1 0 1532 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1713453518
transform 1 0 1508 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1713453518
transform 1 0 1476 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1713453518
transform 1 0 2404 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1713453518
transform 1 0 2388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1713453518
transform 1 0 2388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1713453518
transform 1 0 2332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1713453518
transform 1 0 2164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1713453518
transform 1 0 2156 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1713453518
transform 1 0 2156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1713453518
transform 1 0 2116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1713453518
transform 1 0 2060 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1713453518
transform 1 0 2012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1713453518
transform 1 0 1972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1713453518
transform 1 0 1940 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1713453518
transform 1 0 1940 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1713453518
transform 1 0 1868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1713453518
transform 1 0 2180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1713453518
transform 1 0 2172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1713453518
transform 1 0 2172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1713453518
transform 1 0 2164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1713453518
transform 1 0 2164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1713453518
transform 1 0 2140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1713453518
transform 1 0 2124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1713453518
transform 1 0 2100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1713453518
transform 1 0 2100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1713453518
transform 1 0 2036 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1713453518
transform 1 0 2020 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1713453518
transform 1 0 1932 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1713453518
transform 1 0 1892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1713453518
transform 1 0 1868 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1713453518
transform 1 0 2340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1713453518
transform 1 0 2300 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1713453518
transform 1 0 2300 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1713453518
transform 1 0 2252 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1713453518
transform 1 0 2124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1713453518
transform 1 0 2116 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1713453518
transform 1 0 2084 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1713453518
transform 1 0 2084 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1713453518
transform 1 0 2084 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1713453518
transform 1 0 2076 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1713453518
transform 1 0 1988 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1713453518
transform 1 0 1988 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1713453518
transform 1 0 1980 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1713453518
transform 1 0 1972 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1713453518
transform 1 0 1932 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1713453518
transform 1 0 1924 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1713453518
transform 1 0 1908 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1713453518
transform 1 0 1908 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1713453518
transform 1 0 2132 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1713453518
transform 1 0 2132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1713453518
transform 1 0 2124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1713453518
transform 1 0 2116 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1713453518
transform 1 0 2084 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1713453518
transform 1 0 2044 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1713453518
transform 1 0 2028 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1713453518
transform 1 0 2028 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1713453518
transform 1 0 2028 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1713453518
transform 1 0 1996 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1713453518
transform 1 0 1964 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1713453518
transform 1 0 1964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1713453518
transform 1 0 1900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1713453518
transform 1 0 1868 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1713453518
transform 1 0 1804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1713453518
transform 1 0 1764 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1713453518
transform 1 0 1732 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1713453518
transform 1 0 1644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1713453518
transform 1 0 1540 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1713453518
transform 1 0 2548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1713453518
transform 1 0 2532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1713453518
transform 1 0 2516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1713453518
transform 1 0 2468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1713453518
transform 1 0 2428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1713453518
transform 1 0 2404 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1713453518
transform 1 0 2380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1713453518
transform 1 0 2364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1713453518
transform 1 0 2364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1713453518
transform 1 0 2364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1713453518
transform 1 0 2364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1713453518
transform 1 0 2356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1713453518
transform 1 0 2348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1713453518
transform 1 0 2236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1713453518
transform 1 0 2236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1713453518
transform 1 0 2236 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1713453518
transform 1 0 2228 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1713453518
transform 1 0 2188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1713453518
transform 1 0 2188 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1713453518
transform 1 0 2764 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1713453518
transform 1 0 2748 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1713453518
transform 1 0 2724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1713453518
transform 1 0 2668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1713453518
transform 1 0 2668 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1713453518
transform 1 0 2644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1713453518
transform 1 0 2644 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1713453518
transform 1 0 2620 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1713453518
transform 1 0 2588 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1713453518
transform 1 0 2540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1713453518
transform 1 0 2484 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1713453518
transform 1 0 2476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1713453518
transform 1 0 2476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1713453518
transform 1 0 2380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1713453518
transform 1 0 2380 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1713453518
transform 1 0 2332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1713453518
transform 1 0 2332 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1713453518
transform 1 0 2236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1713453518
transform 1 0 1708 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1713453518
transform 1 0 1660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1713453518
transform 1 0 1620 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1713453518
transform 1 0 1604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1713453518
transform 1 0 1580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1713453518
transform 1 0 1572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1713453518
transform 1 0 1572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1713453518
transform 1 0 1548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1713453518
transform 1 0 1524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1713453518
transform 1 0 1404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1713453518
transform 1 0 1372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1713453518
transform 1 0 1500 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1713453518
transform 1 0 1500 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1713453518
transform 1 0 1492 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1713453518
transform 1 0 1492 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1713453518
transform 1 0 1476 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1713453518
transform 1 0 1468 0 1 1003
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1713453518
transform 1 0 1372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1713453518
transform 1 0 1372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1713453518
transform 1 0 1372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1713453518
transform 1 0 1348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1713453518
transform 1 0 1348 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1713453518
transform 1 0 1348 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1713453518
transform 1 0 1292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1713453518
transform 1 0 1724 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1713453518
transform 1 0 1692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1713453518
transform 1 0 1652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1713453518
transform 1 0 1580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1713453518
transform 1 0 1564 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1713453518
transform 1 0 1556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1713453518
transform 1 0 1556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1713453518
transform 1 0 1500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1713453518
transform 1 0 1468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1713453518
transform 1 0 1460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1713453518
transform 1 0 1452 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1713453518
transform 1 0 1692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1713453518
transform 1 0 1652 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1713453518
transform 1 0 1644 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1713453518
transform 1 0 1636 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1713453518
transform 1 0 1628 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1713453518
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1713453518
transform 1 0 1620 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1713453518
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1713453518
transform 1 0 1588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1713453518
transform 1 0 1572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1713453518
transform 1 0 1564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1713453518
transform 1 0 1548 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1713453518
transform 1 0 1540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1713453518
transform 1 0 1524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1713453518
transform 1 0 1524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1713453518
transform 1 0 1500 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1713453518
transform 1 0 1492 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1713453518
transform 1 0 1444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1713453518
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1713453518
transform 1 0 1428 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1713453518
transform 1 0 1428 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1713453518
transform 1 0 1412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1713453518
transform 1 0 1396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1713453518
transform 1 0 1396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1713453518
transform 1 0 1372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1713453518
transform 1 0 1364 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1713453518
transform 1 0 1316 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1713453518
transform 1 0 1300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1713453518
transform 1 0 2852 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1713453518
transform 1 0 2820 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1713453518
transform 1 0 2412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1713453518
transform 1 0 1108 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1713453518
transform 1 0 1084 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1713453518
transform 1 0 1076 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1713453518
transform 1 0 1052 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1713453518
transform 1 0 1044 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1713453518
transform 1 0 1044 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1713453518
transform 1 0 1044 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1713453518
transform 1 0 1044 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1713453518
transform 1 0 1036 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1713453518
transform 1 0 1036 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1713453518
transform 1 0 1020 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1713453518
transform 1 0 1020 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1713453518
transform 1 0 1012 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1713453518
transform 1 0 988 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1713453518
transform 1 0 884 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1713453518
transform 1 0 868 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1713453518
transform 1 0 1068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1713453518
transform 1 0 1060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1713453518
transform 1 0 1060 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1713453518
transform 1 0 1060 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1713453518
transform 1 0 1044 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1713453518
transform 1 0 1012 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1713453518
transform 1 0 1012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1713453518
transform 1 0 1012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1713453518
transform 1 0 1004 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1713453518
transform 1 0 1004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1713453518
transform 1 0 1004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1713453518
transform 1 0 996 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1713453518
transform 1 0 988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1713453518
transform 1 0 972 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1713453518
transform 1 0 964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1713453518
transform 1 0 2932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1713453518
transform 1 0 2884 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1713453518
transform 1 0 2828 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1713453518
transform 1 0 2756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1713453518
transform 1 0 2732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1713453518
transform 1 0 2428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1713453518
transform 1 0 2252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1713453518
transform 1 0 1364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1713453518
transform 1 0 1060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1713453518
transform 1 0 1012 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1713453518
transform 1 0 1012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1713453518
transform 1 0 964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1713453518
transform 1 0 892 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1713453518
transform 1 0 852 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1713453518
transform 1 0 620 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1713453518
transform 1 0 612 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1713453518
transform 1 0 572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1713453518
transform 1 0 516 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1713453518
transform 1 0 516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1713453518
transform 1 0 484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1713453518
transform 1 0 484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1713453518
transform 1 0 484 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1713453518
transform 1 0 444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1713453518
transform 1 0 428 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1713453518
transform 1 0 412 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1713453518
transform 1 0 404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1713453518
transform 1 0 396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1713453518
transform 1 0 388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1713453518
transform 1 0 500 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1713453518
transform 1 0 460 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1713453518
transform 1 0 444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1713453518
transform 1 0 444 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1713453518
transform 1 0 444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1713453518
transform 1 0 444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1713453518
transform 1 0 420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1713453518
transform 1 0 420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1713453518
transform 1 0 396 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1713453518
transform 1 0 388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1713453518
transform 1 0 388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1713453518
transform 1 0 372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1713453518
transform 1 0 372 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1713453518
transform 1 0 356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1713453518
transform 1 0 356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1713453518
transform 1 0 332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1713453518
transform 1 0 300 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1713453518
transform 1 0 2732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1713453518
transform 1 0 2724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1713453518
transform 1 0 2660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1713453518
transform 1 0 2628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1713453518
transform 1 0 2444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1713453518
transform 1 0 2300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1713453518
transform 1 0 2276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1713453518
transform 1 0 2180 0 1 2985
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1713453518
transform 1 0 2172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1713453518
transform 1 0 2124 0 1 2985
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1713453518
transform 1 0 2116 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1713453518
transform 1 0 1892 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1713453518
transform 1 0 1660 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1713453518
transform 1 0 1644 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1713453518
transform 1 0 3428 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1713453518
transform 1 0 3388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1713453518
transform 1 0 3388 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1713453518
transform 1 0 3380 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1713453518
transform 1 0 3364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1713453518
transform 1 0 3324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1713453518
transform 1 0 3268 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1713453518
transform 1 0 3220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1713453518
transform 1 0 3164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1713453518
transform 1 0 3148 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1713453518
transform 1 0 3148 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1713453518
transform 1 0 1812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1713453518
transform 1 0 1788 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1713453518
transform 1 0 1788 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1713453518
transform 1 0 1772 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1713453518
transform 1 0 1732 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1713453518
transform 1 0 1724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1713453518
transform 1 0 1716 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1713453518
transform 1 0 1548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1713453518
transform 1 0 1444 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1713453518
transform 1 0 1444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1713453518
transform 1 0 1500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1713453518
transform 1 0 1444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1713453518
transform 1 0 1444 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1713453518
transform 1 0 1436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1713453518
transform 1 0 1428 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1713453518
transform 1 0 1420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1713453518
transform 1 0 1412 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1713453518
transform 1 0 1396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1713453518
transform 1 0 1356 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1713453518
transform 1 0 1332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1713453518
transform 1 0 1332 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1713453518
transform 1 0 1332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1713453518
transform 1 0 1316 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1713453518
transform 1 0 1228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1713453518
transform 1 0 1212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1713453518
transform 1 0 1196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1713453518
transform 1 0 1196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1713453518
transform 1 0 1188 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1713453518
transform 1 0 1180 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1713453518
transform 1 0 1180 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1713453518
transform 1 0 1172 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1713453518
transform 1 0 1156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1713453518
transform 1 0 1140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1713453518
transform 1 0 1516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1713453518
transform 1 0 1500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1713453518
transform 1 0 1484 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1713453518
transform 1 0 1468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1713453518
transform 1 0 1460 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1713453518
transform 1 0 1460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1713453518
transform 1 0 1428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1713453518
transform 1 0 1380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1713453518
transform 1 0 1356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1713453518
transform 1 0 1348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1713453518
transform 1 0 1300 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1713453518
transform 1 0 1244 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1713453518
transform 1 0 1212 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1713453518
transform 1 0 1196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1713453518
transform 1 0 1188 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1713453518
transform 1 0 2892 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1713453518
transform 1 0 2828 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1713453518
transform 1 0 2764 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1713453518
transform 1 0 2668 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1713453518
transform 1 0 2492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1713453518
transform 1 0 2404 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1713453518
transform 1 0 2388 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1713453518
transform 1 0 2300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1713453518
transform 1 0 2284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1713453518
transform 1 0 2236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1713453518
transform 1 0 2212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1713453518
transform 1 0 1404 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1713453518
transform 1 0 1404 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1713453518
transform 1 0 1364 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1713453518
transform 1 0 1356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1713453518
transform 1 0 1356 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1713453518
transform 1 0 1348 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1713453518
transform 1 0 1324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1713453518
transform 1 0 1324 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1713453518
transform 1 0 1324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1713453518
transform 1 0 1308 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1713453518
transform 1 0 1268 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1713453518
transform 1 0 1236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1713453518
transform 1 0 1228 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1713453518
transform 1 0 1116 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1713453518
transform 1 0 3364 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1713453518
transform 1 0 3324 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1713453518
transform 1 0 3300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1713453518
transform 1 0 3284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1713453518
transform 1 0 2788 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1713453518
transform 1 0 2716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1713453518
transform 1 0 2580 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1713453518
transform 1 0 2572 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1713453518
transform 1 0 2556 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1713453518
transform 1 0 2540 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1713453518
transform 1 0 2460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1713453518
transform 1 0 2420 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1713453518
transform 1 0 1812 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1713453518
transform 1 0 3420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1713453518
transform 1 0 3412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1713453518
transform 1 0 3196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1713453518
transform 1 0 3012 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1713453518
transform 1 0 2748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1713453518
transform 1 0 2740 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1713453518
transform 1 0 2588 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1713453518
transform 1 0 2484 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1713453518
transform 1 0 2388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1713453518
transform 1 0 2388 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1713453518
transform 1 0 1868 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1713453518
transform 1 0 3404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1713453518
transform 1 0 2900 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1713453518
transform 1 0 2796 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1713453518
transform 1 0 2756 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1713453518
transform 1 0 2716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1713453518
transform 1 0 2620 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1713453518
transform 1 0 2612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1713453518
transform 1 0 2604 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1713453518
transform 1 0 2604 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1713453518
transform 1 0 2572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1713453518
transform 1 0 2483 0 1 1414
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1713453518
transform 1 0 2452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1713453518
transform 1 0 2780 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1713453518
transform 1 0 2772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1713453518
transform 1 0 2740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1713453518
transform 1 0 2740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1713453518
transform 1 0 2628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1713453518
transform 1 0 2572 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1713453518
transform 1 0 2228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1713453518
transform 1 0 1132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1713453518
transform 1 0 1108 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1713453518
transform 1 0 1076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1713453518
transform 1 0 1068 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1713453518
transform 1 0 1068 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1713453518
transform 1 0 1068 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1713453518
transform 1 0 1052 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1713453518
transform 1 0 1044 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1713453518
transform 1 0 1028 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1713453518
transform 1 0 2956 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1713453518
transform 1 0 2876 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1713453518
transform 1 0 2852 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1713453518
transform 1 0 2652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1713453518
transform 1 0 2212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1713453518
transform 1 0 3372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1713453518
transform 1 0 3372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1713453518
transform 1 0 3332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1713453518
transform 1 0 3220 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1713453518
transform 1 0 3204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1713453518
transform 1 0 3084 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1713453518
transform 1 0 2916 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1713453518
transform 1 0 2828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1713453518
transform 1 0 2636 0 1 1885
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1713453518
transform 1 0 2612 0 1 1885
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1713453518
transform 1 0 2572 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1713453518
transform 1 0 2540 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1713453518
transform 1 0 2444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1713453518
transform 1 0 1700 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1713453518
transform 1 0 3404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1713453518
transform 1 0 3332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1713453518
transform 1 0 3292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1713453518
transform 1 0 3180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1713453518
transform 1 0 2980 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1713453518
transform 1 0 2932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1713453518
transform 1 0 2700 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1713453518
transform 1 0 2684 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1713453518
transform 1 0 2652 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1713453518
transform 1 0 2468 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1713453518
transform 1 0 1836 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1713453518
transform 1 0 3276 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1713453518
transform 1 0 3276 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1713453518
transform 1 0 3140 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1713453518
transform 1 0 3044 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1713453518
transform 1 0 3012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1713453518
transform 1 0 2948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1713453518
transform 1 0 2764 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1713453518
transform 1 0 2572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1713453518
transform 1 0 2380 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1713453518
transform 1 0 1652 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1713453518
transform 1 0 3140 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1713453518
transform 1 0 3076 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1713453518
transform 1 0 2956 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1713453518
transform 1 0 2924 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1713453518
transform 1 0 2908 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1713453518
transform 1 0 2892 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1713453518
transform 1 0 2796 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1713453518
transform 1 0 2692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1713453518
transform 1 0 2412 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1713453518
transform 1 0 2140 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1713453518
transform 1 0 1900 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1713453518
transform 1 0 1300 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1713453518
transform 1 0 2836 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1713453518
transform 1 0 2772 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1713453518
transform 1 0 2684 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1713453518
transform 1 0 2556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1713453518
transform 1 0 2172 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1713453518
transform 1 0 1236 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1713453518
transform 1 0 1188 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1713453518
transform 1 0 1148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1713453518
transform 1 0 1084 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1713453518
transform 1 0 1076 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1713453518
transform 1 0 1068 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1713453518
transform 1 0 1052 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1713453518
transform 1 0 1036 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1713453518
transform 1 0 1020 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1713453518
transform 1 0 3124 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1713453518
transform 1 0 3076 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1713453518
transform 1 0 3044 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1713453518
transform 1 0 2996 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1713453518
transform 1 0 2724 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1713453518
transform 1 0 2428 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1713453518
transform 1 0 1948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1713453518
transform 1 0 1732 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1713453518
transform 1 0 1676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1713453518
transform 1 0 1668 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1713453518
transform 1 0 1644 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1713453518
transform 1 0 1524 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1713453518
transform 1 0 2188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1713453518
transform 1 0 2188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1713453518
transform 1 0 2180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1713453518
transform 1 0 2164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1713453518
transform 1 0 2156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1713453518
transform 1 0 2556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1713453518
transform 1 0 2540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1713453518
transform 1 0 2540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1713453518
transform 1 0 1428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1713453518
transform 1 0 524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1713453518
transform 1 0 476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1713453518
transform 1 0 1580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1713453518
transform 1 0 1532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1713453518
transform 1 0 1492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1713453518
transform 1 0 1324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1713453518
transform 1 0 1324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1713453518
transform 1 0 1292 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1713453518
transform 1 0 2660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1713453518
transform 1 0 2644 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1713453518
transform 1 0 2796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1713453518
transform 1 0 2716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1713453518
transform 1 0 3436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1713453518
transform 1 0 3404 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1713453518
transform 1 0 3100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1713453518
transform 1 0 3068 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1713453518
transform 1 0 2980 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1713453518
transform 1 0 2436 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1713453518
transform 1 0 2084 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1713453518
transform 1 0 3156 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1713453518
transform 1 0 3036 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1713453518
transform 1 0 2740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1713453518
transform 1 0 2676 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1713453518
transform 1 0 2300 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1713453518
transform 1 0 3100 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1713453518
transform 1 0 2940 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1713453518
transform 1 0 2900 0 1 2645
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1713453518
transform 1 0 2892 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1713453518
transform 1 0 2668 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1713453518
transform 1 0 2332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1713453518
transform 1 0 2324 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1713453518
transform 1 0 3212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1713453518
transform 1 0 3180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1713453518
transform 1 0 3172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1713453518
transform 1 0 3156 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1713453518
transform 1 0 2868 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1713453518
transform 1 0 2484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1713453518
transform 1 0 2204 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1713453518
transform 1 0 2156 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1713453518
transform 1 0 3372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1713453518
transform 1 0 3324 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1713453518
transform 1 0 3324 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1713453518
transform 1 0 3076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1713453518
transform 1 0 2228 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1713453518
transform 1 0 2196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1713453518
transform 1 0 3284 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1713453518
transform 1 0 3284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1713453518
transform 1 0 2804 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1713453518
transform 1 0 2644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1713453518
transform 1 0 2180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1713453518
transform 1 0 3420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1713453518
transform 1 0 3412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1713453518
transform 1 0 3300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1713453518
transform 1 0 3188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1713453518
transform 1 0 2908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1713453518
transform 1 0 2196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1713453518
transform 1 0 3372 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1713453518
transform 1 0 3364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1713453518
transform 1 0 3324 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1713453518
transform 1 0 3260 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1713453518
transform 1 0 3020 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1713453518
transform 1 0 2236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1713453518
transform 1 0 2172 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1713453518
transform 1 0 2164 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1713453518
transform 1 0 2156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1713453518
transform 1 0 2148 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1713453518
transform 1 0 2068 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1713453518
transform 1 0 2044 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1713453518
transform 1 0 2020 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1713453518
transform 1 0 1644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1713453518
transform 1 0 1380 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1713453518
transform 1 0 1316 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1713453518
transform 1 0 1284 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1713453518
transform 1 0 1284 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1713453518
transform 1 0 1276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1713453518
transform 1 0 1276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1713453518
transform 1 0 1220 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1713453518
transform 1 0 1212 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1713453518
transform 1 0 1204 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1713453518
transform 1 0 1180 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1713453518
transform 1 0 1124 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1713453518
transform 1 0 1092 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1713453518
transform 1 0 1076 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1713453518
transform 1 0 1404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1713453518
transform 1 0 1380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1713453518
transform 1 0 1372 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1713453518
transform 1 0 1356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1713453518
transform 1 0 1284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1713453518
transform 1 0 1268 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1713453518
transform 1 0 1268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1713453518
transform 1 0 1228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1713453518
transform 1 0 1180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1713453518
transform 1 0 1180 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1713453518
transform 1 0 1172 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1713453518
transform 1 0 1148 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1713453518
transform 1 0 1140 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1713453518
transform 1 0 1124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1713453518
transform 1 0 1916 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1713453518
transform 1 0 1876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1713453518
transform 1 0 1844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1713453518
transform 1 0 1812 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1713453518
transform 1 0 1492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1713453518
transform 1 0 3356 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1713453518
transform 1 0 3356 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1713453518
transform 1 0 3348 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1713453518
transform 1 0 3196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1713453518
transform 1 0 2676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1713453518
transform 1 0 2164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1713453518
transform 1 0 1556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1713453518
transform 1 0 1516 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1713453518
transform 1 0 1388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1713453518
transform 1 0 1332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1713453518
transform 1 0 1308 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1713453518
transform 1 0 1276 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1713453518
transform 1 0 1196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1713453518
transform 1 0 1188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1713453518
transform 1 0 1172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1713453518
transform 1 0 1156 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1713453518
transform 1 0 1140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1713453518
transform 1 0 1132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1713453518
transform 1 0 1116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1713453518
transform 1 0 1116 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1713453518
transform 1 0 1108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1713453518
transform 1 0 2044 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1713453518
transform 1 0 1948 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1713453518
transform 1 0 1844 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1713453518
transform 1 0 1972 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1713453518
transform 1 0 1884 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1713453518
transform 1 0 1724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1713453518
transform 1 0 2740 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1713453518
transform 1 0 2700 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1713453518
transform 1 0 2628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1713453518
transform 1 0 2588 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1713453518
transform 1 0 2732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1713453518
transform 1 0 2660 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1713453518
transform 1 0 2916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1713453518
transform 1 0 2876 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1713453518
transform 1 0 3044 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1713453518
transform 1 0 2948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1713453518
transform 1 0 3388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1713453518
transform 1 0 3140 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1713453518
transform 1 0 3076 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1713453518
transform 1 0 2692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1713453518
transform 1 0 3292 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1713453518
transform 1 0 2788 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1713453518
transform 1 0 3316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1713453518
transform 1 0 3020 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1713453518
transform 1 0 3188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1713453518
transform 1 0 3188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1713453518
transform 1 0 2268 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1713453518
transform 1 0 2236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1713453518
transform 1 0 2380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1713453518
transform 1 0 2380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1713453518
transform 1 0 3444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1713453518
transform 1 0 3412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1713453518
transform 1 0 3396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1713453518
transform 1 0 3420 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1713453518
transform 1 0 3252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1713453518
transform 1 0 3380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1713453518
transform 1 0 3356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1713453518
transform 1 0 3412 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1713453518
transform 1 0 3388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1713453518
transform 1 0 3348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1713453518
transform 1 0 3324 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1713453518
transform 1 0 3284 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1713453518
transform 1 0 3204 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1713453518
transform 1 0 2836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1713453518
transform 1 0 3348 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1713453518
transform 1 0 3316 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1713453518
transform 1 0 3308 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1713453518
transform 1 0 3300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1713453518
transform 1 0 3212 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1713453518
transform 1 0 3196 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1713453518
transform 1 0 3412 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1713453518
transform 1 0 3412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1713453518
transform 1 0 3372 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1713453518
transform 1 0 3372 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1713453518
transform 1 0 3316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1713453518
transform 1 0 3196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1713453518
transform 1 0 3028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1713453518
transform 1 0 2804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1713453518
transform 1 0 3244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1713453518
transform 1 0 3180 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1713453518
transform 1 0 3132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1713453518
transform 1 0 3020 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1713453518
transform 1 0 3020 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1713453518
transform 1 0 3348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1713453518
transform 1 0 3204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1713453518
transform 1 0 3188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1713453518
transform 1 0 3084 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1713453518
transform 1 0 3012 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1713453518
transform 1 0 2924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1713453518
transform 1 0 2868 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1713453518
transform 1 0 2772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1713453518
transform 1 0 2732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1713453518
transform 1 0 2780 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1713453518
transform 1 0 2692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1713453518
transform 1 0 2956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1713453518
transform 1 0 2868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1713453518
transform 1 0 3036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1713453518
transform 1 0 2948 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1713453518
transform 1 0 2268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1713453518
transform 1 0 2172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1713453518
transform 1 0 2516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1713453518
transform 1 0 2444 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1713453518
transform 1 0 884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1713453518
transform 1 0 796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1713453518
transform 1 0 1036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1713453518
transform 1 0 956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1713453518
transform 1 0 1084 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1713453518
transform 1 0 988 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1713453518
transform 1 0 1052 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1713453518
transform 1 0 964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1713453518
transform 1 0 988 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1713453518
transform 1 0 900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1713453518
transform 1 0 1036 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1713453518
transform 1 0 956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1713453518
transform 1 0 1044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1713453518
transform 1 0 940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1713453518
transform 1 0 1020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1713453518
transform 1 0 900 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1713453518
transform 1 0 1092 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1713453518
transform 1 0 964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1713453518
transform 1 0 988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1713453518
transform 1 0 876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1713453518
transform 1 0 1084 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1713453518
transform 1 0 988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1713453518
transform 1 0 1012 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1713453518
transform 1 0 916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1713453518
transform 1 0 1052 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1713453518
transform 1 0 956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1713453518
transform 1 0 1028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1713453518
transform 1 0 1004 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1713453518
transform 1 0 1092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1713453518
transform 1 0 1004 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1713453518
transform 1 0 1084 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1713453518
transform 1 0 964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1713453518
transform 1 0 1052 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1713453518
transform 1 0 956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1713453518
transform 1 0 1028 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1713453518
transform 1 0 940 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1713453518
transform 1 0 1012 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1713453518
transform 1 0 916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1713453518
transform 1 0 1068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1713453518
transform 1 0 972 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1713453518
transform 1 0 1092 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1713453518
transform 1 0 996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1713453518
transform 1 0 1044 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1713453518
transform 1 0 948 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1713453518
transform 1 0 1052 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1713453518
transform 1 0 964 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1713453518
transform 1 0 1092 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1713453518
transform 1 0 1004 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1713453518
transform 1 0 1068 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1713453518
transform 1 0 996 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1713453518
transform 1 0 1124 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1713453518
transform 1 0 1036 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1713453518
transform 1 0 1148 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1713453518
transform 1 0 1068 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1713453518
transform 1 0 1100 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1713453518
transform 1 0 956 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1713453518
transform 1 0 1068 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1713453518
transform 1 0 940 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1713453518
transform 1 0 908 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1713453518
transform 1 0 844 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1713453518
transform 1 0 892 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1713453518
transform 1 0 796 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1713453518
transform 1 0 916 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1713453518
transform 1 0 852 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1713453518
transform 1 0 1052 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1713453518
transform 1 0 852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1713453518
transform 1 0 3068 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1713453518
transform 1 0 3020 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1713453518
transform 1 0 2220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1713453518
transform 1 0 2220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1713453518
transform 1 0 2172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1713453518
transform 1 0 2156 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1713453518
transform 1 0 3100 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1713453518
transform 1 0 3100 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1713453518
transform 1 0 2980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1713453518
transform 1 0 2732 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1713453518
transform 1 0 2636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1713453518
transform 1 0 2468 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1713453518
transform 1 0 2132 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1713453518
transform 1 0 2116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1713453518
transform 1 0 2068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1713453518
transform 1 0 1924 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1713453518
transform 1 0 1796 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1713453518
transform 1 0 1740 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1713453518
transform 1 0 1516 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1713453518
transform 1 0 1476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1713453518
transform 1 0 1460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1713453518
transform 1 0 1620 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1713453518
transform 1 0 1532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1713453518
transform 1 0 1468 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1713453518
transform 1 0 636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1713453518
transform 1 0 412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1713453518
transform 1 0 348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1713453518
transform 1 0 236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1713453518
transform 1 0 2764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1713453518
transform 1 0 2764 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1713453518
transform 1 0 2748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1713453518
transform 1 0 2732 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1713453518
transform 1 0 2724 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1713453518
transform 1 0 2692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1713453518
transform 1 0 2684 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1713453518
transform 1 0 2028 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1713453518
transform 1 0 1044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1713453518
transform 1 0 2988 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1713453518
transform 1 0 1988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1713453518
transform 1 0 2084 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1713453518
transform 1 0 1996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1713453518
transform 1 0 2012 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1713453518
transform 1 0 1964 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1713453518
transform 1 0 2252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1713453518
transform 1 0 2052 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1713453518
transform 1 0 2316 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1713453518
transform 1 0 2244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1713453518
transform 1 0 2692 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1713453518
transform 1 0 2340 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1713453518
transform 1 0 2716 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1713453518
transform 1 0 2652 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1713453518
transform 1 0 2644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1713453518
transform 1 0 2628 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1713453518
transform 1 0 2700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1713453518
transform 1 0 2668 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1713453518
transform 1 0 2732 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1713453518
transform 1 0 2708 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1713453518
transform 1 0 2756 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1713453518
transform 1 0 2748 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1713453518
transform 1 0 2660 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1713453518
transform 1 0 2332 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1713453518
transform 1 0 3028 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1713453518
transform 1 0 2740 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1713453518
transform 1 0 2660 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1713453518
transform 1 0 1988 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1713453518
transform 1 0 2060 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1713453518
transform 1 0 1948 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1713453518
transform 1 0 1916 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1713453518
transform 1 0 1940 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1713453518
transform 1 0 1684 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1713453518
transform 1 0 1636 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1713453518
transform 1 0 1636 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1713453518
transform 1 0 1332 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1713453518
transform 1 0 3252 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1713453518
transform 1 0 3204 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1713453518
transform 1 0 3204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1713453518
transform 1 0 3164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1713453518
transform 1 0 2772 0 1 3055
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1713453518
transform 1 0 2580 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1713453518
transform 1 0 2532 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1713453518
transform 1 0 2476 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1713453518
transform 1 0 1748 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1713453518
transform 1 0 1748 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1713453518
transform 1 0 1708 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1713453518
transform 1 0 1692 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1713453518
transform 1 0 1564 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1713453518
transform 1 0 1404 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1713453518
transform 1 0 2348 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1713453518
transform 1 0 2236 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1713453518
transform 1 0 1724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1713453518
transform 1 0 1684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1713453518
transform 1 0 1396 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1713453518
transform 1 0 2692 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1713453518
transform 1 0 2668 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1713453518
transform 1 0 2716 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1713453518
transform 1 0 2700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1713453518
transform 1 0 2932 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1713453518
transform 1 0 2724 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1713453518
transform 1 0 2956 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1713453518
transform 1 0 2932 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1713453518
transform 1 0 3076 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1713453518
transform 1 0 2948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1713453518
transform 1 0 2660 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1713453518
transform 1 0 1580 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1713453518
transform 1 0 3260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1713453518
transform 1 0 3204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1713453518
transform 1 0 3012 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1713453518
transform 1 0 3012 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1713453518
transform 1 0 2972 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1713453518
transform 1 0 2956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1713453518
transform 1 0 2900 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1713453518
transform 1 0 2812 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1713453518
transform 1 0 2580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1713453518
transform 1 0 2356 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1713453518
transform 1 0 1748 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1713453518
transform 1 0 2988 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1713453518
transform 1 0 2964 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1713453518
transform 1 0 2612 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1713453518
transform 1 0 2588 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1713453518
transform 1 0 1692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1713453518
transform 1 0 2716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1713453518
transform 1 0 2628 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1713453518
transform 1 0 2308 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1713453518
transform 1 0 1812 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1713453518
transform 1 0 2652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1713453518
transform 1 0 2572 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1713453518
transform 1 0 2276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1713453518
transform 1 0 1884 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1713453518
transform 1 0 2604 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1713453518
transform 1 0 2604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1713453518
transform 1 0 2692 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1713453518
transform 1 0 2668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1713453518
transform 1 0 2676 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1713453518
transform 1 0 2572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1713453518
transform 1 0 2276 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1713453518
transform 1 0 2204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1713453518
transform 1 0 2708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1713453518
transform 1 0 2700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1713453518
transform 1 0 2636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1713453518
transform 1 0 2596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1713453518
transform 1 0 2612 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1713453518
transform 1 0 2572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1713453518
transform 1 0 2724 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1713453518
transform 1 0 2724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1713453518
transform 1 0 2884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1713453518
transform 1 0 2788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1713453518
transform 1 0 3396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1713453518
transform 1 0 3380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1713453518
transform 1 0 3236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1713453518
transform 1 0 3204 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1713453518
transform 1 0 2860 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1713453518
transform 1 0 2844 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1713453518
transform 1 0 2780 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1713453518
transform 1 0 2676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1713453518
transform 1 0 2580 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1713453518
transform 1 0 2564 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1713453518
transform 1 0 2548 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1713453518
transform 1 0 1908 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1713453518
transform 1 0 2972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1713453518
transform 1 0 2860 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1713453518
transform 1 0 2716 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1713453518
transform 1 0 2684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1713453518
transform 1 0 2972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1713453518
transform 1 0 2884 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1713453518
transform 1 0 2804 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1713453518
transform 1 0 2764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1713453518
transform 1 0 2788 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1713453518
transform 1 0 2780 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1713453518
transform 1 0 2820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1713453518
transform 1 0 2788 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1713453518
transform 1 0 2428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1713453518
transform 1 0 1836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1713453518
transform 1 0 2300 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1713453518
transform 1 0 2300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1713453518
transform 1 0 2284 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1713453518
transform 1 0 2284 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1713453518
transform 1 0 2364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1713453518
transform 1 0 2276 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1713453518
transform 1 0 2532 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1713453518
transform 1 0 2388 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1713453518
transform 1 0 2468 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1713453518
transform 1 0 2436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1713453518
transform 1 0 2668 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1713453518
transform 1 0 2388 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1713453518
transform 1 0 2524 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1713453518
transform 1 0 2412 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1713453518
transform 1 0 2428 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1713453518
transform 1 0 2428 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1713453518
transform 1 0 2388 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1713453518
transform 1 0 2188 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1713453518
transform 1 0 2164 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1713453518
transform 1 0 2116 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1713453518
transform 1 0 2228 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1713453518
transform 1 0 2124 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1713453518
transform 1 0 2172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1713453518
transform 1 0 2164 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1713453518
transform 1 0 2052 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1713453518
transform 1 0 2940 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1713453518
transform 1 0 2908 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1713453518
transform 1 0 2908 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1713453518
transform 1 0 2892 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1713453518
transform 1 0 2188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1713453518
transform 1 0 2148 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1713453518
transform 1 0 2036 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1713453518
transform 1 0 1820 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1713453518
transform 1 0 2644 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1713453518
transform 1 0 2484 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1713453518
transform 1 0 2252 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1713453518
transform 1 0 3244 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1713453518
transform 1 0 3228 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1713453518
transform 1 0 3036 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1713453518
transform 1 0 2812 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1713453518
transform 1 0 2236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1713453518
transform 1 0 1996 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1713453518
transform 1 0 1988 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1713453518
transform 1 0 3044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1713453518
transform 1 0 3012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1713453518
transform 1 0 2508 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1713453518
transform 1 0 2028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1713453518
transform 1 0 2012 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1713453518
transform 1 0 1924 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1713453518
transform 1 0 1868 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1713453518
transform 1 0 1852 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1713453518
transform 1 0 1836 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1713453518
transform 1 0 1924 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1713453518
transform 1 0 1788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1713453518
transform 1 0 1596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1713453518
transform 1 0 3252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1713453518
transform 1 0 3236 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1713453518
transform 1 0 3180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1713453518
transform 1 0 3092 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1713453518
transform 1 0 2556 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1713453518
transform 1 0 2500 0 1 2785
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1713453518
transform 1 0 2308 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1713453518
transform 1 0 1924 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1713453518
transform 1 0 2548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1713453518
transform 1 0 2508 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1713453518
transform 1 0 2508 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1713453518
transform 1 0 3028 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1713453518
transform 1 0 3020 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1713453518
transform 1 0 2972 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1713453518
transform 1 0 2540 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1713453518
transform 1 0 2404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1713453518
transform 1 0 2652 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1713453518
transform 1 0 2652 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1713453518
transform 1 0 2604 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1713453518
transform 1 0 2564 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1713453518
transform 1 0 3276 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1713453518
transform 1 0 3276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1713453518
transform 1 0 3260 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1713453518
transform 1 0 3236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1713453518
transform 1 0 2884 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1713453518
transform 1 0 2604 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1713453518
transform 1 0 2372 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1713453518
transform 1 0 2340 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1713453518
transform 1 0 2740 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1713453518
transform 1 0 2660 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1713453518
transform 1 0 3316 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1713453518
transform 1 0 3284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1713453518
transform 1 0 3236 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1713453518
transform 1 0 2828 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1713453518
transform 1 0 2684 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1713453518
transform 1 0 2356 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1713453518
transform 1 0 2028 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1713453518
transform 1 0 2756 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1713453518
transform 1 0 2732 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1713453518
transform 1 0 2556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1713453518
transform 1 0 2508 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1713453518
transform 1 0 2532 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1713453518
transform 1 0 2532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1713453518
transform 1 0 2516 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1713453518
transform 1 0 2516 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1713453518
transform 1 0 2532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1713453518
transform 1 0 2524 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1713453518
transform 1 0 3260 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1713453518
transform 1 0 3212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1713453518
transform 1 0 3204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1713453518
transform 1 0 3132 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1713453518
transform 1 0 2516 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1713453518
transform 1 0 2508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1713453518
transform 1 0 1924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1713453518
transform 1 0 1884 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1713453518
transform 1 0 1876 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1713453518
transform 1 0 2500 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1713453518
transform 1 0 2500 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1713453518
transform 1 0 2540 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1713453518
transform 1 0 2420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1713453518
transform 1 0 2364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1713453518
transform 1 0 2308 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1713453518
transform 1 0 2452 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1713453518
transform 1 0 2316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1713453518
transform 1 0 2860 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1713453518
transform 1 0 2788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1713453518
transform 1 0 2788 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1713453518
transform 1 0 2652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1713453518
transform 1 0 2484 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1713453518
transform 1 0 2436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1713453518
transform 1 0 2564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1713453518
transform 1 0 2564 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1713453518
transform 1 0 2532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1713453518
transform 1 0 2524 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1713453518
transform 1 0 2620 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1713453518
transform 1 0 2548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1713453518
transform 1 0 2548 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1713453518
transform 1 0 2332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1713453518
transform 1 0 2156 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1713453518
transform 1 0 2684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1713453518
transform 1 0 2596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1713453518
transform 1 0 2588 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1713453518
transform 1 0 2884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1713453518
transform 1 0 2868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1713453518
transform 1 0 2692 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1713453518
transform 1 0 2572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1713453518
transform 1 0 2540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1713453518
transform 1 0 2492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1713453518
transform 1 0 2116 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1713453518
transform 1 0 2100 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1713453518
transform 1 0 2100 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1713453518
transform 1 0 2676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1713453518
transform 1 0 2532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1713453518
transform 1 0 2892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1713453518
transform 1 0 2756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1713453518
transform 1 0 2676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1713453518
transform 1 0 2628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1713453518
transform 1 0 2620 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1713453518
transform 1 0 1804 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1713453518
transform 1 0 2564 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1713453518
transform 1 0 2420 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1713453518
transform 1 0 2388 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1713453518
transform 1 0 2308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1713453518
transform 1 0 2228 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1713453518
transform 1 0 2244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1713453518
transform 1 0 2236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1713453518
transform 1 0 2196 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1713453518
transform 1 0 2188 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1713453518
transform 1 0 2084 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1713453518
transform 1 0 2292 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1713453518
transform 1 0 2252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1713453518
transform 1 0 2460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1713453518
transform 1 0 2444 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1713453518
transform 1 0 2428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1713453518
transform 1 0 2204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1713453518
transform 1 0 2100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1713453518
transform 1 0 2100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1713453518
transform 1 0 2444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1713453518
transform 1 0 2332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1713453518
transform 1 0 2244 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1713453518
transform 1 0 2516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1713453518
transform 1 0 2412 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1713453518
transform 1 0 2388 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1713453518
transform 1 0 2276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1713453518
transform 1 0 1916 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1713453518
transform 1 0 1900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1713453518
transform 1 0 2332 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1713453518
transform 1 0 2260 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1713453518
transform 1 0 2260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1713453518
transform 1 0 2340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1713453518
transform 1 0 2300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1713453518
transform 1 0 2316 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1713453518
transform 1 0 2292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1713453518
transform 1 0 2548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1713453518
transform 1 0 2500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1713453518
transform 1 0 2444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1713453518
transform 1 0 2252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1713453518
transform 1 0 2236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1713453518
transform 1 0 2372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1713453518
transform 1 0 2300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1713453518
transform 1 0 2284 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1713453518
transform 1 0 2564 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1713453518
transform 1 0 2452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1713453518
transform 1 0 2404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1713453518
transform 1 0 2308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1713453518
transform 1 0 2212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1713453518
transform 1 0 2372 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1713453518
transform 1 0 2348 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1713453518
transform 1 0 2324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1713453518
transform 1 0 2556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1713453518
transform 1 0 2524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1713453518
transform 1 0 2444 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1713453518
transform 1 0 2324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1713453518
transform 1 0 2268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1713453518
transform 1 0 2316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1713453518
transform 1 0 2316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1713453518
transform 1 0 2276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1713453518
transform 1 0 2588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1713453518
transform 1 0 2484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1713453518
transform 1 0 2356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1713453518
transform 1 0 2140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1713453518
transform 1 0 1932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1713453518
transform 1 0 2388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1713453518
transform 1 0 2388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1713453518
transform 1 0 2380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1713453518
transform 1 0 2348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1713453518
transform 1 0 2404 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1713453518
transform 1 0 2356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1713453518
transform 1 0 2428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1713453518
transform 1 0 2404 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1713453518
transform 1 0 2948 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1713453518
transform 1 0 2916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1713453518
transform 1 0 2796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1713453518
transform 1 0 2524 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1713453518
transform 1 0 2380 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1713453518
transform 1 0 2052 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1713453518
transform 1 0 2036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1713453518
transform 1 0 2444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1713453518
transform 1 0 2404 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1713453518
transform 1 0 2404 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1713453518
transform 1 0 2572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1713453518
transform 1 0 2468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1713453518
transform 1 0 2452 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1713453518
transform 1 0 2428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1713453518
transform 1 0 2084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1713453518
transform 1 0 2076 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1713453518
transform 1 0 2540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1713453518
transform 1 0 2508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1713453518
transform 1 0 2484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1713453518
transform 1 0 2260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1713453518
transform 1 0 2244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1713453518
transform 1 0 1812 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1713453518
transform 1 0 1780 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1713453518
transform 1 0 1740 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1713453518
transform 1 0 1732 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1713453518
transform 1 0 1612 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1713453518
transform 1 0 1788 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1713453518
transform 1 0 1652 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1713453518
transform 1 0 1612 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1713453518
transform 1 0 2340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1713453518
transform 1 0 2244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1713453518
transform 1 0 2228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1713453518
transform 1 0 2188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1713453518
transform 1 0 2020 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1713453518
transform 1 0 2340 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1713453518
transform 1 0 2284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1713453518
transform 1 0 2252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1713453518
transform 1 0 2900 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1713453518
transform 1 0 2860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1713453518
transform 1 0 2836 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1713453518
transform 1 0 2476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1713453518
transform 1 0 2276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1713453518
transform 1 0 2060 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1713453518
transform 1 0 2012 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1713453518
transform 1 0 2388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1713453518
transform 1 0 2356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1713453518
transform 1 0 2012 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1713453518
transform 1 0 1972 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1713453518
transform 1 0 1972 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1713453518
transform 1 0 1972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1713453518
transform 1 0 1948 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1713453518
transform 1 0 1940 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1713453518
transform 1 0 2036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1713453518
transform 1 0 1948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1713453518
transform 1 0 1988 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1713453518
transform 1 0 1948 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1713453518
transform 1 0 2252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1713453518
transform 1 0 2020 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1713453518
transform 1 0 2068 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1713453518
transform 1 0 2044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1713453518
transform 1 0 2020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1713453518
transform 1 0 2020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1713453518
transform 1 0 1980 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1713453518
transform 1 0 2044 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1713453518
transform 1 0 2028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1713453518
transform 1 0 2012 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1713453518
transform 1 0 2012 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1713453518
transform 1 0 1948 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1713453518
transform 1 0 1852 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1713453518
transform 1 0 2052 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1713453518
transform 1 0 1852 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1713453518
transform 1 0 1484 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1713453518
transform 1 0 2348 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1713453518
transform 1 0 2244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1713453518
transform 1 0 2340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1713453518
transform 1 0 2284 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1713453518
transform 1 0 2260 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1713453518
transform 1 0 1924 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1713453518
transform 1 0 1716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1713453518
transform 1 0 2372 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1713453518
transform 1 0 2372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1713453518
transform 1 0 2116 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1713453518
transform 1 0 2308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1713453518
transform 1 0 2308 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1713453518
transform 1 0 2372 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1713453518
transform 1 0 2372 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1713453518
transform 1 0 2156 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1713453518
transform 1 0 2132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1713453518
transform 1 0 2092 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1713453518
transform 1 0 2052 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1713453518
transform 1 0 2052 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1713453518
transform 1 0 2164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1713453518
transform 1 0 2012 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1713453518
transform 1 0 1884 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1713453518
transform 1 0 2364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1713453518
transform 1 0 2156 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1713453518
transform 1 0 2396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1713453518
transform 1 0 2348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1713453518
transform 1 0 2348 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1713453518
transform 1 0 2468 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1713453518
transform 1 0 2372 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1713453518
transform 1 0 2132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1713453518
transform 1 0 1916 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1713453518
transform 1 0 1916 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1713453518
transform 1 0 1852 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1713453518
transform 1 0 1812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1713453518
transform 1 0 1964 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1713453518
transform 1 0 1964 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1713453518
transform 1 0 1932 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1713453518
transform 1 0 1932 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1713453518
transform 1 0 2004 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1713453518
transform 1 0 1972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1713453518
transform 1 0 1852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1713453518
transform 1 0 1996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1713453518
transform 1 0 1996 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1713453518
transform 1 0 1972 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1713453518
transform 1 0 1964 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1713453518
transform 1 0 2028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1713453518
transform 1 0 1988 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1713453518
transform 1 0 1996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1713453518
transform 1 0 1948 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1713453518
transform 1 0 2076 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1713453518
transform 1 0 2012 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1713453518
transform 1 0 2252 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1713453518
transform 1 0 2100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1713453518
transform 1 0 2060 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1713453518
transform 1 0 2100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1713453518
transform 1 0 1964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1713453518
transform 1 0 2052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1713453518
transform 1 0 1876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1713453518
transform 1 0 1900 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1713453518
transform 1 0 1732 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1713453518
transform 1 0 1652 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1713453518
transform 1 0 1652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1713453518
transform 1 0 1564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1713453518
transform 1 0 1564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1713453518
transform 1 0 1756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1713453518
transform 1 0 1756 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1713453518
transform 1 0 1724 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1713453518
transform 1 0 1724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1713453518
transform 1 0 1748 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1713453518
transform 1 0 1668 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1713453518
transform 1 0 1668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1713453518
transform 1 0 1740 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1713453518
transform 1 0 1740 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1713453518
transform 1 0 1660 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1713453518
transform 1 0 2228 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1713453518
transform 1 0 1988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1713453518
transform 1 0 1820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1713453518
transform 1 0 2084 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1713453518
transform 1 0 2076 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1713453518
transform 1 0 1988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1713453518
transform 1 0 2044 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1713453518
transform 1 0 2020 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1713453518
transform 1 0 2068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1713453518
transform 1 0 2052 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1713453518
transform 1 0 2100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1713453518
transform 1 0 2100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1713453518
transform 1 0 2060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1713453518
transform 1 0 2100 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1713453518
transform 1 0 2076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1713453518
transform 1 0 2052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1713453518
transform 1 0 2044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1713453518
transform 1 0 2028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1713453518
transform 1 0 2124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1713453518
transform 1 0 1924 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1713453518
transform 1 0 1948 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1713453518
transform 1 0 1884 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1713453518
transform 1 0 1892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1713453518
transform 1 0 1876 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1713453518
transform 1 0 1860 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1713453518
transform 1 0 1852 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1713453518
transform 1 0 1852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1713453518
transform 1 0 1876 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1713453518
transform 1 0 1820 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1713453518
transform 1 0 1796 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1713453518
transform 1 0 1892 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1713453518
transform 1 0 1876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1713453518
transform 1 0 1876 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1713453518
transform 1 0 2124 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1713453518
transform 1 0 2076 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1713453518
transform 1 0 1988 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1713453518
transform 1 0 2196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1713453518
transform 1 0 2132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1713453518
transform 1 0 2100 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1713453518
transform 1 0 1940 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1713453518
transform 1 0 1892 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1713453518
transform 1 0 2148 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1713453518
transform 1 0 1900 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1713453518
transform 1 0 2228 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1713453518
transform 1 0 2124 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1713453518
transform 1 0 2156 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1713453518
transform 1 0 2124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1713453518
transform 1 0 2092 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1713453518
transform 1 0 2092 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1713453518
transform 1 0 2412 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1713453518
transform 1 0 2060 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1713453518
transform 1 0 2076 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1713453518
transform 1 0 1556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1713453518
transform 1 0 1540 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1713453518
transform 1 0 1500 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1713453518
transform 1 0 1252 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1713453518
transform 1 0 1252 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1713453518
transform 1 0 1548 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1713453518
transform 1 0 1444 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1713453518
transform 1 0 2396 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1713453518
transform 1 0 2316 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1713453518
transform 1 0 2940 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1713453518
transform 1 0 2444 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1713453518
transform 1 0 2932 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1713453518
transform 1 0 2860 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1713453518
transform 1 0 2796 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1713453518
transform 1 0 2324 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1713453518
transform 1 0 1228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1713453518
transform 1 0 2948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1713453518
transform 1 0 2708 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1713453518
transform 1 0 2644 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1713453518
transform 1 0 2396 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1713453518
transform 1 0 1196 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1713453518
transform 1 0 2220 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1713453518
transform 1 0 2108 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1713453518
transform 1 0 1308 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1713453518
transform 1 0 1260 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1713453518
transform 1 0 2324 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1713453518
transform 1 0 1932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1713453518
transform 1 0 1540 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1713453518
transform 1 0 1356 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1713453518
transform 1 0 1356 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1713453518
transform 1 0 2316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1713453518
transform 1 0 2132 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1713453518
transform 1 0 2220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1713453518
transform 1 0 2140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1713453518
transform 1 0 2172 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1713453518
transform 1 0 2012 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1713453518
transform 1 0 1820 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1713453518
transform 1 0 1788 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1713453518
transform 1 0 1660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1713453518
transform 1 0 1148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1713453518
transform 1 0 2276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1713453518
transform 1 0 2100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1713453518
transform 1 0 1740 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1713453518
transform 1 0 1660 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1713453518
transform 1 0 1612 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1713453518
transform 1 0 2252 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1713453518
transform 1 0 2220 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1713453518
transform 1 0 2156 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1713453518
transform 1 0 1460 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1713453518
transform 1 0 2788 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1713453518
transform 1 0 2660 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1713453518
transform 1 0 2332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1713453518
transform 1 0 1964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1713453518
transform 1 0 1692 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1713453518
transform 1 0 2188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1713453518
transform 1 0 2148 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1713453518
transform 1 0 1532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1713453518
transform 1 0 1492 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1713453518
transform 1 0 1492 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1713453518
transform 1 0 1460 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1713453518
transform 1 0 1452 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1713453518
transform 1 0 2172 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1713453518
transform 1 0 2156 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1713453518
transform 1 0 2100 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1713453518
transform 1 0 2004 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1713453518
transform 1 0 1604 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1713453518
transform 1 0 1588 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1713453518
transform 1 0 1548 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1713453518
transform 1 0 1292 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1713453518
transform 1 0 2180 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1713453518
transform 1 0 1932 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1713453518
transform 1 0 1524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1713453518
transform 1 0 1404 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1713453518
transform 1 0 1132 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1713453518
transform 1 0 1916 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1713453518
transform 1 0 1908 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1713453518
transform 1 0 1908 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1713453518
transform 1 0 1908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1713453518
transform 1 0 2084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1713453518
transform 1 0 1980 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1713453518
transform 1 0 1940 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1713453518
transform 1 0 1924 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1713453518
transform 1 0 2100 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1713453518
transform 1 0 2076 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1713453518
transform 1 0 2100 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1713453518
transform 1 0 2092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1713453518
transform 1 0 2092 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1713453518
transform 1 0 2036 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1713453518
transform 1 0 1196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1713453518
transform 1 0 3404 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1713453518
transform 1 0 3388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1713453518
transform 1 0 3364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1713453518
transform 1 0 3332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1713453518
transform 1 0 3116 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1713453518
transform 1 0 2908 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1713453518
transform 1 0 2892 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1713453518
transform 1 0 2572 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1713453518
transform 1 0 2556 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1713453518
transform 1 0 2532 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1713453518
transform 1 0 2436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1713453518
transform 1 0 2028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1713453518
transform 1 0 1908 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1713453518
transform 1 0 2164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1713453518
transform 1 0 2140 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1713453518
transform 1 0 2116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1713453518
transform 1 0 2116 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1713453518
transform 1 0 2052 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1713453518
transform 1 0 1716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1713453518
transform 1 0 1604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1713453518
transform 1 0 1260 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1713453518
transform 1 0 2204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1713453518
transform 1 0 2204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1713453518
transform 1 0 2156 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1713453518
transform 1 0 1788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1713453518
transform 1 0 1724 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1713453518
transform 1 0 1428 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1713453518
transform 1 0 1340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1713453518
transform 1 0 2196 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1713453518
transform 1 0 2124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1713453518
transform 1 0 2180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1713453518
transform 1 0 2156 0 1 1495
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1713453518
transform 1 0 2236 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1713453518
transform 1 0 2132 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1713453518
transform 1 0 1924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1713453518
transform 1 0 1524 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1713453518
transform 1 0 2228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1713453518
transform 1 0 2020 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1713453518
transform 1 0 1676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1713453518
transform 1 0 1564 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1713453518
transform 1 0 1516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1713453518
transform 1 0 2132 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1713453518
transform 1 0 1708 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1713453518
transform 1 0 1684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1713453518
transform 1 0 1452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1713453518
transform 1 0 2204 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1713453518
transform 1 0 2204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1713453518
transform 1 0 1708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1713453518
transform 1 0 1708 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1713453518
transform 1 0 1500 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1713453518
transform 1 0 1916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1713453518
transform 1 0 1908 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1713453518
transform 1 0 2156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1713453518
transform 1 0 1884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1713453518
transform 1 0 1740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1713453518
transform 1 0 1724 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1713453518
transform 1 0 1340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1713453518
transform 1 0 2140 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1713453518
transform 1 0 1932 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1713453518
transform 1 0 1748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1713453518
transform 1 0 1684 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1713453518
transform 1 0 1300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1713453518
transform 1 0 1868 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1713453518
transform 1 0 1764 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1713453518
transform 1 0 1532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1713453518
transform 1 0 1340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1713453518
transform 1 0 1876 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1713453518
transform 1 0 1860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1713453518
transform 1 0 1956 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1713453518
transform 1 0 1892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1713453518
transform 1 0 2604 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1713453518
transform 1 0 2532 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1713453518
transform 1 0 2012 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1713453518
transform 1 0 1924 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1713453518
transform 1 0 1580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1713453518
transform 1 0 2540 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1713453518
transform 1 0 2508 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1713453518
transform 1 0 2156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1713453518
transform 1 0 2116 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1713453518
transform 1 0 1972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1713453518
transform 1 0 1628 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1713453518
transform 1 0 1836 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1713453518
transform 1 0 1820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1713453518
transform 1 0 1676 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1713453518
transform 1 0 1652 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1713453518
transform 1 0 1604 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1713453518
transform 1 0 1460 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1713453518
transform 1 0 1460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1713453518
transform 1 0 2092 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1713453518
transform 1 0 1892 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1713453518
transform 1 0 1740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1713453518
transform 1 0 1724 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1713453518
transform 1 0 1692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1713453518
transform 1 0 1428 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1713453518
transform 1 0 2932 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1713453518
transform 1 0 2836 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1713453518
transform 1 0 3092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1713453518
transform 1 0 2972 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1713453518
transform 1 0 3052 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1713453518
transform 1 0 2980 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1713453518
transform 1 0 3436 0 1 1755
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1713453518
transform 1 0 3100 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1713453518
transform 1 0 3444 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1713453518
transform 1 0 3372 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1713453518
transform 1 0 3412 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1713453518
transform 1 0 3396 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1713453518
transform 1 0 3428 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1713453518
transform 1 0 3428 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1713453518
transform 1 0 3404 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1713453518
transform 1 0 3068 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1713453518
transform 1 0 3420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1713453518
transform 1 0 3404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1713453518
transform 1 0 3364 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1713453518
transform 1 0 3244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1713453518
transform 1 0 3404 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1713453518
transform 1 0 3380 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1713453518
transform 1 0 3364 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1713453518
transform 1 0 3348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1713453518
transform 1 0 2852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1713453518
transform 1 0 2772 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1713453518
transform 1 0 2764 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1713453518
transform 1 0 2764 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1713453518
transform 1 0 2732 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1713453518
transform 1 0 2724 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1713453518
transform 1 0 2684 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1713453518
transform 1 0 2420 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1713453518
transform 1 0 2364 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1713453518
transform 1 0 2308 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1713453518
transform 1 0 1844 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1713453518
transform 1 0 3404 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1713453518
transform 1 0 3332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1713453518
transform 1 0 3284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1713453518
transform 1 0 3284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1713453518
transform 1 0 3244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1713453518
transform 1 0 3236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1713453518
transform 1 0 3340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1713453518
transform 1 0 3340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1713453518
transform 1 0 3324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1713453518
transform 1 0 3324 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1713453518
transform 1 0 3412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1713453518
transform 1 0 3356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1713453518
transform 1 0 3316 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1713453518
transform 1 0 3212 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1713453518
transform 1 0 3188 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1713453518
transform 1 0 3188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1713453518
transform 1 0 3164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1713453518
transform 1 0 2852 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1713453518
transform 1 0 2836 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1713453518
transform 1 0 2812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1713453518
transform 1 0 2812 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1713453518
transform 1 0 2796 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1713453518
transform 1 0 2580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1713453518
transform 1 0 2420 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1713453518
transform 1 0 2380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1713453518
transform 1 0 2268 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1713453518
transform 1 0 1796 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1713453518
transform 1 0 3204 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1713453518
transform 1 0 3164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1713453518
transform 1 0 3188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1713453518
transform 1 0 3156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1713453518
transform 1 0 3180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1713453518
transform 1 0 2892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1713453518
transform 1 0 2860 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1713453518
transform 1 0 2980 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1713453518
transform 1 0 2956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1713453518
transform 1 0 2956 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1713453518
transform 1 0 2972 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1713453518
transform 1 0 2868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1713453518
transform 1 0 3020 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1713453518
transform 1 0 3012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1713453518
transform 1 0 3012 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1713453518
transform 1 0 3012 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1713453518
transform 1 0 3052 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1713453518
transform 1 0 3052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1713453518
transform 1 0 3004 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1713453518
transform 1 0 2988 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1713453518
transform 1 0 2916 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1713453518
transform 1 0 2884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1713453518
transform 1 0 2940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1713453518
transform 1 0 2868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1713453518
transform 1 0 2868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1713453518
transform 1 0 2908 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1713453518
transform 1 0 2804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1713453518
transform 1 0 2804 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1713453518
transform 1 0 3164 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1713453518
transform 1 0 3164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1713453518
transform 1 0 3052 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1713453518
transform 1 0 2996 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1713453518
transform 1 0 2876 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1713453518
transform 1 0 3020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1713453518
transform 1 0 3020 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1713453518
transform 1 0 2988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1713453518
transform 1 0 2868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1713453518
transform 1 0 2860 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1713453518
transform 1 0 2876 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1713453518
transform 1 0 2780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1713453518
transform 1 0 2764 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1713453518
transform 1 0 3420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1713453518
transform 1 0 3196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1713453518
transform 1 0 3228 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1713453518
transform 1 0 3156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1713453518
transform 1 0 3140 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1713453518
transform 1 0 3140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1713453518
transform 1 0 3132 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1713453518
transform 1 0 3132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1713453518
transform 1 0 3092 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1713453518
transform 1 0 2812 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1713453518
transform 1 0 2756 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1713453518
transform 1 0 2692 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1713453518
transform 1 0 2692 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1713453518
transform 1 0 2500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1713453518
transform 1 0 1772 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1713453518
transform 1 0 3172 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1713453518
transform 1 0 3076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1713453518
transform 1 0 3068 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1713453518
transform 1 0 3068 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1713453518
transform 1 0 3084 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1713453518
transform 1 0 2956 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1713453518
transform 1 0 2908 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1713453518
transform 1 0 3028 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1713453518
transform 1 0 2988 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1713453518
transform 1 0 2980 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1713453518
transform 1 0 3396 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1713453518
transform 1 0 3316 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1713453518
transform 1 0 3340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1713453518
transform 1 0 3300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1713453518
transform 1 0 3340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1713453518
transform 1 0 3340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1713453518
transform 1 0 3404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1713453518
transform 1 0 3404 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1713453518
transform 1 0 3340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1713453518
transform 1 0 3316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1713453518
transform 1 0 3444 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1713453518
transform 1 0 3444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1713453518
transform 1 0 3420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1713453518
transform 1 0 3356 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1713453518
transform 1 0 3436 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1713453518
transform 1 0 3388 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1713453518
transform 1 0 2396 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1713453518
transform 1 0 2348 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1713453518
transform 1 0 2348 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1713453518
transform 1 0 3380 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1713453518
transform 1 0 3364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1713453518
transform 1 0 3348 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1713453518
transform 1 0 3364 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1713453518
transform 1 0 3292 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1713453518
transform 1 0 3212 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1713453518
transform 1 0 3420 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1713453518
transform 1 0 3372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1713453518
transform 1 0 3388 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1713453518
transform 1 0 3364 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1713453518
transform 1 0 3380 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1713453518
transform 1 0 3332 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1713453518
transform 1 0 3316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1713453518
transform 1 0 3404 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1713453518
transform 1 0 3316 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1713453518
transform 1 0 3316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1713453518
transform 1 0 2964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1713453518
transform 1 0 2556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1713453518
transform 1 0 2964 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1713453518
transform 1 0 2956 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1713453518
transform 1 0 2948 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1713453518
transform 1 0 2940 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1713453518
transform 1 0 2972 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1713453518
transform 1 0 2972 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1713453518
transform 1 0 2940 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1713453518
transform 1 0 2916 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1713453518
transform 1 0 2948 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1713453518
transform 1 0 2796 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1713453518
transform 1 0 2004 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1713453518
transform 1 0 3292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1713453518
transform 1 0 2956 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1713453518
transform 1 0 3244 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1713453518
transform 1 0 3236 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1713453518
transform 1 0 3276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1713453518
transform 1 0 3252 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1713453518
transform 1 0 3292 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1713453518
transform 1 0 3220 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1713453518
transform 1 0 3220 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1713453518
transform 1 0 3260 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1713453518
transform 1 0 3140 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1713453518
transform 1 0 3124 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1713453518
transform 1 0 2892 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1713453518
transform 1 0 2884 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1713453518
transform 1 0 2884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1713453518
transform 1 0 2868 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1713453518
transform 1 0 2852 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1713453518
transform 1 0 3028 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1713453518
transform 1 0 2924 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1713453518
transform 1 0 2908 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1713453518
transform 1 0 2908 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1713453518
transform 1 0 2764 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1713453518
transform 1 0 2900 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1713453518
transform 1 0 2884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1713453518
transform 1 0 3052 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1713453518
transform 1 0 2932 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1713453518
transform 1 0 3196 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1713453518
transform 1 0 3060 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1713453518
transform 1 0 3028 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1713453518
transform 1 0 3116 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1713453518
transform 1 0 3060 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1713453518
transform 1 0 3196 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1713453518
transform 1 0 3180 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1713453518
transform 1 0 3108 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1713453518
transform 1 0 3180 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1713453518
transform 1 0 3148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1713453518
transform 1 0 3164 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1713453518
transform 1 0 2868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1713453518
transform 1 0 2964 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1713453518
transform 1 0 2948 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1713453518
transform 1 0 2932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1713453518
transform 1 0 2836 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1713453518
transform 1 0 2772 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1713453518
transform 1 0 2748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1713453518
transform 1 0 2716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1713453518
transform 1 0 2684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1713453518
transform 1 0 2636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1713453518
transform 1 0 2548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1713453518
transform 1 0 2020 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1713453518
transform 1 0 2812 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1713453518
transform 1 0 2788 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1713453518
transform 1 0 2740 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1713453518
transform 1 0 2772 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1713453518
transform 1 0 2684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1713453518
transform 1 0 2604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1713453518
transform 1 0 2588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1713453518
transform 1 0 2212 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1713453518
transform 1 0 2532 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1713453518
transform 1 0 2532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1713453518
transform 1 0 2548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1713453518
transform 1 0 2532 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1713453518
transform 1 0 2524 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1713453518
transform 1 0 2508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1713453518
transform 1 0 3372 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1713453518
transform 1 0 3220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1713453518
transform 1 0 2492 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1713453518
transform 1 0 2692 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1713453518
transform 1 0 2556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1713453518
transform 1 0 3044 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1713453518
transform 1 0 2868 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1713453518
transform 1 0 2780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1713453518
transform 1 0 2580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1713453518
transform 1 0 2540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3699
timestamp 1713453518
transform 1 0 2556 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1713453518
transform 1 0 2556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1713453518
transform 1 0 2692 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3702
timestamp 1713453518
transform 1 0 2596 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1713453518
transform 1 0 2540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1713453518
transform 1 0 2732 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1713453518
transform 1 0 2652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1713453518
transform 1 0 2572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3707
timestamp 1713453518
transform 1 0 2644 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3708
timestamp 1713453518
transform 1 0 2564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1713453518
transform 1 0 3220 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1713453518
transform 1 0 3220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1713453518
transform 1 0 2604 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1713453518
transform 1 0 2948 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1713453518
transform 1 0 2916 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1713453518
transform 1 0 2940 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1713453518
transform 1 0 2940 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1713453518
transform 1 0 2916 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1713453518
transform 1 0 2852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1713453518
transform 1 0 3036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1713453518
transform 1 0 2852 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1713453518
transform 1 0 2836 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1713453518
transform 1 0 2844 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1713453518
transform 1 0 2780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1713453518
transform 1 0 2716 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1713453518
transform 1 0 2612 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1713453518
transform 1 0 2100 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1713453518
transform 1 0 3100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1713453518
transform 1 0 2972 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1713453518
transform 1 0 2892 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1713453518
transform 1 0 3196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1713453518
transform 1 0 3196 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1713453518
transform 1 0 2996 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1713453518
transform 1 0 2956 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1713453518
transform 1 0 2908 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1713453518
transform 1 0 2852 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1713453518
transform 1 0 2820 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1713453518
transform 1 0 2724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1713453518
transform 1 0 3036 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1713453518
transform 1 0 2964 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1713453518
transform 1 0 2956 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1713453518
transform 1 0 3148 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1713453518
transform 1 0 3100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1713453518
transform 1 0 3092 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1713453518
transform 1 0 3092 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1713453518
transform 1 0 3068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1713453518
transform 1 0 3068 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1713453518
transform 1 0 3428 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1713453518
transform 1 0 3052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1713453518
transform 1 0 3100 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1713453518
transform 1 0 2956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1713453518
transform 1 0 2748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1713453518
transform 1 0 3412 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1713453518
transform 1 0 3404 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3753
timestamp 1713453518
transform 1 0 3412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1713453518
transform 1 0 3388 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1713453518
transform 1 0 3452 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1713453518
transform 1 0 3420 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1713453518
transform 1 0 3420 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1713453518
transform 1 0 3420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1713453518
transform 1 0 3452 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1713453518
transform 1 0 3420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1713453518
transform 1 0 3412 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1713453518
transform 1 0 2924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1713453518
transform 1 0 3020 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1713453518
transform 1 0 2916 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1713453518
transform 1 0 2916 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3766
timestamp 1713453518
transform 1 0 2996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1713453518
transform 1 0 2932 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1713453518
transform 1 0 2892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1713453518
transform 1 0 3428 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1713453518
transform 1 0 3420 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1713453518
transform 1 0 3404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1713453518
transform 1 0 3428 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1713453518
transform 1 0 3380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1713453518
transform 1 0 3420 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1713453518
transform 1 0 3332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1713453518
transform 1 0 3324 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1713453518
transform 1 0 3420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1713453518
transform 1 0 3388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1713453518
transform 1 0 3388 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1713453518
transform 1 0 3364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1713453518
transform 1 0 3292 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1713453518
transform 1 0 3196 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1713453518
transform 1 0 3396 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1713453518
transform 1 0 3364 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3785
timestamp 1713453518
transform 1 0 3356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1713453518
transform 1 0 3380 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1713453518
transform 1 0 3380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1713453518
transform 1 0 3332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1713453518
transform 1 0 3300 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1713453518
transform 1 0 3404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1713453518
transform 1 0 3372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1713453518
transform 1 0 3340 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1713453518
transform 1 0 3396 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1713453518
transform 1 0 3316 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1713453518
transform 1 0 3292 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1713453518
transform 1 0 3260 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1713453518
transform 1 0 3236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1713453518
transform 1 0 3348 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1713453518
transform 1 0 3332 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1713453518
transform 1 0 3332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1713453518
transform 1 0 2188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1713453518
transform 1 0 2060 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1713453518
transform 1 0 2276 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1713453518
transform 1 0 2260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1713453518
transform 1 0 2188 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1713453518
transform 1 0 2188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1713453518
transform 1 0 2764 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3808
timestamp 1713453518
transform 1 0 2764 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1713453518
transform 1 0 2100 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1713453518
transform 1 0 1340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1713453518
transform 1 0 3164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1713453518
transform 1 0 3044 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1713453518
transform 1 0 3068 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1713453518
transform 1 0 3068 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1713453518
transform 1 0 3332 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1713453518
transform 1 0 3060 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1713453518
transform 1 0 3436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1713453518
transform 1 0 3364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1713453518
transform 1 0 3436 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1713453518
transform 1 0 3380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1713453518
transform 1 0 3372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1713453518
transform 1 0 3364 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1713453518
transform 1 0 3300 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1713453518
transform 1 0 3388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1713453518
transform 1 0 3356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3826
timestamp 1713453518
transform 1 0 3324 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1713453518
transform 1 0 3420 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1713453518
transform 1 0 3420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1713453518
transform 1 0 3324 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1713453518
transform 1 0 3300 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1713453518
transform 1 0 2884 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1713453518
transform 1 0 2956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1713453518
transform 1 0 2876 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1713453518
transform 1 0 2876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1713453518
transform 1 0 2972 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1713453518
transform 1 0 2892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1713453518
transform 1 0 2836 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1713453518
transform 1 0 3268 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1713453518
transform 1 0 3236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1713453518
transform 1 0 3236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1713453518
transform 1 0 3044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1713453518
transform 1 0 2980 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1713453518
transform 1 0 3052 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1713453518
transform 1 0 2828 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1713453518
transform 1 0 2828 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1713453518
transform 1 0 2812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1713453518
transform 1 0 2788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1713453518
transform 1 0 2844 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1713453518
transform 1 0 2828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1713453518
transform 1 0 2804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1713453518
transform 1 0 2940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1713453518
transform 1 0 2940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1713453518
transform 1 0 2996 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1713453518
transform 1 0 2972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1713453518
transform 1 0 2908 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1713453518
transform 1 0 3276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1713453518
transform 1 0 3276 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1713453518
transform 1 0 3164 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1713453518
transform 1 0 3148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1713453518
transform 1 0 3068 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1713453518
transform 1 0 2988 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1713453518
transform 1 0 3084 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1713453518
transform 1 0 2932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1713453518
transform 1 0 2932 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1713453518
transform 1 0 3012 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1713453518
transform 1 0 2964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1713453518
transform 1 0 2860 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1713453518
transform 1 0 2756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1713453518
transform 1 0 2564 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1713453518
transform 1 0 2788 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1713453518
transform 1 0 2764 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1713453518
transform 1 0 2740 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1713453518
transform 1 0 2724 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1713453518
transform 1 0 2820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1713453518
transform 1 0 2764 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1713453518
transform 1 0 2868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1713453518
transform 1 0 2772 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1713453518
transform 1 0 2748 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1713453518
transform 1 0 2748 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1713453518
transform 1 0 2708 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1713453518
transform 1 0 2676 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1713453518
transform 1 0 2724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1713453518
transform 1 0 2708 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1713453518
transform 1 0 2692 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1713453518
transform 1 0 2548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1713453518
transform 1 0 2604 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1713453518
transform 1 0 2468 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1713453518
transform 1 0 2452 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1713453518
transform 1 0 2564 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1713453518
transform 1 0 2452 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1713453518
transform 1 0 2436 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1713453518
transform 1 0 2716 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1713453518
transform 1 0 2676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1713453518
transform 1 0 2612 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1713453518
transform 1 0 2604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1713453518
transform 1 0 2580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1713453518
transform 1 0 2660 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1713453518
transform 1 0 2620 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1713453518
transform 1 0 2788 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1713453518
transform 1 0 2604 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1713453518
transform 1 0 2452 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1713453518
transform 1 0 2644 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1713453518
transform 1 0 2644 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_3904
timestamp 1713453518
transform 1 0 2596 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1713453518
transform 1 0 2300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1713453518
transform 1 0 2564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1713453518
transform 1 0 2428 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1713453518
transform 1 0 2308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1713453518
transform 1 0 2612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3910
timestamp 1713453518
transform 1 0 2492 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1713453518
transform 1 0 2356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1713453518
transform 1 0 2900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1713453518
transform 1 0 2796 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1713453518
transform 1 0 2612 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1713453518
transform 1 0 2868 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3916
timestamp 1713453518
transform 1 0 2860 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1713453518
transform 1 0 2980 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1713453518
transform 1 0 2820 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1713453518
transform 1 0 2740 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1713453518
transform 1 0 2932 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1713453518
transform 1 0 2876 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1713453518
transform 1 0 2708 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3923
timestamp 1713453518
transform 1 0 2852 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1713453518
transform 1 0 2804 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3925
timestamp 1713453518
transform 1 0 2924 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3926
timestamp 1713453518
transform 1 0 2868 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1713453518
transform 1 0 2836 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3928
timestamp 1713453518
transform 1 0 2860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1713453518
transform 1 0 2852 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1713453518
transform 1 0 2836 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1713453518
transform 1 0 2772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1713453518
transform 1 0 2004 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1713453518
transform 1 0 1996 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3934
timestamp 1713453518
transform 1 0 2012 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3935
timestamp 1713453518
transform 1 0 1892 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1713453518
transform 1 0 1884 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3937
timestamp 1713453518
transform 1 0 1884 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1713453518
transform 1 0 1804 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3939
timestamp 1713453518
transform 1 0 1772 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1713453518
transform 1 0 1924 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1713453518
transform 1 0 1900 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3942
timestamp 1713453518
transform 1 0 1836 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3943
timestamp 1713453518
transform 1 0 1804 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1713453518
transform 1 0 2180 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1713453518
transform 1 0 1988 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3946
timestamp 1713453518
transform 1 0 1988 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3947
timestamp 1713453518
transform 1 0 2508 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1713453518
transform 1 0 2420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1713453518
transform 1 0 2548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1713453518
transform 1 0 2468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1713453518
transform 1 0 2588 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3952
timestamp 1713453518
transform 1 0 2556 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1713453518
transform 1 0 2676 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1713453518
transform 1 0 2636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1713453518
transform 1 0 2684 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1713453518
transform 1 0 2644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1713453518
transform 1 0 2596 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1713453518
transform 1 0 2596 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1713453518
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1713453518
transform 1 0 2508 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3961
timestamp 1713453518
transform 1 0 2668 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1713453518
transform 1 0 2660 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1713453518
transform 1 0 2516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3964
timestamp 1713453518
transform 1 0 2900 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3965
timestamp 1713453518
transform 1 0 2708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1713453518
transform 1 0 2564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3967
timestamp 1713453518
transform 1 0 2572 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1713453518
transform 1 0 2516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1713453518
transform 1 0 2468 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1713453518
transform 1 0 2372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1713453518
transform 1 0 2532 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1713453518
transform 1 0 2516 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1713453518
transform 1 0 2428 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3974
timestamp 1713453518
transform 1 0 2596 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3975
timestamp 1713453518
transform 1 0 2540 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1713453518
transform 1 0 2516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1713453518
transform 1 0 2492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1713453518
transform 1 0 2436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1713453518
transform 1 0 2428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3980
timestamp 1713453518
transform 1 0 2452 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1713453518
transform 1 0 2412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3982
timestamp 1713453518
transform 1 0 2452 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1713453518
transform 1 0 2404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1713453518
transform 1 0 2340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1713453518
transform 1 0 2428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1713453518
transform 1 0 2380 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3987
timestamp 1713453518
transform 1 0 2284 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1713453518
transform 1 0 2484 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1713453518
transform 1 0 2380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1713453518
transform 1 0 2332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1713453518
transform 1 0 2436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1713453518
transform 1 0 2436 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1713453518
transform 1 0 2356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1713453518
transform 1 0 2420 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3995
timestamp 1713453518
transform 1 0 2380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1713453518
transform 1 0 2324 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1713453518
transform 1 0 2412 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1713453518
transform 1 0 2412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1713453518
transform 1 0 2524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1713453518
transform 1 0 2508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1713453518
transform 1 0 2500 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1713453518
transform 1 0 2340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1713453518
transform 1 0 2308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1713453518
transform 1 0 2596 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1713453518
transform 1 0 2420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4006
timestamp 1713453518
transform 1 0 2316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1713453518
transform 1 0 1532 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1713453518
transform 1 0 932 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1713453518
transform 1 0 1540 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4010
timestamp 1713453518
transform 1 0 1508 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1713453518
transform 1 0 1596 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4012
timestamp 1713453518
transform 1 0 1516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1713453518
transform 1 0 1628 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1713453518
transform 1 0 1628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1713453518
transform 1 0 3220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1713453518
transform 1 0 3212 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1713453518
transform 1 0 3196 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1713453518
transform 1 0 3172 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1713453518
transform 1 0 3172 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1713453518
transform 1 0 2964 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1713453518
transform 1 0 1828 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4022
timestamp 1713453518
transform 1 0 1708 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1713453518
transform 1 0 1708 0 1 2895
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1713453518
transform 1 0 1660 0 1 2895
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1713453518
transform 1 0 1660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1713453518
transform 1 0 1684 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1713453518
transform 1 0 1068 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4028
timestamp 1713453518
transform 1 0 1796 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4029
timestamp 1713453518
transform 1 0 1516 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1713453518
transform 1 0 1628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1713453518
transform 1 0 1508 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1713453518
transform 1 0 2132 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1713453518
transform 1 0 2108 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1713453518
transform 1 0 2092 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1713453518
transform 1 0 2068 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1713453518
transform 1 0 2012 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4037
timestamp 1713453518
transform 1 0 1932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1713453518
transform 1 0 1852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4039
timestamp 1713453518
transform 1 0 1820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4040
timestamp 1713453518
transform 1 0 1620 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4041
timestamp 1713453518
transform 1 0 1620 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1713453518
transform 1 0 1652 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1713453518
transform 1 0 1636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1713453518
transform 1 0 1364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1713453518
transform 1 0 1324 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1713453518
transform 1 0 1308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1713453518
transform 1 0 1308 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1713453518
transform 1 0 1244 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1713453518
transform 1 0 1204 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1713453518
transform 1 0 1188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1713453518
transform 1 0 1972 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1713453518
transform 1 0 1972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4053
timestamp 1713453518
transform 1 0 1772 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1713453518
transform 1 0 1772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1713453518
transform 1 0 3196 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4056
timestamp 1713453518
transform 1 0 3148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1713453518
transform 1 0 3140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1713453518
transform 1 0 3140 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1713453518
transform 1 0 3140 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1713453518
transform 1 0 2916 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1713453518
transform 1 0 1828 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1713453518
transform 1 0 1788 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1713453518
transform 1 0 1372 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1713453518
transform 1 0 1332 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1713453518
transform 1 0 1316 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1713453518
transform 1 0 1268 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1713453518
transform 1 0 1228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1713453518
transform 1 0 1276 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4069
timestamp 1713453518
transform 1 0 1268 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1713453518
transform 1 0 1220 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1713453518
transform 1 0 1172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1713453518
transform 1 0 1508 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1713453518
transform 1 0 892 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1713453518
transform 1 0 1572 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1713453518
transform 1 0 1484 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1713453518
transform 1 0 1492 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4077
timestamp 1713453518
transform 1 0 1492 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4078
timestamp 1713453518
transform 1 0 1428 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4079
timestamp 1713453518
transform 1 0 1412 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1713453518
transform 1 0 1204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1713453518
transform 1 0 1524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4082
timestamp 1713453518
transform 1 0 1492 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1713453518
transform 1 0 3228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4084
timestamp 1713453518
transform 1 0 3204 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4085
timestamp 1713453518
transform 1 0 2996 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1713453518
transform 1 0 2916 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4087
timestamp 1713453518
transform 1 0 2028 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1713453518
transform 1 0 1580 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1713453518
transform 1 0 1596 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4090
timestamp 1713453518
transform 1 0 1172 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1713453518
transform 1 0 1156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1713453518
transform 1 0 1140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4093
timestamp 1713453518
transform 1 0 1132 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4094
timestamp 1713453518
transform 1 0 1132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1713453518
transform 1 0 1092 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1713453518
transform 1 0 1052 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1713453518
transform 1 0 1844 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1713453518
transform 1 0 1548 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1713453518
transform 1 0 1628 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1713453518
transform 1 0 1556 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1713453518
transform 1 0 1652 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4102
timestamp 1713453518
transform 1 0 1636 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1713453518
transform 1 0 1372 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1713453518
transform 1 0 1356 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1713453518
transform 1 0 1356 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4106
timestamp 1713453518
transform 1 0 1292 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1713453518
transform 1 0 1268 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1713453518
transform 1 0 1260 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1713453518
transform 1 0 1204 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1713453518
transform 1 0 1148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1713453518
transform 1 0 1476 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4112
timestamp 1713453518
transform 1 0 908 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1713453518
transform 1 0 1956 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1713453518
transform 1 0 1452 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1713453518
transform 1 0 1468 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1713453518
transform 1 0 1460 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4117
timestamp 1713453518
transform 1 0 1396 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1713453518
transform 1 0 1388 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1713453518
transform 1 0 1380 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4120
timestamp 1713453518
transform 1 0 1308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1713453518
transform 1 0 1732 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1713453518
transform 1 0 1500 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1713453518
transform 1 0 3116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4124
timestamp 1713453518
transform 1 0 3092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4125
timestamp 1713453518
transform 1 0 3084 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4126
timestamp 1713453518
transform 1 0 2796 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1713453518
transform 1 0 2700 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4128
timestamp 1713453518
transform 1 0 2428 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4129
timestamp 1713453518
transform 1 0 1812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1713453518
transform 1 0 1860 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4131
timestamp 1713453518
transform 1 0 1244 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4132
timestamp 1713453518
transform 1 0 1300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4133
timestamp 1713453518
transform 1 0 1276 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4134
timestamp 1713453518
transform 1 0 1180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1713453518
transform 1 0 1148 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1713453518
transform 1 0 1100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4137
timestamp 1713453518
transform 1 0 1100 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4138
timestamp 1713453518
transform 1 0 1084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4139
timestamp 1713453518
transform 1 0 1028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4140
timestamp 1713453518
transform 1 0 2012 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1713453518
transform 1 0 1932 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1713453518
transform 1 0 2100 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4143
timestamp 1713453518
transform 1 0 1940 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4144
timestamp 1713453518
transform 1 0 2124 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4145
timestamp 1713453518
transform 1 0 2108 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4146
timestamp 1713453518
transform 1 0 1444 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4147
timestamp 1713453518
transform 1 0 2396 0 1 2955
box -2 -2 2 2
use M2_M1  M2_M1_4148
timestamp 1713453518
transform 1 0 2396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1713453518
transform 1 0 2364 0 1 2955
box -2 -2 2 2
use M2_M1  M2_M1_4150
timestamp 1713453518
transform 1 0 2060 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4151
timestamp 1713453518
transform 1 0 2012 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4152
timestamp 1713453518
transform 1 0 2012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1713453518
transform 1 0 1956 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4154
timestamp 1713453518
transform 1 0 1388 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4155
timestamp 1713453518
transform 1 0 1356 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4156
timestamp 1713453518
transform 1 0 1308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4157
timestamp 1713453518
transform 1 0 1300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4158
timestamp 1713453518
transform 1 0 1292 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4159
timestamp 1713453518
transform 1 0 1244 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4160
timestamp 1713453518
transform 1 0 1860 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4161
timestamp 1713453518
transform 1 0 1108 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1713453518
transform 1 0 2812 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4163
timestamp 1713453518
transform 1 0 1820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4164
timestamp 1713453518
transform 1 0 1868 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4165
timestamp 1713453518
transform 1 0 1828 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4166
timestamp 1713453518
transform 1 0 1924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4167
timestamp 1713453518
transform 1 0 1924 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4168
timestamp 1713453518
transform 1 0 2252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4169
timestamp 1713453518
transform 1 0 1996 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4170
timestamp 1713453518
transform 1 0 2012 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4171
timestamp 1713453518
transform 1 0 2012 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4172
timestamp 1713453518
transform 1 0 1572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4173
timestamp 1713453518
transform 1 0 1500 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1713453518
transform 1 0 1492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4175
timestamp 1713453518
transform 1 0 1460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4176
timestamp 1713453518
transform 1 0 1308 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4177
timestamp 1713453518
transform 1 0 1284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4178
timestamp 1713453518
transform 1 0 1220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4179
timestamp 1713453518
transform 1 0 1148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4180
timestamp 1713453518
transform 1 0 1404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4181
timestamp 1713453518
transform 1 0 1276 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4182
timestamp 1713453518
transform 1 0 2972 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4183
timestamp 1713453518
transform 1 0 1468 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4184
timestamp 1713453518
transform 1 0 1316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4185
timestamp 1713453518
transform 1 0 1268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4186
timestamp 1713453518
transform 1 0 1252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4187
timestamp 1713453518
transform 1 0 1084 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4188
timestamp 1713453518
transform 1 0 1076 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4189
timestamp 1713453518
transform 1 0 1044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4190
timestamp 1713453518
transform 1 0 2828 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4191
timestamp 1713453518
transform 1 0 2820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4192
timestamp 1713453518
transform 1 0 2868 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4193
timestamp 1713453518
transform 1 0 2836 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1713453518
transform 1 0 2868 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_4195
timestamp 1713453518
transform 1 0 2836 0 1 2985
box -2 -2 2 2
use M2_M1  M2_M1_4196
timestamp 1713453518
transform 1 0 2812 0 1 2985
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1713453518
transform 1 0 2812 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1713453518
transform 1 0 1300 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4199
timestamp 1713453518
transform 1 0 1284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1713453518
transform 1 0 1284 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1713453518
transform 1 0 1260 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4202
timestamp 1713453518
transform 1 0 1268 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4203
timestamp 1713453518
transform 1 0 1268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4204
timestamp 1713453518
transform 1 0 2548 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4205
timestamp 1713453518
transform 1 0 1116 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1713453518
transform 1 0 3140 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4207
timestamp 1713453518
transform 1 0 2516 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4208
timestamp 1713453518
transform 1 0 2468 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4209
timestamp 1713453518
transform 1 0 2468 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4210
timestamp 1713453518
transform 1 0 2428 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4211
timestamp 1713453518
transform 1 0 2100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4212
timestamp 1713453518
transform 1 0 2636 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4213
timestamp 1713453518
transform 1 0 2524 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1713453518
transform 1 0 2972 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4215
timestamp 1713453518
transform 1 0 2548 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4216
timestamp 1713453518
transform 1 0 2284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4217
timestamp 1713453518
transform 1 0 1716 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1713453518
transform 1 0 1436 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4219
timestamp 1713453518
transform 1 0 1148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4220
timestamp 1713453518
transform 1 0 1132 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4221
timestamp 1713453518
transform 1 0 1124 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1713453518
transform 1 0 1084 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1713453518
transform 1 0 1084 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4224
timestamp 1713453518
transform 1 0 1060 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4225
timestamp 1713453518
transform 1 0 1060 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4226
timestamp 1713453518
transform 1 0 3252 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1713453518
transform 1 0 3124 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1713453518
transform 1 0 3148 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_4229
timestamp 1713453518
transform 1 0 3132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1713453518
transform 1 0 3124 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_4231
timestamp 1713453518
transform 1 0 3116 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1713453518
transform 1 0 3084 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4233
timestamp 1713453518
transform 1 0 3068 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1713453518
transform 1 0 2204 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1713453518
transform 1 0 2204 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4236
timestamp 1713453518
transform 1 0 2148 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1713453518
transform 1 0 1404 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1713453518
transform 1 0 3172 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4239
timestamp 1713453518
transform 1 0 1348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4240
timestamp 1713453518
transform 1 0 1436 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4241
timestamp 1713453518
transform 1 0 1420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4242
timestamp 1713453518
transform 1 0 1284 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4243
timestamp 1713453518
transform 1 0 1268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4244
timestamp 1713453518
transform 1 0 1292 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4245
timestamp 1713453518
transform 1 0 1292 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4246
timestamp 1713453518
transform 1 0 1532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4247
timestamp 1713453518
transform 1 0 1516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1713453518
transform 1 0 1508 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1713453518
transform 1 0 1332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1713453518
transform 1 0 1268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4251
timestamp 1713453518
transform 1 0 1236 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4252
timestamp 1713453518
transform 1 0 1220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1713453518
transform 1 0 1188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4254
timestamp 1713453518
transform 1 0 1172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4255
timestamp 1713453518
transform 1 0 2564 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4256
timestamp 1713453518
transform 1 0 1148 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4257
timestamp 1713453518
transform 1 0 3332 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4258
timestamp 1713453518
transform 1 0 2540 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4259
timestamp 1713453518
transform 1 0 2564 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1713453518
transform 1 0 2548 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4261
timestamp 1713453518
transform 1 0 2572 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1713453518
transform 1 0 2388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1713453518
transform 1 0 2748 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4264
timestamp 1713453518
transform 1 0 2644 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4265
timestamp 1713453518
transform 1 0 3196 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4266
timestamp 1713453518
transform 1 0 3164 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4267
timestamp 1713453518
transform 1 0 3164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4268
timestamp 1713453518
transform 1 0 3124 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1713453518
transform 1 0 2940 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4270
timestamp 1713453518
transform 1 0 2796 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4271
timestamp 1713453518
transform 1 0 2636 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4272
timestamp 1713453518
transform 1 0 2596 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4273
timestamp 1713453518
transform 1 0 2476 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_4274
timestamp 1713453518
transform 1 0 2476 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1713453518
transform 1 0 2452 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_4276
timestamp 1713453518
transform 1 0 1860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1713453518
transform 1 0 1756 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4278
timestamp 1713453518
transform 1 0 1188 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4279
timestamp 1713453518
transform 1 0 2948 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1713453518
transform 1 0 2820 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4281
timestamp 1713453518
transform 1 0 2676 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4282
timestamp 1713453518
transform 1 0 3364 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1713453518
transform 1 0 3196 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_4284
timestamp 1713453518
transform 1 0 3196 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_4285
timestamp 1713453518
transform 1 0 2940 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1713453518
transform 1 0 2764 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4287
timestamp 1713453518
transform 1 0 3372 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4288
timestamp 1713453518
transform 1 0 3348 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4289
timestamp 1713453518
transform 1 0 3012 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4290
timestamp 1713453518
transform 1 0 2420 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4291
timestamp 1713453518
transform 1 0 1180 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4292
timestamp 1713453518
transform 1 0 1164 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1713453518
transform 1 0 1156 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4294
timestamp 1713453518
transform 1 0 1036 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1713453518
transform 1 0 1124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1713453518
transform 1 0 1020 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4297
timestamp 1713453518
transform 1 0 1020 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4298
timestamp 1713453518
transform 1 0 988 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4299
timestamp 1713453518
transform 1 0 988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1713453518
transform 1 0 3316 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4301
timestamp 1713453518
transform 1 0 3316 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1713453518
transform 1 0 3340 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4303
timestamp 1713453518
transform 1 0 3324 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1713453518
transform 1 0 3308 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1713453518
transform 1 0 3284 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1713453518
transform 1 0 3228 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4307
timestamp 1713453518
transform 1 0 3068 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1713453518
transform 1 0 2644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4309
timestamp 1713453518
transform 1 0 2620 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4310
timestamp 1713453518
transform 1 0 2476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1713453518
transform 1 0 1388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4312
timestamp 1713453518
transform 1 0 2764 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1713453518
transform 1 0 2748 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1713453518
transform 1 0 2740 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1713453518
transform 1 0 2732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4316
timestamp 1713453518
transform 1 0 2692 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1713453518
transform 1 0 2580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4318
timestamp 1713453518
transform 1 0 1276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4319
timestamp 1713453518
transform 1 0 3244 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4320
timestamp 1713453518
transform 1 0 3236 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1713453518
transform 1 0 3212 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4322
timestamp 1713453518
transform 1 0 3196 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4323
timestamp 1713453518
transform 1 0 3196 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4324
timestamp 1713453518
transform 1 0 3124 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4325
timestamp 1713453518
transform 1 0 3084 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4326
timestamp 1713453518
transform 1 0 3076 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4327
timestamp 1713453518
transform 1 0 3076 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4328
timestamp 1713453518
transform 1 0 2516 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1713453518
transform 1 0 1124 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1713453518
transform 1 0 3116 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4331
timestamp 1713453518
transform 1 0 2492 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1713453518
transform 1 0 2516 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1713453518
transform 1 0 2500 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4334
timestamp 1713453518
transform 1 0 2524 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1713453518
transform 1 0 2316 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1713453518
transform 1 0 2732 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1713453518
transform 1 0 2628 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4338
timestamp 1713453518
transform 1 0 2884 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1713453518
transform 1 0 2844 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1713453518
transform 1 0 2828 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4341
timestamp 1713453518
transform 1 0 3388 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_4342
timestamp 1713453518
transform 1 0 3364 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_4343
timestamp 1713453518
transform 1 0 3052 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_4344
timestamp 1713453518
transform 1 0 2924 0 1 3305
box -2 -2 2 2
use M2_M1  M2_M1_4345
timestamp 1713453518
transform 1 0 2924 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_4346
timestamp 1713453518
transform 1 0 3348 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4347
timestamp 1713453518
transform 1 0 3300 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4348
timestamp 1713453518
transform 1 0 2540 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4349
timestamp 1713453518
transform 1 0 2436 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1713453518
transform 1 0 2260 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4351
timestamp 1713453518
transform 1 0 1276 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4352
timestamp 1713453518
transform 1 0 1140 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4353
timestamp 1713453518
transform 1 0 1140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1713453518
transform 1 0 1116 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4355
timestamp 1713453518
transform 1 0 1076 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4356
timestamp 1713453518
transform 1 0 1020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4357
timestamp 1713453518
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4358
timestamp 1713453518
transform 1 0 3388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_4359
timestamp 1713453518
transform 1 0 3124 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_4360
timestamp 1713453518
transform 1 0 3156 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_4361
timestamp 1713453518
transform 1 0 3156 0 1 3245
box -2 -2 2 2
use M2_M1  M2_M1_4362
timestamp 1713453518
transform 1 0 3156 0 1 3345
box -2 -2 2 2
use M2_M1  M2_M1_4363
timestamp 1713453518
transform 1 0 3132 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_4364
timestamp 1713453518
transform 1 0 2780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4365
timestamp 1713453518
transform 1 0 2748 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4366
timestamp 1713453518
transform 1 0 2716 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4367
timestamp 1713453518
transform 1 0 2484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4368
timestamp 1713453518
transform 1 0 2468 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1713453518
transform 1 0 2444 0 1 1445
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1713453518
transform 1 0 1308 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1713453518
transform 1 0 2804 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_4372
timestamp 1713453518
transform 1 0 2804 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1713453518
transform 1 0 2804 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4374
timestamp 1713453518
transform 1 0 2788 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_4375
timestamp 1713453518
transform 1 0 2460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1713453518
transform 1 0 1260 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1713453518
transform 1 0 2564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4378
timestamp 1713453518
transform 1 0 1068 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4379
timestamp 1713453518
transform 1 0 3236 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1713453518
transform 1 0 2540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1713453518
transform 1 0 2452 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4382
timestamp 1713453518
transform 1 0 2140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4383
timestamp 1713453518
transform 1 0 2628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4384
timestamp 1713453518
transform 1 0 2532 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4385
timestamp 1713453518
transform 1 0 3100 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4386
timestamp 1713453518
transform 1 0 3092 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4387
timestamp 1713453518
transform 1 0 3020 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4388
timestamp 1713453518
transform 1 0 3020 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4389
timestamp 1713453518
transform 1 0 3004 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4390
timestamp 1713453518
transform 1 0 2924 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4391
timestamp 1713453518
transform 1 0 2796 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4392
timestamp 1713453518
transform 1 0 2660 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4393
timestamp 1713453518
transform 1 0 2596 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4394
timestamp 1713453518
transform 1 0 2580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4395
timestamp 1713453518
transform 1 0 2348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1713453518
transform 1 0 3332 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_4397
timestamp 1713453518
transform 1 0 3300 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4398
timestamp 1713453518
transform 1 0 3052 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_4399
timestamp 1713453518
transform 1 0 2668 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_4400
timestamp 1713453518
transform 1 0 1516 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1713453518
transform 1 0 2276 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1713453518
transform 1 0 1508 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1713453518
transform 1 0 3292 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4404
timestamp 1713453518
transform 1 0 3244 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1713453518
transform 1 0 2356 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_4406
timestamp 1713453518
transform 1 0 2356 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_4407
timestamp 1713453518
transform 1 0 3324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4408
timestamp 1713453518
transform 1 0 3212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4409
timestamp 1713453518
transform 1 0 3236 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_4410
timestamp 1713453518
transform 1 0 3212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4411
timestamp 1713453518
transform 1 0 3212 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_4412
timestamp 1713453518
transform 1 0 3180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_4413
timestamp 1713453518
transform 1 0 1548 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4414
timestamp 1713453518
transform 1 0 1436 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4415
timestamp 1713453518
transform 1 0 1476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4416
timestamp 1713453518
transform 1 0 1316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4417
timestamp 1713453518
transform 1 0 1324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4418
timestamp 1713453518
transform 1 0 1292 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4419
timestamp 1713453518
transform 1 0 1916 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4420
timestamp 1713453518
transform 1 0 1092 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4421
timestamp 1713453518
transform 1 0 3268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1713453518
transform 1 0 1876 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4423
timestamp 1713453518
transform 1 0 2028 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4424
timestamp 1713453518
transform 1 0 1884 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1713453518
transform 1 0 2076 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4426
timestamp 1713453518
transform 1 0 1996 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1713453518
transform 1 0 2444 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4428
timestamp 1713453518
transform 1 0 2124 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1713453518
transform 1 0 3332 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4430
timestamp 1713453518
transform 1 0 3308 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4431
timestamp 1713453518
transform 1 0 3132 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_4432
timestamp 1713453518
transform 1 0 2436 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1713453518
transform 1 0 1628 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4434
timestamp 1713453518
transform 1 0 1540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4435
timestamp 1713453518
transform 1 0 1492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4436
timestamp 1713453518
transform 1 0 1556 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1713453518
transform 1 0 1124 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4438
timestamp 1713453518
transform 1 0 1524 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4439
timestamp 1713453518
transform 1 0 1516 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4440
timestamp 1713453518
transform 1 0 1444 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4441
timestamp 1713453518
transform 1 0 1388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4442
timestamp 1713453518
transform 1 0 1372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4443
timestamp 1713453518
transform 1 0 1372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1713453518
transform 1 0 3364 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1713453518
transform 1 0 3236 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4446
timestamp 1713453518
transform 1 0 3252 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4447
timestamp 1713453518
transform 1 0 3236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1713453518
transform 1 0 3212 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_4449
timestamp 1713453518
transform 1 0 3092 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4450
timestamp 1713453518
transform 1 0 3036 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4451
timestamp 1713453518
transform 1 0 3012 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1713453518
transform 1 0 1644 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4453
timestamp 1713453518
transform 1 0 1364 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1713453518
transform 1 0 1604 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4455
timestamp 1713453518
transform 1 0 1388 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1713453518
transform 1 0 1396 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4457
timestamp 1713453518
transform 1 0 1396 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4458
timestamp 1713453518
transform 1 0 1564 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4459
timestamp 1713453518
transform 1 0 1348 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4460
timestamp 1713453518
transform 1 0 1348 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4461
timestamp 1713453518
transform 1 0 1348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4462
timestamp 1713453518
transform 1 0 1324 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1713453518
transform 1 0 1188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1713453518
transform 1 0 1852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1713453518
transform 1 0 1052 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4466
timestamp 1713453518
transform 1 0 3268 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4467
timestamp 1713453518
transform 1 0 1812 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4468
timestamp 1713453518
transform 1 0 1820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4469
timestamp 1713453518
transform 1 0 1820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4470
timestamp 1713453518
transform 1 0 1924 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4471
timestamp 1713453518
transform 1 0 1836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1713453518
transform 1 0 2460 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1713453518
transform 1 0 1892 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4474
timestamp 1713453518
transform 1 0 3300 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1713453518
transform 1 0 3284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4476
timestamp 1713453518
transform 1 0 3284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1713453518
transform 1 0 3268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4478
timestamp 1713453518
transform 1 0 3252 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4479
timestamp 1713453518
transform 1 0 3252 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4480
timestamp 1713453518
transform 1 0 3156 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1713453518
transform 1 0 3140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4482
timestamp 1713453518
transform 1 0 2884 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4483
timestamp 1713453518
transform 1 0 2796 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1713453518
transform 1 0 2556 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4485
timestamp 1713453518
transform 1 0 2508 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1713453518
transform 1 0 1692 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1713453518
transform 1 0 2628 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4488
timestamp 1713453518
transform 1 0 2532 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4489
timestamp 1713453518
transform 1 0 1540 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1713453518
transform 1 0 3412 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1713453518
transform 1 0 3348 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4492
timestamp 1713453518
transform 1 0 3156 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_4493
timestamp 1713453518
transform 1 0 2540 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_4494
timestamp 1713453518
transform 1 0 1468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1713453518
transform 1 0 1724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1713453518
transform 1 0 1700 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4497
timestamp 1713453518
transform 1 0 1596 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4498
timestamp 1713453518
transform 1 0 1572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4499
timestamp 1713453518
transform 1 0 1644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1713453518
transform 1 0 1116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1713453518
transform 1 0 1508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4502
timestamp 1713453518
transform 1 0 1508 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1713453518
transform 1 0 1228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4504
timestamp 1713453518
transform 1 0 1228 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4505
timestamp 1713453518
transform 1 0 1228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4506
timestamp 1713453518
transform 1 0 1172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4507
timestamp 1713453518
transform 1 0 3420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4508
timestamp 1713453518
transform 1 0 3260 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4509
timestamp 1713453518
transform 1 0 3276 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4510
timestamp 1713453518
transform 1 0 3260 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4511
timestamp 1713453518
transform 1 0 3236 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_4512
timestamp 1713453518
transform 1 0 3148 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4513
timestamp 1713453518
transform 1 0 3092 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1713453518
transform 1 0 2796 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4515
timestamp 1713453518
transform 1 0 1548 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1713453518
transform 1 0 1420 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1713453518
transform 1 0 1428 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4518
timestamp 1713453518
transform 1 0 1340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4519
timestamp 1713453518
transform 1 0 1308 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4520
timestamp 1713453518
transform 1 0 1292 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1713453518
transform 1 0 1588 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1713453518
transform 1 0 1548 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1713453518
transform 1 0 1484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4524
timestamp 1713453518
transform 1 0 1204 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4525
timestamp 1713453518
transform 1 0 1188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1713453518
transform 1 0 1188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1713453518
transform 1 0 1276 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1713453518
transform 1 0 1180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4529
timestamp 1713453518
transform 1 0 2020 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4530
timestamp 1713453518
transform 1 0 1044 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4531
timestamp 1713453518
transform 1 0 2892 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1713453518
transform 1 0 1988 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1713453518
transform 1 0 2028 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1713453518
transform 1 0 2004 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4535
timestamp 1713453518
transform 1 0 2028 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4536
timestamp 1713453518
transform 1 0 2004 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4537
timestamp 1713453518
transform 1 0 2364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4538
timestamp 1713453518
transform 1 0 2100 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4539
timestamp 1713453518
transform 1 0 3020 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4540
timestamp 1713453518
transform 1 0 2892 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4541
timestamp 1713453518
transform 1 0 2692 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1713453518
transform 1 0 2444 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4543
timestamp 1713453518
transform 1 0 1748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4544
timestamp 1713453518
transform 1 0 1892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4545
timestamp 1713453518
transform 1 0 1860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1713453518
transform 1 0 1788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4547
timestamp 1713453518
transform 1 0 1548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4548
timestamp 1713453518
transform 1 0 1724 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1713453518
transform 1 0 1156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4550
timestamp 1713453518
transform 1 0 1508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1713453518
transform 1 0 1508 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4552
timestamp 1713453518
transform 1 0 1492 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4553
timestamp 1713453518
transform 1 0 1476 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4554
timestamp 1713453518
transform 1 0 1348 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4555
timestamp 1713453518
transform 1 0 1244 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4556
timestamp 1713453518
transform 1 0 1236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4557
timestamp 1713453518
transform 1 0 2988 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4558
timestamp 1713453518
transform 1 0 2860 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4559
timestamp 1713453518
transform 1 0 2876 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4560
timestamp 1713453518
transform 1 0 2860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4561
timestamp 1713453518
transform 1 0 2852 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_4562
timestamp 1713453518
transform 1 0 2796 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4563
timestamp 1713453518
transform 1 0 2756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1713453518
transform 1 0 2644 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4565
timestamp 1713453518
transform 1 0 1828 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4566
timestamp 1713453518
transform 1 0 1636 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1713453518
transform 1 0 1724 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4568
timestamp 1713453518
transform 1 0 1628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1713453518
transform 1 0 1580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4570
timestamp 1713453518
transform 1 0 1564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1713453518
transform 1 0 1596 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4572
timestamp 1713453518
transform 1 0 1572 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1713453518
transform 1 0 1540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4574
timestamp 1713453518
transform 1 0 1500 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4575
timestamp 1713453518
transform 1 0 1492 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4576
timestamp 1713453518
transform 1 0 1460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4577
timestamp 1713453518
transform 1 0 1292 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1713453518
transform 1 0 1292 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1713453518
transform 1 0 1532 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1713453518
transform 1 0 1452 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1713453518
transform 1 0 2196 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4582
timestamp 1713453518
transform 1 0 1092 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1713453518
transform 1 0 2828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4584
timestamp 1713453518
transform 1 0 2172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4585
timestamp 1713453518
transform 1 0 2124 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4586
timestamp 1713453518
transform 1 0 2124 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4587
timestamp 1713453518
transform 1 0 2092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4588
timestamp 1713453518
transform 1 0 2084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4589
timestamp 1713453518
transform 1 0 2316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4590
timestamp 1713453518
transform 1 0 2100 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4591
timestamp 1713453518
transform 1 0 2932 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1713453518
transform 1 0 2892 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4593
timestamp 1713453518
transform 1 0 2828 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4594
timestamp 1713453518
transform 1 0 2348 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4595
timestamp 1713453518
transform 1 0 1740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4596
timestamp 1713453518
transform 1 0 1868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4597
timestamp 1713453518
transform 1 0 1772 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1713453518
transform 1 0 1644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4599
timestamp 1713453518
transform 1 0 1604 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1713453518
transform 1 0 1652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4601
timestamp 1713453518
transform 1 0 1140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4602
timestamp 1713453518
transform 1 0 1588 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4603
timestamp 1713453518
transform 1 0 1572 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4604
timestamp 1713453518
transform 1 0 1396 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1713453518
transform 1 0 1372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4606
timestamp 1713453518
transform 1 0 3012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4607
timestamp 1713453518
transform 1 0 2796 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1713453518
transform 1 0 2812 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4609
timestamp 1713453518
transform 1 0 2796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4610
timestamp 1713453518
transform 1 0 2788 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1713453518
transform 1 0 2756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4612
timestamp 1713453518
transform 1 0 1756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1713453518
transform 1 0 1620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4614
timestamp 1713453518
transform 1 0 1716 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4615
timestamp 1713453518
transform 1 0 1340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4616
timestamp 1713453518
transform 1 0 1356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4617
timestamp 1713453518
transform 1 0 1316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1713453518
transform 1 0 1308 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4619
timestamp 1713453518
transform 1 0 1268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1713453518
transform 1 0 1268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1713453518
transform 1 0 1260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4622
timestamp 1713453518
transform 1 0 1236 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4623
timestamp 1713453518
transform 1 0 1332 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4624
timestamp 1713453518
transform 1 0 1308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4625
timestamp 1713453518
transform 1 0 1212 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4626
timestamp 1713453518
transform 1 0 1204 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4627
timestamp 1713453518
transform 1 0 1756 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4628
timestamp 1713453518
transform 1 0 1748 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1713453518
transform 1 0 1716 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4630
timestamp 1713453518
transform 1 0 1596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4631
timestamp 1713453518
transform 1 0 1508 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4632
timestamp 1713453518
transform 1 0 1212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1713453518
transform 1 0 1172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4634
timestamp 1713453518
transform 1 0 1172 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4635
timestamp 1713453518
transform 1 0 2100 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4636
timestamp 1713453518
transform 1 0 1068 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4637
timestamp 1713453518
transform 1 0 3028 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1713453518
transform 1 0 2060 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4639
timestamp 1713453518
transform 1 0 2092 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4640
timestamp 1713453518
transform 1 0 2076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4641
timestamp 1713453518
transform 1 0 2148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4642
timestamp 1713453518
transform 1 0 2140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4643
timestamp 1713453518
transform 1 0 2316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1713453518
transform 1 0 2156 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1713453518
transform 1 0 2540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4646
timestamp 1713453518
transform 1 0 2460 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4647
timestamp 1713453518
transform 1 0 2276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4648
timestamp 1713453518
transform 1 0 3316 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4649
timestamp 1713453518
transform 1 0 3076 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4650
timestamp 1713453518
transform 1 0 2908 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_4651
timestamp 1713453518
transform 1 0 2564 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4652
timestamp 1713453518
transform 1 0 1460 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4653
timestamp 1713453518
transform 1 0 2012 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1713453518
transform 1 0 1716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1713453518
transform 1 0 1644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1713453518
transform 1 0 1116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4657
timestamp 1713453518
transform 1 0 3148 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1713453518
transform 1 0 3004 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4659
timestamp 1713453518
transform 1 0 3020 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1713453518
transform 1 0 3004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4661
timestamp 1713453518
transform 1 0 2964 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_4662
timestamp 1713453518
transform 1 0 2940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4663
timestamp 1713453518
transform 1 0 1428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4664
timestamp 1713453518
transform 1 0 1428 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1713453518
transform 1 0 1428 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4666
timestamp 1713453518
transform 1 0 1396 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4667
timestamp 1713453518
transform 1 0 1812 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4668
timestamp 1713453518
transform 1 0 1012 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1713453518
transform 1 0 3300 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4670
timestamp 1713453518
transform 1 0 1788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4671
timestamp 1713453518
transform 1 0 1812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4672
timestamp 1713453518
transform 1 0 1796 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1713453518
transform 1 0 1940 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1713453518
transform 1 0 1860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4675
timestamp 1713453518
transform 1 0 2460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4676
timestamp 1713453518
transform 1 0 1876 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4677
timestamp 1713453518
transform 1 0 3340 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1713453518
transform 1 0 3316 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4679
timestamp 1713453518
transform 1 0 3092 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_4680
timestamp 1713453518
transform 1 0 2796 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1713453518
transform 1 0 2772 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_4682
timestamp 1713453518
transform 1 0 2044 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4683
timestamp 1713453518
transform 1 0 1772 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4684
timestamp 1713453518
transform 1 0 1668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4685
timestamp 1713453518
transform 1 0 1564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1713453518
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1713453518
transform 1 0 1076 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4688
timestamp 1713453518
transform 1 0 3412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4689
timestamp 1713453518
transform 1 0 3292 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1713453518
transform 1 0 3316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4691
timestamp 1713453518
transform 1 0 3260 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4692
timestamp 1713453518
transform 1 0 3228 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_4693
timestamp 1713453518
transform 1 0 3116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4694
timestamp 1713453518
transform 1 0 3340 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4695
timestamp 1713453518
transform 1 0 3332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1713453518
transform 1 0 3300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1713453518
transform 1 0 3268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1713453518
transform 1 0 3252 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4699
timestamp 1713453518
transform 1 0 3252 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4700
timestamp 1713453518
transform 1 0 3140 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_4701
timestamp 1713453518
transform 1 0 3140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4702
timestamp 1713453518
transform 1 0 3132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4703
timestamp 1713453518
transform 1 0 3108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1713453518
transform 1 0 3108 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1713453518
transform 1 0 3108 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1713453518
transform 1 0 3100 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4707
timestamp 1713453518
transform 1 0 2508 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1713453518
transform 1 0 1028 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4709
timestamp 1713453518
transform 1 0 3284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1713453518
transform 1 0 2468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4711
timestamp 1713453518
transform 1 0 2404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4712
timestamp 1713453518
transform 1 0 2372 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1713453518
transform 1 0 2572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1713453518
transform 1 0 2468 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1713453518
transform 1 0 3172 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4716
timestamp 1713453518
transform 1 0 3172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4717
timestamp 1713453518
transform 1 0 3116 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1713453518
transform 1 0 3108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1713453518
transform 1 0 2996 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4720
timestamp 1713453518
transform 1 0 2940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1713453518
transform 1 0 2876 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1713453518
transform 1 0 2708 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1713453518
transform 1 0 2684 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4724
timestamp 1713453518
transform 1 0 2684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4725
timestamp 1713453518
transform 1 0 2452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1713453518
transform 1 0 1836 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1713453518
transform 1 0 2908 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1713453518
transform 1 0 2764 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1713453518
transform 1 0 2756 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1713453518
transform 1 0 3348 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4731
timestamp 1713453518
transform 1 0 3324 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4732
timestamp 1713453518
transform 1 0 3132 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4733
timestamp 1713453518
transform 1 0 2892 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1713453518
transform 1 0 2356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4735
timestamp 1713453518
transform 1 0 1836 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4736
timestamp 1713453518
transform 1 0 1724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1713453518
transform 1 0 1604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4738
timestamp 1713453518
transform 1 0 1732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4739
timestamp 1713453518
transform 1 0 1124 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1713453518
transform 1 0 3412 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4741
timestamp 1713453518
transform 1 0 3244 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1713453518
transform 1 0 3260 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1713453518
transform 1 0 3244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4744
timestamp 1713453518
transform 1 0 3228 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4745
timestamp 1713453518
transform 1 0 3180 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1713453518
transform 1 0 1772 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4747
timestamp 1713453518
transform 1 0 1700 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4748
timestamp 1713453518
transform 1 0 1612 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_4749
timestamp 1713453518
transform 1 0 1532 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4750
timestamp 1713453518
transform 1 0 1204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1713453518
transform 1 0 1204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4752
timestamp 1713453518
transform 1 0 1188 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1713453518
transform 1 0 2420 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1713453518
transform 1 0 1068 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1713453518
transform 1 0 3228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4756
timestamp 1713453518
transform 1 0 2348 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4757
timestamp 1713453518
transform 1 0 2420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1713453518
transform 1 0 2404 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4759
timestamp 1713453518
transform 1 0 2428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4760
timestamp 1713453518
transform 1 0 2148 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4761
timestamp 1713453518
transform 1 0 2524 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1713453518
transform 1 0 2508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4763
timestamp 1713453518
transform 1 0 2892 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4764
timestamp 1713453518
transform 1 0 2604 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1713453518
transform 1 0 1892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4766
timestamp 1713453518
transform 1 0 3316 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4767
timestamp 1713453518
transform 1 0 3284 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4768
timestamp 1713453518
transform 1 0 2908 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4769
timestamp 1713453518
transform 1 0 2644 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4770
timestamp 1713453518
transform 1 0 1420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4771
timestamp 1713453518
transform 1 0 2388 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1713453518
transform 1 0 1820 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4773
timestamp 1713453518
transform 1 0 1716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1713453518
transform 1 0 1716 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4775
timestamp 1713453518
transform 1 0 3412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4776
timestamp 1713453518
transform 1 0 3196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4777
timestamp 1713453518
transform 1 0 3228 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1713453518
transform 1 0 3204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4779
timestamp 1713453518
transform 1 0 3164 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4780
timestamp 1713453518
transform 1 0 3164 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4781
timestamp 1713453518
transform 1 0 1852 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4782
timestamp 1713453518
transform 1 0 1676 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1713453518
transform 1 0 1348 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4784
timestamp 1713453518
transform 1 0 1324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1713453518
transform 1 0 1332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4786
timestamp 1713453518
transform 1 0 1260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4787
timestamp 1713453518
transform 1 0 2356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4788
timestamp 1713453518
transform 1 0 1084 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1713453518
transform 1 0 2980 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4790
timestamp 1713453518
transform 1 0 2316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4791
timestamp 1713453518
transform 1 0 2244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4792
timestamp 1713453518
transform 1 0 2044 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4793
timestamp 1713453518
transform 1 0 2516 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1713453518
transform 1 0 2316 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4795
timestamp 1713453518
transform 1 0 3340 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4796
timestamp 1713453518
transform 1 0 3300 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1713453518
transform 1 0 2796 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1713453518
transform 1 0 2548 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4799
timestamp 1713453518
transform 1 0 1700 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4800
timestamp 1713453518
transform 1 0 1940 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4801
timestamp 1713453518
transform 1 0 1924 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4802
timestamp 1713453518
transform 1 0 1796 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4803
timestamp 1713453518
transform 1 0 1756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4804
timestamp 1713453518
transform 1 0 1844 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4805
timestamp 1713453518
transform 1 0 1164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4806
timestamp 1713453518
transform 1 0 1788 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4807
timestamp 1713453518
transform 1 0 1652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4808
timestamp 1713453518
transform 1 0 1588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4809
timestamp 1713453518
transform 1 0 1476 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4810
timestamp 1713453518
transform 1 0 1468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4811
timestamp 1713453518
transform 1 0 1444 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4812
timestamp 1713453518
transform 1 0 3348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4813
timestamp 1713453518
transform 1 0 3012 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4814
timestamp 1713453518
transform 1 0 3092 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4815
timestamp 1713453518
transform 1 0 3060 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4816
timestamp 1713453518
transform 1 0 3092 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1713453518
transform 1 0 2940 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4818
timestamp 1713453518
transform 1 0 2852 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_4819
timestamp 1713453518
transform 1 0 2852 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1713453518
transform 1 0 1772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4821
timestamp 1713453518
transform 1 0 1612 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4822
timestamp 1713453518
transform 1 0 1644 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4823
timestamp 1713453518
transform 1 0 1580 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4824
timestamp 1713453518
transform 1 0 1548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4825
timestamp 1713453518
transform 1 0 1540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4826
timestamp 1713453518
transform 1 0 1556 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4827
timestamp 1713453518
transform 1 0 1524 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4828
timestamp 1713453518
transform 1 0 1708 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4829
timestamp 1713453518
transform 1 0 1612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4830
timestamp 1713453518
transform 1 0 1476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1713453518
transform 1 0 1460 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1713453518
transform 1 0 1444 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4833
timestamp 1713453518
transform 1 0 1548 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4834
timestamp 1713453518
transform 1 0 1476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4835
timestamp 1713453518
transform 1 0 2372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1713453518
transform 1 0 1092 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1713453518
transform 1 0 3284 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4838
timestamp 1713453518
transform 1 0 2348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4839
timestamp 1713453518
transform 1 0 2260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4840
timestamp 1713453518
transform 1 0 2156 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4841
timestamp 1713453518
transform 1 0 2500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4842
timestamp 1713453518
transform 1 0 2324 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4843
timestamp 1713453518
transform 1 0 2716 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4844
timestamp 1713453518
transform 1 0 2604 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4845
timestamp 1713453518
transform 1 0 1764 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4846
timestamp 1713453518
transform 1 0 3316 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4847
timestamp 1713453518
transform 1 0 3284 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4848
timestamp 1713453518
transform 1 0 3132 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_4849
timestamp 1713453518
transform 1 0 2588 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_4850
timestamp 1713453518
transform 1 0 1804 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1713453518
transform 1 0 1844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4852
timestamp 1713453518
transform 1 0 1196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4853
timestamp 1713453518
transform 1 0 3356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4854
timestamp 1713453518
transform 1 0 3300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4855
timestamp 1713453518
transform 1 0 3316 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1713453518
transform 1 0 3244 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_4857
timestamp 1713453518
transform 1 0 3228 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4858
timestamp 1713453518
transform 1 0 3228 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1713453518
transform 1 0 3180 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4860
timestamp 1713453518
transform 1 0 3180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1713453518
transform 1 0 1724 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4862
timestamp 1713453518
transform 1 0 1580 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4863
timestamp 1713453518
transform 1 0 1764 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4864
timestamp 1713453518
transform 1 0 1700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4865
timestamp 1713453518
transform 1 0 1604 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4866
timestamp 1713453518
transform 1 0 1564 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4867
timestamp 1713453518
transform 1 0 1668 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1713453518
transform 1 0 1668 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1713453518
transform 1 0 1676 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4870
timestamp 1713453518
transform 1 0 1676 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4871
timestamp 1713453518
transform 1 0 1596 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4872
timestamp 1713453518
transform 1 0 1580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4873
timestamp 1713453518
transform 1 0 1412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4874
timestamp 1713453518
transform 1 0 1556 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_4875
timestamp 1713453518
transform 1 0 1508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4876
timestamp 1713453518
transform 1 0 2340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4877
timestamp 1713453518
transform 1 0 1060 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4878
timestamp 1713453518
transform 1 0 3068 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4879
timestamp 1713453518
transform 1 0 2316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4880
timestamp 1713453518
transform 1 0 2252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1713453518
transform 1 0 2124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1713453518
transform 1 0 2436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4883
timestamp 1713453518
transform 1 0 2308 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1713453518
transform 1 0 2596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4885
timestamp 1713453518
transform 1 0 2412 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4886
timestamp 1713453518
transform 1 0 1740 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1713453518
transform 1 0 3268 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1713453518
transform 1 0 3204 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4889
timestamp 1713453518
transform 1 0 2988 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1713453518
transform 1 0 2468 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_4891
timestamp 1713453518
transform 1 0 1780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4892
timestamp 1713453518
transform 1 0 2196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1713453518
transform 1 0 1868 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4894
timestamp 1713453518
transform 1 0 1756 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1713453518
transform 1 0 1692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4896
timestamp 1713453518
transform 1 0 1812 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1713453518
transform 1 0 1124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4898
timestamp 1713453518
transform 1 0 1652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4899
timestamp 1713453518
transform 1 0 1652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4900
timestamp 1713453518
transform 1 0 1628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1713453518
transform 1 0 1532 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4902
timestamp 1713453518
transform 1 0 1332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4903
timestamp 1713453518
transform 1 0 1252 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4904
timestamp 1713453518
transform 1 0 1244 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1713453518
transform 1 0 1180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4906
timestamp 1713453518
transform 1 0 3260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1713453518
transform 1 0 3044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4908
timestamp 1713453518
transform 1 0 3060 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4909
timestamp 1713453518
transform 1 0 3044 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4910
timestamp 1713453518
transform 1 0 3020 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1713453518
transform 1 0 2908 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1713453518
transform 1 0 1700 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4913
timestamp 1713453518
transform 1 0 1596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1713453518
transform 1 0 1764 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4915
timestamp 1713453518
transform 1 0 1572 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4916
timestamp 1713453518
transform 1 0 1556 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4917
timestamp 1713453518
transform 1 0 1556 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1713453518
transform 1 0 1612 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4919
timestamp 1713453518
transform 1 0 1516 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4920
timestamp 1713453518
transform 1 0 1508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1713453518
transform 1 0 1500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4922
timestamp 1713453518
transform 1 0 1316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4923
timestamp 1713453518
transform 1 0 1316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4924
timestamp 1713453518
transform 1 0 1492 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_4925
timestamp 1713453518
transform 1 0 1420 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4926
timestamp 1713453518
transform 1 0 1908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4927
timestamp 1713453518
transform 1 0 1052 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4928
timestamp 1713453518
transform 1 0 2636 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4929
timestamp 1713453518
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4930
timestamp 1713453518
transform 1 0 1908 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1713453518
transform 1 0 1892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1713453518
transform 1 0 2012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1713453518
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4934
timestamp 1713453518
transform 1 0 2380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1713453518
transform 1 0 1972 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4936
timestamp 1713453518
transform 1 0 2596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1713453518
transform 1 0 2324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4938
timestamp 1713453518
transform 1 0 1756 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4939
timestamp 1713453518
transform 1 0 2980 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4940
timestamp 1713453518
transform 1 0 2852 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4941
timestamp 1713453518
transform 1 0 2756 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4942
timestamp 1713453518
transform 1 0 2452 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1713453518
transform 1 0 2404 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4944
timestamp 1713453518
transform 1 0 1652 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4945
timestamp 1713453518
transform 1 0 2028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4946
timestamp 1713453518
transform 1 0 1868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4947
timestamp 1713453518
transform 1 0 1772 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1713453518
transform 1 0 1684 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4949
timestamp 1713453518
transform 1 0 1788 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4950
timestamp 1713453518
transform 1 0 1100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4951
timestamp 1713453518
transform 1 0 1676 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4952
timestamp 1713453518
transform 1 0 1668 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4953
timestamp 1713453518
transform 1 0 1316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4954
timestamp 1713453518
transform 1 0 1300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4955
timestamp 1713453518
transform 1 0 1292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4956
timestamp 1713453518
transform 1 0 2964 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1713453518
transform 1 0 2676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1713453518
transform 1 0 2756 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1713453518
transform 1 0 2708 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4960
timestamp 1713453518
transform 1 0 2756 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1713453518
transform 1 0 2756 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_4962
timestamp 1713453518
transform 1 0 1700 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1713453518
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4964
timestamp 1713453518
transform 1 0 1604 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4965
timestamp 1713453518
transform 1 0 1292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4966
timestamp 1713453518
transform 1 0 1132 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4967
timestamp 1713453518
transform 1 0 1092 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4968
timestamp 1713453518
transform 1 0 1276 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4969
timestamp 1713453518
transform 1 0 1252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1713453518
transform 1 0 1244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4971
timestamp 1713453518
transform 1 0 1188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4972
timestamp 1713453518
transform 1 0 1244 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4973
timestamp 1713453518
transform 1 0 1172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4974
timestamp 1713453518
transform 1 0 1692 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1713453518
transform 1 0 1652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4976
timestamp 1713453518
transform 1 0 1556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4977
timestamp 1713453518
transform 1 0 1532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4978
timestamp 1713453518
transform 1 0 1236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4979
timestamp 1713453518
transform 1 0 1228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4980
timestamp 1713453518
transform 1 0 1180 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1713453518
transform 1 0 1180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4982
timestamp 1713453518
transform 1 0 1156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4983
timestamp 1713453518
transform 1 0 1156 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_4984
timestamp 1713453518
transform 1 0 1852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4985
timestamp 1713453518
transform 1 0 1012 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4986
timestamp 1713453518
transform 1 0 2812 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4987
timestamp 1713453518
transform 1 0 1804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4988
timestamp 1713453518
transform 1 0 1964 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4989
timestamp 1713453518
transform 1 0 1828 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1713453518
transform 1 0 1948 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4991
timestamp 1713453518
transform 1 0 1916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4992
timestamp 1713453518
transform 1 0 2316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4993
timestamp 1713453518
transform 1 0 2028 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4994
timestamp 1713453518
transform 1 0 3412 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1713453518
transform 1 0 3356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4996
timestamp 1713453518
transform 1 0 3340 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1713453518
transform 1 0 2788 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4998
timestamp 1713453518
transform 1 0 2668 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4999
timestamp 1713453518
transform 1 0 2620 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5000
timestamp 1713453518
transform 1 0 2564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5001
timestamp 1713453518
transform 1 0 2524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1713453518
transform 1 0 2468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5003
timestamp 1713453518
transform 1 0 2444 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5004
timestamp 1713453518
transform 1 0 2236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5005
timestamp 1713453518
transform 1 0 1796 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5006
timestamp 1713453518
transform 1 0 2884 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5007
timestamp 1713453518
transform 1 0 2836 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1713453518
transform 1 0 2636 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_5009
timestamp 1713453518
transform 1 0 2444 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_5010
timestamp 1713453518
transform 1 0 1460 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5011
timestamp 1713453518
transform 1 0 1700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5012
timestamp 1713453518
transform 1 0 1684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5013
timestamp 1713453518
transform 1 0 1764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5014
timestamp 1713453518
transform 1 0 1084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5015
timestamp 1713453518
transform 1 0 2940 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5016
timestamp 1713453518
transform 1 0 2804 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5017
timestamp 1713453518
transform 1 0 2820 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5018
timestamp 1713453518
transform 1 0 2788 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5019
timestamp 1713453518
transform 1 0 2756 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5020
timestamp 1713453518
transform 1 0 2724 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5021
timestamp 1713453518
transform 1 0 1420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5022
timestamp 1713453518
transform 1 0 1420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5023
timestamp 1713453518
transform 1 0 1412 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1713453518
transform 1 0 1308 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5025
timestamp 1713453518
transform 1 0 1228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5026
timestamp 1713453518
transform 1 0 1108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5027
timestamp 1713453518
transform 1 0 1100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5028
timestamp 1713453518
transform 1 0 1252 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5029
timestamp 1713453518
transform 1 0 1196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1713453518
transform 1 0 2052 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1713453518
transform 1 0 1084 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5032
timestamp 1713453518
transform 1 0 3284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1713453518
transform 1 0 2012 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5034
timestamp 1713453518
transform 1 0 2036 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5035
timestamp 1713453518
transform 1 0 2028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5036
timestamp 1713453518
transform 1 0 2020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5037
timestamp 1713453518
transform 1 0 2004 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5038
timestamp 1713453518
transform 1 0 2324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5039
timestamp 1713453518
transform 1 0 2100 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1713453518
transform 1 0 2604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5041
timestamp 1713453518
transform 1 0 2532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1713453518
transform 1 0 2500 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1713453518
transform 1 0 3300 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_5044
timestamp 1713453518
transform 1 0 3236 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5045
timestamp 1713453518
transform 1 0 3108 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5046
timestamp 1713453518
transform 1 0 2596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5047
timestamp 1713453518
transform 1 0 2588 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1713453518
transform 1 0 2076 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5049
timestamp 1713453518
transform 1 0 1812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5050
timestamp 1713453518
transform 1 0 1764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5051
timestamp 1713453518
transform 1 0 1084 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5052
timestamp 1713453518
transform 1 0 3268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1713453518
transform 1 0 3268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5054
timestamp 1713453518
transform 1 0 3300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5055
timestamp 1713453518
transform 1 0 3292 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1713453518
transform 1 0 3420 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1713453518
transform 1 0 3300 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_5058
timestamp 1713453518
transform 1 0 3364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5059
timestamp 1713453518
transform 1 0 3364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5060
timestamp 1713453518
transform 1 0 1212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5061
timestamp 1713453518
transform 1 0 1180 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_5062
timestamp 1713453518
transform 1 0 1284 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1713453518
transform 1 0 1204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1713453518
transform 1 0 1132 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1713453518
transform 1 0 1140 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5066
timestamp 1713453518
transform 1 0 1100 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5067
timestamp 1713453518
transform 1 0 1100 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1713453518
transform 1 0 1092 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5069
timestamp 1713453518
transform 1 0 1076 0 1 685
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1713453518
transform 1 0 1068 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_5071
timestamp 1713453518
transform 1 0 1212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1713453518
transform 1 0 1180 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5073
timestamp 1713453518
transform 1 0 3404 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5074
timestamp 1713453518
transform 1 0 3388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1713453518
transform 1 0 3372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5076
timestamp 1713453518
transform 1 0 3372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1713453518
transform 1 0 3356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5078
timestamp 1713453518
transform 1 0 3228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5079
timestamp 1713453518
transform 1 0 3148 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5080
timestamp 1713453518
transform 1 0 3140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5081
timestamp 1713453518
transform 1 0 3132 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1713453518
transform 1 0 2260 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5083
timestamp 1713453518
transform 1 0 988 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5084
timestamp 1713453518
transform 1 0 3092 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5085
timestamp 1713453518
transform 1 0 2236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5086
timestamp 1713453518
transform 1 0 2260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5087
timestamp 1713453518
transform 1 0 2244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1713453518
transform 1 0 2268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1713453518
transform 1 0 2108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1713453518
transform 1 0 2348 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1713453518
transform 1 0 2332 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1713453518
transform 1 0 2300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5093
timestamp 1713453518
transform 1 0 2300 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5094
timestamp 1713453518
transform 1 0 2636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5095
timestamp 1713453518
transform 1 0 2548 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1713453518
transform 1 0 2420 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1713453518
transform 1 0 3204 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5098
timestamp 1713453518
transform 1 0 3060 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1713453518
transform 1 0 2940 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5100
timestamp 1713453518
transform 1 0 2476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1713453518
transform 1 0 2444 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1713453518
transform 1 0 2140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1713453518
transform 1 0 1812 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5104
timestamp 1713453518
transform 1 0 1700 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1713453518
transform 1 0 1684 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5106
timestamp 1713453518
transform 1 0 1700 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5107
timestamp 1713453518
transform 1 0 1068 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1713453518
transform 1 0 3124 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1713453518
transform 1 0 3068 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1713453518
transform 1 0 3292 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1713453518
transform 1 0 3180 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5112
timestamp 1713453518
transform 1 0 3332 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5113
timestamp 1713453518
transform 1 0 3300 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1713453518
transform 1 0 3324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5115
timestamp 1713453518
transform 1 0 3300 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5116
timestamp 1713453518
transform 1 0 1220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5117
timestamp 1713453518
transform 1 0 1196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5118
timestamp 1713453518
transform 1 0 1260 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5119
timestamp 1713453518
transform 1 0 1188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5120
timestamp 1713453518
transform 1 0 1188 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_5121
timestamp 1713453518
transform 1 0 1188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5122
timestamp 1713453518
transform 1 0 1196 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5123
timestamp 1713453518
transform 1 0 1188 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_5124
timestamp 1713453518
transform 1 0 1180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5125
timestamp 1713453518
transform 1 0 1164 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5126
timestamp 1713453518
transform 1 0 1156 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5127
timestamp 1713453518
transform 1 0 1180 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_5128
timestamp 1713453518
transform 1 0 1164 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5129
timestamp 1713453518
transform 1 0 1804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5130
timestamp 1713453518
transform 1 0 1132 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5131
timestamp 1713453518
transform 1 0 3012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5132
timestamp 1713453518
transform 1 0 1764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5133
timestamp 1713453518
transform 1 0 1796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5134
timestamp 1713453518
transform 1 0 1780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1713453518
transform 1 0 1828 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5136
timestamp 1713453518
transform 1 0 1828 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5137
timestamp 1713453518
transform 1 0 2332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5138
timestamp 1713453518
transform 1 0 1884 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5139
timestamp 1713453518
transform 1 0 2612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5140
timestamp 1713453518
transform 1 0 2276 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5141
timestamp 1713453518
transform 1 0 1772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5142
timestamp 1713453518
transform 1 0 2884 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5143
timestamp 1713453518
transform 1 0 2852 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5144
timestamp 1713453518
transform 1 0 2852 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_5145
timestamp 1713453518
transform 1 0 2412 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_5146
timestamp 1713453518
transform 1 0 1476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1713453518
transform 1 0 2204 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5148
timestamp 1713453518
transform 1 0 1668 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5149
timestamp 1713453518
transform 1 0 1636 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5150
timestamp 1713453518
transform 1 0 1636 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_5151
timestamp 1713453518
transform 1 0 2972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5152
timestamp 1713453518
transform 1 0 2956 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5153
timestamp 1713453518
transform 1 0 3092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5154
timestamp 1713453518
transform 1 0 3052 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5155
timestamp 1713453518
transform 1 0 3212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5156
timestamp 1713453518
transform 1 0 3124 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1713453518
transform 1 0 1716 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5158
timestamp 1713453518
transform 1 0 1676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5159
timestamp 1713453518
transform 1 0 1396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5160
timestamp 1713453518
transform 1 0 1372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5161
timestamp 1713453518
transform 1 0 1380 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5162
timestamp 1713453518
transform 1 0 1300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1713453518
transform 1 0 1332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5164
timestamp 1713453518
transform 1 0 1308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1713453518
transform 1 0 2212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5166
timestamp 1713453518
transform 1 0 1020 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5167
timestamp 1713453518
transform 1 0 2740 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5168
timestamp 1713453518
transform 1 0 2180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5169
timestamp 1713453518
transform 1 0 2164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5170
timestamp 1713453518
transform 1 0 2084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5171
timestamp 1713453518
transform 1 0 2300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5172
timestamp 1713453518
transform 1 0 2180 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1713453518
transform 1 0 3164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5174
timestamp 1713453518
transform 1 0 2700 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5175
timestamp 1713453518
transform 1 0 2604 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5176
timestamp 1713453518
transform 1 0 2500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5177
timestamp 1713453518
transform 1 0 2420 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5178
timestamp 1713453518
transform 1 0 2420 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5179
timestamp 1713453518
transform 1 0 2356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5180
timestamp 1713453518
transform 1 0 2348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5181
timestamp 1713453518
transform 1 0 2324 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5182
timestamp 1713453518
transform 1 0 2260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5183
timestamp 1713453518
transform 1 0 2012 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1713453518
transform 1 0 2460 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5185
timestamp 1713453518
transform 1 0 2276 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1713453518
transform 1 0 1756 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5187
timestamp 1713453518
transform 1 0 2796 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1713453518
transform 1 0 2788 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5189
timestamp 1713453518
transform 1 0 2636 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5190
timestamp 1713453518
transform 1 0 2340 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_5191
timestamp 1713453518
transform 1 0 1788 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5192
timestamp 1713453518
transform 1 0 2116 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5193
timestamp 1713453518
transform 1 0 2012 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5194
timestamp 1713453518
transform 1 0 1956 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5195
timestamp 1713453518
transform 1 0 1716 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5196
timestamp 1713453518
transform 1 0 1972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5197
timestamp 1713453518
transform 1 0 1084 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5198
timestamp 1713453518
transform 1 0 1260 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5199
timestamp 1713453518
transform 1 0 1140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1713453518
transform 1 0 1132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5201
timestamp 1713453518
transform 1 0 1084 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5202
timestamp 1713453518
transform 1 0 1196 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5203
timestamp 1713453518
transform 1 0 1140 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5204
timestamp 1713453518
transform 1 0 1132 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5205
timestamp 1713453518
transform 1 0 1116 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5206
timestamp 1713453518
transform 1 0 1668 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5207
timestamp 1713453518
transform 1 0 1596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5208
timestamp 1713453518
transform 1 0 1580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5209
timestamp 1713453518
transform 1 0 1372 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1713453518
transform 1 0 2820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5211
timestamp 1713453518
transform 1 0 2708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5212
timestamp 1713453518
transform 1 0 2724 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5213
timestamp 1713453518
transform 1 0 2708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5214
timestamp 1713453518
transform 1 0 2748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5215
timestamp 1713453518
transform 1 0 2700 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1713453518
transform 1 0 1740 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1713453518
transform 1 0 1516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1713453518
transform 1 0 1772 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5219
timestamp 1713453518
transform 1 0 1604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5220
timestamp 1713453518
transform 1 0 1540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5221
timestamp 1713453518
transform 1 0 1540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5222
timestamp 1713453518
transform 1 0 1596 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5223
timestamp 1713453518
transform 1 0 1596 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5224
timestamp 1713453518
transform 1 0 1676 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1713453518
transform 1 0 1660 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1713453518
transform 1 0 1572 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1713453518
transform 1 0 1436 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1713453518
transform 1 0 1516 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_5229
timestamp 1713453518
transform 1 0 1452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5230
timestamp 1713453518
transform 1 0 2204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1713453518
transform 1 0 1044 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5232
timestamp 1713453518
transform 1 0 2692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5233
timestamp 1713453518
transform 1 0 2180 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1713453518
transform 1 0 2188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5235
timestamp 1713453518
transform 1 0 2188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5236
timestamp 1713453518
transform 1 0 2164 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1713453518
transform 1 0 2148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5238
timestamp 1713453518
transform 1 0 2340 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1713453518
transform 1 0 2212 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1713453518
transform 1 0 3188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5241
timestamp 1713453518
transform 1 0 2740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1713453518
transform 1 0 2708 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1713453518
transform 1 0 2660 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5244
timestamp 1713453518
transform 1 0 2476 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1713453518
transform 1 0 2476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5246
timestamp 1713453518
transform 1 0 2460 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5247
timestamp 1713453518
transform 1 0 2444 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1713453518
transform 1 0 2404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1713453518
transform 1 0 2364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5250
timestamp 1713453518
transform 1 0 2324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1713453518
transform 1 0 1852 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1713453518
transform 1 0 2580 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5253
timestamp 1713453518
transform 1 0 2380 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5254
timestamp 1713453518
transform 1 0 1748 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1713453518
transform 1 0 2780 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5256
timestamp 1713453518
transform 1 0 2756 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5257
timestamp 1713453518
transform 1 0 2684 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5258
timestamp 1713453518
transform 1 0 2476 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1713453518
transform 1 0 1804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5260
timestamp 1713453518
transform 1 0 2092 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5261
timestamp 1713453518
transform 1 0 1820 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5262
timestamp 1713453518
transform 1 0 1772 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5263
timestamp 1713453518
transform 1 0 1668 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1713453518
transform 1 0 1796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5265
timestamp 1713453518
transform 1 0 1156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1713453518
transform 1 0 1628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1713453518
transform 1 0 1620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5268
timestamp 1713453518
transform 1 0 1580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1713453518
transform 1 0 1580 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5270
timestamp 1713453518
transform 1 0 1436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5271
timestamp 1713453518
transform 1 0 1428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1713453518
transform 1 0 2820 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5273
timestamp 1713453518
transform 1 0 2676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1713453518
transform 1 0 2700 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5275
timestamp 1713453518
transform 1 0 2684 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5276
timestamp 1713453518
transform 1 0 2676 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5277
timestamp 1713453518
transform 1 0 2676 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_5278
timestamp 1713453518
transform 1 0 1740 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1713453518
transform 1 0 1516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1713453518
transform 1 0 1764 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5281
timestamp 1713453518
transform 1 0 1692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5282
timestamp 1713453518
transform 1 0 1636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1713453518
transform 1 0 1596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5284
timestamp 1713453518
transform 1 0 1660 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5285
timestamp 1713453518
transform 1 0 1628 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1713453518
transform 1 0 1716 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5287
timestamp 1713453518
transform 1 0 1700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5288
timestamp 1713453518
transform 1 0 1660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1713453518
transform 1 0 1588 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1713453518
transform 1 0 1452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1713453518
transform 1 0 1356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5292
timestamp 1713453518
transform 1 0 1572 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_5293
timestamp 1713453518
transform 1 0 1460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5294
timestamp 1713453518
transform 1 0 2308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1713453518
transform 1 0 1036 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1713453518
transform 1 0 2788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5297
timestamp 1713453518
transform 1 0 2276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5298
timestamp 1713453518
transform 1 0 2284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1713453518
transform 1 0 2284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5300
timestamp 1713453518
transform 1 0 2244 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1713453518
transform 1 0 2132 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5302
timestamp 1713453518
transform 1 0 2364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5303
timestamp 1713453518
transform 1 0 2308 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5304
timestamp 1713453518
transform 1 0 3084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1713453518
transform 1 0 2564 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1713453518
transform 1 0 2548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5307
timestamp 1713453518
transform 1 0 2492 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1713453518
transform 1 0 2404 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5309
timestamp 1713453518
transform 1 0 2340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5310
timestamp 1713453518
transform 1 0 2308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5311
timestamp 1713453518
transform 1 0 2212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5312
timestamp 1713453518
transform 1 0 2204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1713453518
transform 1 0 1852 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5314
timestamp 1713453518
transform 1 0 2516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5315
timestamp 1713453518
transform 1 0 2332 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1713453518
transform 1 0 1660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5317
timestamp 1713453518
transform 1 0 2948 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5318
timestamp 1713453518
transform 1 0 2884 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5319
timestamp 1713453518
transform 1 0 2572 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5320
timestamp 1713453518
transform 1 0 2428 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_5321
timestamp 1713453518
transform 1 0 1780 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5322
timestamp 1713453518
transform 1 0 2068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5323
timestamp 1713453518
transform 1 0 1860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5324
timestamp 1713453518
transform 1 0 1812 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5325
timestamp 1713453518
transform 1 0 1652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5326
timestamp 1713453518
transform 1 0 1820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5327
timestamp 1713453518
transform 1 0 1068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5328
timestamp 1713453518
transform 1 0 1652 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5329
timestamp 1713453518
transform 1 0 1644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5330
timestamp 1713453518
transform 1 0 1604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5331
timestamp 1713453518
transform 1 0 1604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1713453518
transform 1 0 1540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5333
timestamp 1713453518
transform 1 0 1452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5334
timestamp 1713453518
transform 1 0 1452 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1713453518
transform 1 0 1380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5336
timestamp 1713453518
transform 1 0 1340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1713453518
transform 1 0 2932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5338
timestamp 1713453518
transform 1 0 2756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5339
timestamp 1713453518
transform 1 0 2772 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5340
timestamp 1713453518
transform 1 0 2756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1713453518
transform 1 0 2732 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1713453518
transform 1 0 2668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5343
timestamp 1713453518
transform 1 0 2620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5344
timestamp 1713453518
transform 1 0 2620 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1713453518
transform 1 0 1700 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1713453518
transform 1 0 1636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5347
timestamp 1713453518
transform 1 0 1764 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5348
timestamp 1713453518
transform 1 0 1676 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5349
timestamp 1713453518
transform 1 0 1628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5350
timestamp 1713453518
transform 1 0 1588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1713453518
transform 1 0 1652 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1713453518
transform 1 0 1620 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5353
timestamp 1713453518
transform 1 0 1724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5354
timestamp 1713453518
transform 1 0 1724 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5355
timestamp 1713453518
transform 1 0 1700 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5356
timestamp 1713453518
transform 1 0 1620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5357
timestamp 1713453518
transform 1 0 1588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5358
timestamp 1713453518
transform 1 0 1564 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5359
timestamp 1713453518
transform 1 0 1324 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5360
timestamp 1713453518
transform 1 0 1316 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5361
timestamp 1713453518
transform 1 0 1292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5362
timestamp 1713453518
transform 1 0 1276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5363
timestamp 1713453518
transform 1 0 1556 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_5364
timestamp 1713453518
transform 1 0 1508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1713453518
transform 1 0 1828 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1713453518
transform 1 0 988 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1713453518
transform 1 0 2932 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1713453518
transform 1 0 1804 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5369
timestamp 1713453518
transform 1 0 2004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5370
timestamp 1713453518
transform 1 0 1772 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1713453518
transform 1 0 1780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5372
timestamp 1713453518
transform 1 0 1764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5373
timestamp 1713453518
transform 1 0 1804 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5374
timestamp 1713453518
transform 1 0 1796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5375
timestamp 1713453518
transform 1 0 1772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1713453518
transform 1 0 1772 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5377
timestamp 1713453518
transform 1 0 1732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5378
timestamp 1713453518
transform 1 0 1716 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1713453518
transform 1 0 1700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5380
timestamp 1713453518
transform 1 0 1500 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_5381
timestamp 1713453518
transform 1 0 1572 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5382
timestamp 1713453518
transform 1 0 1484 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5383
timestamp 1713453518
transform 1 0 2036 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5384
timestamp 1713453518
transform 1 0 1980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5385
timestamp 1713453518
transform 1 0 1972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5386
timestamp 1713453518
transform 1 0 1964 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5387
timestamp 1713453518
transform 1 0 1892 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1713453518
transform 1 0 1644 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5389
timestamp 1713453518
transform 1 0 2180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5390
timestamp 1713453518
transform 1 0 2004 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5391
timestamp 1713453518
transform 1 0 2060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5392
timestamp 1713453518
transform 1 0 1756 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5393
timestamp 1713453518
transform 1 0 1684 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5394
timestamp 1713453518
transform 1 0 1668 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1713453518
transform 1 0 1724 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5396
timestamp 1713453518
transform 1 0 1316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5397
timestamp 1713453518
transform 1 0 3124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5398
timestamp 1713453518
transform 1 0 2852 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5399
timestamp 1713453518
transform 1 0 2844 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5400
timestamp 1713453518
transform 1 0 2772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5401
timestamp 1713453518
transform 1 0 2508 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5402
timestamp 1713453518
transform 1 0 2228 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5403
timestamp 1713453518
transform 1 0 1788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5404
timestamp 1713453518
transform 1 0 1740 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5405
timestamp 1713453518
transform 1 0 1684 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5406
timestamp 1713453518
transform 1 0 1660 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5407
timestamp 1713453518
transform 1 0 1404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1713453518
transform 1 0 1372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1713453518
transform 1 0 1372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1713453518
transform 1 0 1356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1713453518
transform 1 0 2916 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5412
timestamp 1713453518
transform 1 0 2916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5413
timestamp 1713453518
transform 1 0 3012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5414
timestamp 1713453518
transform 1 0 2972 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5415
timestamp 1713453518
transform 1 0 2596 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5416
timestamp 1713453518
transform 1 0 2508 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1713453518
transform 1 0 2380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5418
timestamp 1713453518
transform 1 0 2300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5419
timestamp 1713453518
transform 1 0 3044 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5420
timestamp 1713453518
transform 1 0 3012 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1713453518
transform 1 0 2844 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5422
timestamp 1713453518
transform 1 0 2820 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5423
timestamp 1713453518
transform 1 0 1524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5424
timestamp 1713453518
transform 1 0 2652 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5425
timestamp 1713453518
transform 1 0 2460 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1713453518
transform 1 0 2372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5427
timestamp 1713453518
transform 1 0 2316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1713453518
transform 1 0 2316 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5429
timestamp 1713453518
transform 1 0 2316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5430
timestamp 1713453518
transform 1 0 2260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5431
timestamp 1713453518
transform 1 0 2260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5432
timestamp 1713453518
transform 1 0 2452 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5433
timestamp 1713453518
transform 1 0 2428 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_5434
timestamp 1713453518
transform 1 0 2364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5435
timestamp 1713453518
transform 1 0 2356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5436
timestamp 1713453518
transform 1 0 1508 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5437
timestamp 1713453518
transform 1 0 1300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5438
timestamp 1713453518
transform 1 0 1268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5439
timestamp 1713453518
transform 1 0 1252 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_5440
timestamp 1713453518
transform 1 0 1244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5441
timestamp 1713453518
transform 1 0 1244 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1713453518
transform 1 0 1220 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_5443
timestamp 1713453518
transform 1 0 1156 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5444
timestamp 1713453518
transform 1 0 1156 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5445
timestamp 1713453518
transform 1 0 1188 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5446
timestamp 1713453518
transform 1 0 1132 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5447
timestamp 1713453518
transform 1 0 1116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5448
timestamp 1713453518
transform 1 0 1436 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1713453518
transform 1 0 1404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1713453518
transform 1 0 1716 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5451
timestamp 1713453518
transform 1 0 1636 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5452
timestamp 1713453518
transform 1 0 1492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1713453518
transform 1 0 1468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1713453518
transform 1 0 1372 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5455
timestamp 1713453518
transform 1 0 1220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1713453518
transform 1 0 2684 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1713453518
transform 1 0 2476 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5458
timestamp 1713453518
transform 1 0 2444 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1713453518
transform 1 0 2324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1713453518
transform 1 0 1868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5461
timestamp 1713453518
transform 1 0 1052 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5462
timestamp 1713453518
transform 1 0 2004 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5463
timestamp 1713453518
transform 1 0 1852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5464
timestamp 1713453518
transform 1 0 2068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1713453518
transform 1 0 1972 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5466
timestamp 1713453518
transform 1 0 2180 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1713453518
transform 1 0 1988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5468
timestamp 1713453518
transform 1 0 1996 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1713453518
transform 1 0 1940 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5470
timestamp 1713453518
transform 1 0 1836 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5471
timestamp 1713453518
transform 1 0 1716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1713453518
transform 1 0 1836 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1713453518
transform 1 0 1084 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5474
timestamp 1713453518
transform 1 0 3220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1713453518
transform 1 0 2564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5476
timestamp 1713453518
transform 1 0 2532 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1713453518
transform 1 0 2444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5478
timestamp 1713453518
transform 1 0 1980 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1713453518
transform 1 0 1812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5480
timestamp 1713453518
transform 1 0 2276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1713453518
transform 1 0 2052 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1713453518
transform 1 0 2036 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5483
timestamp 1713453518
transform 1 0 1956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1713453518
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1713453518
transform 1 0 1740 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1713453518
transform 1 0 1524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1713453518
transform 1 0 1940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1713453518
transform 1 0 1412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1713453518
transform 1 0 2484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5490
timestamp 1713453518
transform 1 0 1964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5491
timestamp 1713453518
transform 1 0 1956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5492
timestamp 1713453518
transform 1 0 1892 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5493
timestamp 1713453518
transform 1 0 1844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1713453518
transform 1 0 1404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5495
timestamp 1713453518
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5496
timestamp 1713453518
transform 1 0 1420 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5497
timestamp 1713453518
transform 1 0 1268 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1713453518
transform 1 0 1172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1713453518
transform 1 0 1148 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1713453518
transform 1 0 1220 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5501
timestamp 1713453518
transform 1 0 1204 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5502
timestamp 1713453518
transform 1 0 1156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1713453518
transform 1 0 1124 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1713453518
transform 1 0 1396 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_5505
timestamp 1713453518
transform 1 0 1348 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5506
timestamp 1713453518
transform 1 0 1428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5507
timestamp 1713453518
transform 1 0 1364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5508
timestamp 1713453518
transform 1 0 1252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1713453518
transform 1 0 1236 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5510
timestamp 1713453518
transform 1 0 1836 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1713453518
transform 1 0 1812 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5512
timestamp 1713453518
transform 1 0 1788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5513
timestamp 1713453518
transform 1 0 1756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5514
timestamp 1713453518
transform 1 0 1676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5515
timestamp 1713453518
transform 1 0 1452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5516
timestamp 1713453518
transform 1 0 1932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1713453518
transform 1 0 1092 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5518
timestamp 1713453518
transform 1 0 1948 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5519
timestamp 1713453518
transform 1 0 1908 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1713453518
transform 1 0 2132 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5521
timestamp 1713453518
transform 1 0 1916 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1713453518
transform 1 0 2172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5523
timestamp 1713453518
transform 1 0 2116 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1713453518
transform 1 0 2220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1713453518
transform 1 0 2116 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1713453518
transform 1 0 2140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1713453518
transform 1 0 2100 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1713453518
transform 1 0 2092 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1713453518
transform 1 0 1756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5530
timestamp 1713453518
transform 1 0 1716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1713453518
transform 1 0 1052 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5532
timestamp 1713453518
transform 1 0 3084 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5533
timestamp 1713453518
transform 1 0 2916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1713453518
transform 1 0 2476 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5535
timestamp 1713453518
transform 1 0 2052 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5536
timestamp 1713453518
transform 1 0 1924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5537
timestamp 1713453518
transform 1 0 2140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1713453518
transform 1 0 2124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5539
timestamp 1713453518
transform 1 0 2340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5540
timestamp 1713453518
transform 1 0 2148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5541
timestamp 1713453518
transform 1 0 3220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5542
timestamp 1713453518
transform 1 0 3220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1713453518
transform 1 0 3180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5544
timestamp 1713453518
transform 1 0 3148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5545
timestamp 1713453518
transform 1 0 3124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1713453518
transform 1 0 3108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5547
timestamp 1713453518
transform 1 0 3092 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5548
timestamp 1713453518
transform 1 0 3092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5549
timestamp 1713453518
transform 1 0 3092 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5550
timestamp 1713453518
transform 1 0 3212 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5551
timestamp 1713453518
transform 1 0 3164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5552
timestamp 1713453518
transform 1 0 2084 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1713453518
transform 1 0 1948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5554
timestamp 1713453518
transform 1 0 1932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5555
timestamp 1713453518
transform 1 0 1828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5556
timestamp 1713453518
transform 1 0 1284 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5557
timestamp 1713453518
transform 1 0 1908 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5558
timestamp 1713453518
transform 1 0 1444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5559
timestamp 1713453518
transform 1 0 1428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1713453518
transform 1 0 1428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5561
timestamp 1713453518
transform 1 0 1444 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5562
timestamp 1713453518
transform 1 0 1284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5563
timestamp 1713453518
transform 1 0 1108 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_5564
timestamp 1713453518
transform 1 0 1108 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5565
timestamp 1713453518
transform 1 0 1084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5566
timestamp 1713453518
transform 1 0 1084 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_5567
timestamp 1713453518
transform 1 0 1428 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_5568
timestamp 1713453518
transform 1 0 1372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5569
timestamp 1713453518
transform 1 0 1436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1713453518
transform 1 0 1396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5571
timestamp 1713453518
transform 1 0 1092 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5572
timestamp 1713453518
transform 1 0 1092 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5573
timestamp 1713453518
transform 1 0 1364 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5574
timestamp 1713453518
transform 1 0 1340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5575
timestamp 1713453518
transform 1 0 1332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5576
timestamp 1713453518
transform 1 0 1252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1713453518
transform 1 0 1236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5578
timestamp 1713453518
transform 1 0 1236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5579
timestamp 1713453518
transform 1 0 1196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5580
timestamp 1713453518
transform 1 0 1948 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5581
timestamp 1713453518
transform 1 0 1924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5582
timestamp 1713453518
transform 1 0 1828 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5583
timestamp 1713453518
transform 1 0 1716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5584
timestamp 1713453518
transform 1 0 3324 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5585
timestamp 1713453518
transform 1 0 3284 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5586
timestamp 1713453518
transform 1 0 1620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5587
timestamp 1713453518
transform 1 0 1460 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5588
timestamp 1713453518
transform 1 0 1860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1713453518
transform 1 0 1036 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5590
timestamp 1713453518
transform 1 0 1868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5591
timestamp 1713453518
transform 1 0 1836 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5592
timestamp 1713453518
transform 1 0 1996 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5593
timestamp 1713453518
transform 1 0 1836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5594
timestamp 1713453518
transform 1 0 2156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5595
timestamp 1713453518
transform 1 0 1956 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5596
timestamp 1713453518
transform 1 0 1972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5597
timestamp 1713453518
transform 1 0 1972 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1713453518
transform 1 0 1924 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5599
timestamp 1713453518
transform 1 0 1828 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5600
timestamp 1713453518
transform 1 0 1764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5601
timestamp 1713453518
transform 1 0 1716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5602
timestamp 1713453518
transform 1 0 1812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5603
timestamp 1713453518
transform 1 0 1020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5604
timestamp 1713453518
transform 1 0 2092 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1713453518
transform 1 0 2052 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5606
timestamp 1713453518
transform 1 0 2396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5607
timestamp 1713453518
transform 1 0 2132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5608
timestamp 1713453518
transform 1 0 3412 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5609
timestamp 1713453518
transform 1 0 3404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5610
timestamp 1713453518
transform 1 0 2052 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5611
timestamp 1713453518
transform 1 0 1884 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5612
timestamp 1713453518
transform 1 0 1868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5613
timestamp 1713453518
transform 1 0 1812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1713453518
transform 1 0 1060 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1713453518
transform 1 0 1860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5616
timestamp 1713453518
transform 1 0 1324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5617
timestamp 1713453518
transform 1 0 1316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5618
timestamp 1713453518
transform 1 0 1308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5619
timestamp 1713453518
transform 1 0 1332 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5620
timestamp 1713453518
transform 1 0 1268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5621
timestamp 1713453518
transform 1 0 1284 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5622
timestamp 1713453518
transform 1 0 1172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5623
timestamp 1713453518
transform 1 0 1156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5624
timestamp 1713453518
transform 1 0 1340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1713453518
transform 1 0 1316 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5626
timestamp 1713453518
transform 1 0 1452 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1713453518
transform 1 0 1356 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5628
timestamp 1713453518
transform 1 0 1252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5629
timestamp 1713453518
transform 1 0 1868 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5630
timestamp 1713453518
transform 1 0 1836 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5631
timestamp 1713453518
transform 1 0 3292 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1713453518
transform 1 0 3252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1713453518
transform 1 0 1748 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5634
timestamp 1713453518
transform 1 0 1684 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5635
timestamp 1713453518
transform 1 0 2084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5636
timestamp 1713453518
transform 1 0 876 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_5637
timestamp 1713453518
transform 1 0 2236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5638
timestamp 1713453518
transform 1 0 2068 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5639
timestamp 1713453518
transform 1 0 2244 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1713453518
transform 1 0 2244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1713453518
transform 1 0 2212 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5642
timestamp 1713453518
transform 1 0 1820 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5643
timestamp 1713453518
transform 1 0 2332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1713453518
transform 1 0 2220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5645
timestamp 1713453518
transform 1 0 2468 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1713453518
transform 1 0 2428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1713453518
transform 1 0 3436 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1713453518
transform 1 0 3420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5649
timestamp 1713453518
transform 1 0 1836 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5650
timestamp 1713453518
transform 1 0 1628 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1713453518
transform 1 0 1940 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1713453518
transform 1 0 1828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5653
timestamp 1713453518
transform 1 0 1596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5654
timestamp 1713453518
transform 1 0 1604 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5655
timestamp 1713453518
transform 1 0 1580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5656
timestamp 1713453518
transform 1 0 1548 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1713453518
transform 1 0 1524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1713453518
transform 1 0 2052 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1713453518
transform 1 0 2028 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1713453518
transform 1 0 1956 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5661
timestamp 1713453518
transform 1 0 1748 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1713453518
transform 1 0 3300 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5663
timestamp 1713453518
transform 1 0 3236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5664
timestamp 1713453518
transform 1 0 1740 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5665
timestamp 1713453518
transform 1 0 1724 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1713453518
transform 1 0 1740 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1713453518
transform 1 0 1732 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5668
timestamp 1713453518
transform 1 0 3332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5669
timestamp 1713453518
transform 1 0 3332 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5670
timestamp 1713453518
transform 1 0 3420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5671
timestamp 1713453518
transform 1 0 3404 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1713453518
transform 1 0 2820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5673
timestamp 1713453518
transform 1 0 2804 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1713453518
transform 1 0 1372 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_5675
timestamp 1713453518
transform 1 0 1316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1713453518
transform 1 0 932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5677
timestamp 1713453518
transform 1 0 2924 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5678
timestamp 1713453518
transform 1 0 2852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5679
timestamp 1713453518
transform 1 0 892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5680
timestamp 1713453518
transform 1 0 868 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1713453518
transform 1 0 3172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1713453518
transform 1 0 3148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5683
timestamp 1713453518
transform 1 0 3412 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5684
timestamp 1713453518
transform 1 0 3388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5685
timestamp 1713453518
transform 1 0 3180 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5686
timestamp 1713453518
transform 1 0 3156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5687
timestamp 1713453518
transform 1 0 3412 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5688
timestamp 1713453518
transform 1 0 3388 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5689
timestamp 1713453518
transform 1 0 3260 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1713453518
transform 1 0 3172 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_5691
timestamp 1713453518
transform 1 0 3188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1713453518
transform 1 0 2564 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1713453518
transform 1 0 2620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1713453518
transform 1 0 2516 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1713453518
transform 1 0 2508 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1713453518
transform 1 0 2356 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5697
timestamp 1713453518
transform 1 0 3308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5698
timestamp 1713453518
transform 1 0 3220 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5699
timestamp 1713453518
transform 1 0 3292 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1713453518
transform 1 0 3244 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5701
timestamp 1713453518
transform 1 0 3236 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5702
timestamp 1713453518
transform 1 0 3228 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_5703
timestamp 1713453518
transform 1 0 3244 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5704
timestamp 1713453518
transform 1 0 3244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5705
timestamp 1713453518
transform 1 0 2380 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5706
timestamp 1713453518
transform 1 0 2156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1713453518
transform 1 0 2156 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5708
timestamp 1713453518
transform 1 0 2124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5709
timestamp 1713453518
transform 1 0 2108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5710
timestamp 1713453518
transform 1 0 2108 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5711
timestamp 1713453518
transform 1 0 2244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1713453518
transform 1 0 2188 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5713
timestamp 1713453518
transform 1 0 2068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5714
timestamp 1713453518
transform 1 0 1972 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5715
timestamp 1713453518
transform 1 0 1876 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5716
timestamp 1713453518
transform 1 0 2196 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5717
timestamp 1713453518
transform 1 0 2148 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5718
timestamp 1713453518
transform 1 0 2156 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5719
timestamp 1713453518
transform 1 0 2124 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5720
timestamp 1713453518
transform 1 0 2052 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1713453518
transform 1 0 1980 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5722
timestamp 1713453518
transform 1 0 2108 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_5723
timestamp 1713453518
transform 1 0 2084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5724
timestamp 1713453518
transform 1 0 1948 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5725
timestamp 1713453518
transform 1 0 3140 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5726
timestamp 1713453518
transform 1 0 3028 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5727
timestamp 1713453518
transform 1 0 3044 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5728
timestamp 1713453518
transform 1 0 3012 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5729
timestamp 1713453518
transform 1 0 2860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5730
timestamp 1713453518
transform 1 0 2708 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5731
timestamp 1713453518
transform 1 0 2588 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5732
timestamp 1713453518
transform 1 0 1956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5733
timestamp 1713453518
transform 1 0 3092 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5734
timestamp 1713453518
transform 1 0 3036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5735
timestamp 1713453518
transform 1 0 2908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5736
timestamp 1713453518
transform 1 0 2724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5737
timestamp 1713453518
transform 1 0 2620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5738
timestamp 1713453518
transform 1 0 2172 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5739
timestamp 1713453518
transform 1 0 3004 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5740
timestamp 1713453518
transform 1 0 2900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5741
timestamp 1713453518
transform 1 0 2764 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5742
timestamp 1713453518
transform 1 0 2716 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5743
timestamp 1713453518
transform 1 0 2692 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5744
timestamp 1713453518
transform 1 0 2612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5745
timestamp 1713453518
transform 1 0 3132 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5746
timestamp 1713453518
transform 1 0 3084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5747
timestamp 1713453518
transform 1 0 2156 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5748
timestamp 1713453518
transform 1 0 2004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5749
timestamp 1713453518
transform 1 0 2004 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5750
timestamp 1713453518
transform 1 0 2180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5751
timestamp 1713453518
transform 1 0 2164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5752
timestamp 1713453518
transform 1 0 2044 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5753
timestamp 1713453518
transform 1 0 2036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5754
timestamp 1713453518
transform 1 0 1908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5755
timestamp 1713453518
transform 1 0 1884 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5756
timestamp 1713453518
transform 1 0 1980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1713453518
transform 1 0 1964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5758
timestamp 1713453518
transform 1 0 1892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5759
timestamp 1713453518
transform 1 0 2444 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5760
timestamp 1713453518
transform 1 0 2116 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5761
timestamp 1713453518
transform 1 0 2076 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5762
timestamp 1713453518
transform 1 0 2060 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5763
timestamp 1713453518
transform 1 0 2068 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_5764
timestamp 1713453518
transform 1 0 2028 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5765
timestamp 1713453518
transform 1 0 2028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5766
timestamp 1713453518
transform 1 0 1988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5767
timestamp 1713453518
transform 1 0 2060 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5768
timestamp 1713453518
transform 1 0 2028 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5769
timestamp 1713453518
transform 1 0 2052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5770
timestamp 1713453518
transform 1 0 2044 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5771
timestamp 1713453518
transform 1 0 2036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5772
timestamp 1713453518
transform 1 0 1972 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5773
timestamp 1713453518
transform 1 0 1940 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5774
timestamp 1713453518
transform 1 0 636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5775
timestamp 1713453518
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5776
timestamp 1713453518
transform 1 0 556 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5777
timestamp 1713453518
transform 1 0 660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5778
timestamp 1713453518
transform 1 0 612 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5779
timestamp 1713453518
transform 1 0 436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5780
timestamp 1713453518
transform 1 0 308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5781
timestamp 1713453518
transform 1 0 820 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5782
timestamp 1713453518
transform 1 0 692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5783
timestamp 1713453518
transform 1 0 444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1713453518
transform 1 0 404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5785
timestamp 1713453518
transform 1 0 636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5786
timestamp 1713453518
transform 1 0 476 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5787
timestamp 1713453518
transform 1 0 148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5788
timestamp 1713453518
transform 1 0 132 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5789
timestamp 1713453518
transform 1 0 300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1713453518
transform 1 0 260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5791
timestamp 1713453518
transform 1 0 196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5792
timestamp 1713453518
transform 1 0 156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5793
timestamp 1713453518
transform 1 0 244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5794
timestamp 1713453518
transform 1 0 236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5795
timestamp 1713453518
transform 1 0 332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5796
timestamp 1713453518
transform 1 0 292 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5797
timestamp 1713453518
transform 1 0 356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1713453518
transform 1 0 308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5799
timestamp 1713453518
transform 1 0 324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5800
timestamp 1713453518
transform 1 0 276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5801
timestamp 1713453518
transform 1 0 292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1713453518
transform 1 0 252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1713453518
transform 1 0 812 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5804
timestamp 1713453518
transform 1 0 508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5805
timestamp 1713453518
transform 1 0 756 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5806
timestamp 1713453518
transform 1 0 316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5807
timestamp 1713453518
transform 1 0 812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5808
timestamp 1713453518
transform 1 0 196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5809
timestamp 1713453518
transform 1 0 340 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5810
timestamp 1713453518
transform 1 0 284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5811
timestamp 1713453518
transform 1 0 356 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1713453518
transform 1 0 316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5813
timestamp 1713453518
transform 1 0 348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5814
timestamp 1713453518
transform 1 0 276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5815
timestamp 1713453518
transform 1 0 348 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1713453518
transform 1 0 300 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5817
timestamp 1713453518
transform 1 0 516 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5818
timestamp 1713453518
transform 1 0 460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5819
timestamp 1713453518
transform 1 0 284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5820
timestamp 1713453518
transform 1 0 244 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5821
timestamp 1713453518
transform 1 0 356 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5822
timestamp 1713453518
transform 1 0 300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5823
timestamp 1713453518
transform 1 0 412 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5824
timestamp 1713453518
transform 1 0 364 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5825
timestamp 1713453518
transform 1 0 396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5826
timestamp 1713453518
transform 1 0 356 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5827
timestamp 1713453518
transform 1 0 348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5828
timestamp 1713453518
transform 1 0 308 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5829
timestamp 1713453518
transform 1 0 724 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5830
timestamp 1713453518
transform 1 0 684 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5831
timestamp 1713453518
transform 1 0 724 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_5832
timestamp 1713453518
transform 1 0 684 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_5833
timestamp 1713453518
transform 1 0 476 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_5834
timestamp 1713453518
transform 1 0 428 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_5835
timestamp 1713453518
transform 1 0 420 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5836
timestamp 1713453518
transform 1 0 380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5837
timestamp 1713453518
transform 1 0 308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_5838
timestamp 1713453518
transform 1 0 268 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_5839
timestamp 1713453518
transform 1 0 332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5840
timestamp 1713453518
transform 1 0 284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5841
timestamp 1713453518
transform 1 0 316 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5842
timestamp 1713453518
transform 1 0 276 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1713453518
transform 1 0 716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5844
timestamp 1713453518
transform 1 0 676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5845
timestamp 1713453518
transform 1 0 252 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5846
timestamp 1713453518
transform 1 0 212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5847
timestamp 1713453518
transform 1 0 148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1713453518
transform 1 0 140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5849
timestamp 1713453518
transform 1 0 372 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5850
timestamp 1713453518
transform 1 0 300 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5851
timestamp 1713453518
transform 1 0 628 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_5852
timestamp 1713453518
transform 1 0 596 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5853
timestamp 1713453518
transform 1 0 556 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5854
timestamp 1713453518
transform 1 0 444 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5855
timestamp 1713453518
transform 1 0 444 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1713453518
transform 1 0 268 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5857
timestamp 1713453518
transform 1 0 268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5858
timestamp 1713453518
transform 1 0 252 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5859
timestamp 1713453518
transform 1 0 244 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_5860
timestamp 1713453518
transform 1 0 236 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5861
timestamp 1713453518
transform 1 0 228 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5862
timestamp 1713453518
transform 1 0 220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5863
timestamp 1713453518
transform 1 0 204 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1713453518
transform 1 0 196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5865
timestamp 1713453518
transform 1 0 572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5866
timestamp 1713453518
transform 1 0 516 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5867
timestamp 1713453518
transform 1 0 492 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5868
timestamp 1713453518
transform 1 0 476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5869
timestamp 1713453518
transform 1 0 468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5870
timestamp 1713453518
transform 1 0 388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5871
timestamp 1713453518
transform 1 0 532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5872
timestamp 1713453518
transform 1 0 340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5873
timestamp 1713453518
transform 1 0 436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5874
timestamp 1713453518
transform 1 0 396 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5875
timestamp 1713453518
transform 1 0 324 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5876
timestamp 1713453518
transform 1 0 164 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5877
timestamp 1713453518
transform 1 0 372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1713453518
transform 1 0 308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5879
timestamp 1713453518
transform 1 0 492 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5880
timestamp 1713453518
transform 1 0 396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1713453518
transform 1 0 372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5882
timestamp 1713453518
transform 1 0 332 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1713453518
transform 1 0 332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1713453518
transform 1 0 164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1713453518
transform 1 0 148 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5886
timestamp 1713453518
transform 1 0 108 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1713453518
transform 1 0 364 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5888
timestamp 1713453518
transform 1 0 132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5889
timestamp 1713453518
transform 1 0 588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5890
timestamp 1713453518
transform 1 0 356 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_5891
timestamp 1713453518
transform 1 0 572 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5892
timestamp 1713453518
transform 1 0 556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5893
timestamp 1713453518
transform 1 0 556 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5894
timestamp 1713453518
transform 1 0 548 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_5895
timestamp 1713453518
transform 1 0 532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5896
timestamp 1713453518
transform 1 0 492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5897
timestamp 1713453518
transform 1 0 484 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5898
timestamp 1713453518
transform 1 0 476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5899
timestamp 1713453518
transform 1 0 572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5900
timestamp 1713453518
transform 1 0 572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1713453518
transform 1 0 588 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5902
timestamp 1713453518
transform 1 0 564 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5903
timestamp 1713453518
transform 1 0 548 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5904
timestamp 1713453518
transform 1 0 468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5905
timestamp 1713453518
transform 1 0 252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5906
timestamp 1713453518
transform 1 0 252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5907
timestamp 1713453518
transform 1 0 236 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5908
timestamp 1713453518
transform 1 0 220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5909
timestamp 1713453518
transform 1 0 444 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5910
timestamp 1713453518
transform 1 0 236 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5911
timestamp 1713453518
transform 1 0 556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5912
timestamp 1713453518
transform 1 0 452 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1713453518
transform 1 0 540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5914
timestamp 1713453518
transform 1 0 540 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5915
timestamp 1713453518
transform 1 0 364 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1713453518
transform 1 0 300 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5917
timestamp 1713453518
transform 1 0 380 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5918
timestamp 1713453518
transform 1 0 340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5919
timestamp 1713453518
transform 1 0 500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5920
timestamp 1713453518
transform 1 0 492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5921
timestamp 1713453518
transform 1 0 484 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5922
timestamp 1713453518
transform 1 0 460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5923
timestamp 1713453518
transform 1 0 444 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5924
timestamp 1713453518
transform 1 0 572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1713453518
transform 1 0 540 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5926
timestamp 1713453518
transform 1 0 540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1713453518
transform 1 0 652 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5928
timestamp 1713453518
transform 1 0 612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5929
timestamp 1713453518
transform 1 0 596 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1713453518
transform 1 0 588 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_5931
timestamp 1713453518
transform 1 0 588 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5932
timestamp 1713453518
transform 1 0 580 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5933
timestamp 1713453518
transform 1 0 428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5934
timestamp 1713453518
transform 1 0 236 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5935
timestamp 1713453518
transform 1 0 676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5936
timestamp 1713453518
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1713453518
transform 1 0 652 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5938
timestamp 1713453518
transform 1 0 644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5939
timestamp 1713453518
transform 1 0 628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5940
timestamp 1713453518
transform 1 0 588 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5941
timestamp 1713453518
transform 1 0 556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5942
timestamp 1713453518
transform 1 0 556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5943
timestamp 1713453518
transform 1 0 676 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5944
timestamp 1713453518
transform 1 0 604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1713453518
transform 1 0 628 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5946
timestamp 1713453518
transform 1 0 620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5947
timestamp 1713453518
transform 1 0 596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1713453518
transform 1 0 540 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5949
timestamp 1713453518
transform 1 0 540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5950
timestamp 1713453518
transform 1 0 460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5951
timestamp 1713453518
transform 1 0 260 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5952
timestamp 1713453518
transform 1 0 636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5953
timestamp 1713453518
transform 1 0 452 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5954
timestamp 1713453518
transform 1 0 635 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1713453518
transform 1 0 556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5956
timestamp 1713453518
transform 1 0 420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5957
timestamp 1713453518
transform 1 0 236 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5958
timestamp 1713453518
transform 1 0 580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5959
timestamp 1713453518
transform 1 0 412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5960
timestamp 1713453518
transform 1 0 580 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5961
timestamp 1713453518
transform 1 0 548 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5962
timestamp 1713453518
transform 1 0 404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5963
timestamp 1713453518
transform 1 0 180 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5964
timestamp 1713453518
transform 1 0 676 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5965
timestamp 1713453518
transform 1 0 396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1713453518
transform 1 0 684 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5967
timestamp 1713453518
transform 1 0 644 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5968
timestamp 1713453518
transform 1 0 652 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5969
timestamp 1713453518
transform 1 0 588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5970
timestamp 1713453518
transform 1 0 564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5971
timestamp 1713453518
transform 1 0 548 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5972
timestamp 1713453518
transform 1 0 596 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5973
timestamp 1713453518
transform 1 0 596 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5974
timestamp 1713453518
transform 1 0 588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5975
timestamp 1713453518
transform 1 0 628 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5976
timestamp 1713453518
transform 1 0 612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5977
timestamp 1713453518
transform 1 0 516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5978
timestamp 1713453518
transform 1 0 516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5979
timestamp 1713453518
transform 1 0 452 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5980
timestamp 1713453518
transform 1 0 716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5981
timestamp 1713453518
transform 1 0 628 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5982
timestamp 1713453518
transform 1 0 620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5983
timestamp 1713453518
transform 1 0 620 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5984
timestamp 1713453518
transform 1 0 572 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1713453518
transform 1 0 420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5986
timestamp 1713453518
transform 1 0 396 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5987
timestamp 1713453518
transform 1 0 604 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5988
timestamp 1713453518
transform 1 0 412 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5989
timestamp 1713453518
transform 1 0 628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5990
timestamp 1713453518
transform 1 0 604 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1713453518
transform 1 0 700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5992
timestamp 1713453518
transform 1 0 684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5993
timestamp 1713453518
transform 1 0 652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5994
timestamp 1713453518
transform 1 0 644 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5995
timestamp 1713453518
transform 1 0 620 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5996
timestamp 1713453518
transform 1 0 612 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5997
timestamp 1713453518
transform 1 0 388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1713453518
transform 1 0 364 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5999
timestamp 1713453518
transform 1 0 740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6000
timestamp 1713453518
transform 1 0 380 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6001
timestamp 1713453518
transform 1 0 740 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6002
timestamp 1713453518
transform 1 0 692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6003
timestamp 1713453518
transform 1 0 348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6004
timestamp 1713453518
transform 1 0 252 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6005
timestamp 1713453518
transform 1 0 644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6006
timestamp 1713453518
transform 1 0 340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6007
timestamp 1713453518
transform 1 0 668 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6008
timestamp 1713453518
transform 1 0 644 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6009
timestamp 1713453518
transform 1 0 436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6010
timestamp 1713453518
transform 1 0 252 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_6011
timestamp 1713453518
transform 1 0 692 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6012
timestamp 1713453518
transform 1 0 412 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6013
timestamp 1713453518
transform 1 0 716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6014
timestamp 1713453518
transform 1 0 692 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6015
timestamp 1713453518
transform 1 0 724 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6016
timestamp 1713453518
transform 1 0 540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6017
timestamp 1713453518
transform 1 0 540 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6018
timestamp 1713453518
transform 1 0 492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6019
timestamp 1713453518
transform 1 0 780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6020
timestamp 1713453518
transform 1 0 740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6021
timestamp 1713453518
transform 1 0 676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6022
timestamp 1713453518
transform 1 0 588 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6023
timestamp 1713453518
transform 1 0 588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6024
timestamp 1713453518
transform 1 0 588 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_6025
timestamp 1713453518
transform 1 0 748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6026
timestamp 1713453518
transform 1 0 684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6027
timestamp 1713453518
transform 1 0 652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6028
timestamp 1713453518
transform 1 0 636 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6029
timestamp 1713453518
transform 1 0 628 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_6030
timestamp 1713453518
transform 1 0 572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6031
timestamp 1713453518
transform 1 0 460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6032
timestamp 1713453518
transform 1 0 260 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1713453518
transform 1 0 596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6034
timestamp 1713453518
transform 1 0 452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6035
timestamp 1713453518
transform 1 0 724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6036
timestamp 1713453518
transform 1 0 644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6037
timestamp 1713453518
transform 1 0 644 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1713453518
transform 1 0 644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6039
timestamp 1713453518
transform 1 0 604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6040
timestamp 1713453518
transform 1 0 572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1713453518
transform 1 0 596 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1713453518
transform 1 0 580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6043
timestamp 1713453518
transform 1 0 460 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6044
timestamp 1713453518
transform 1 0 260 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_6045
timestamp 1713453518
transform 1 0 700 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6046
timestamp 1713453518
transform 1 0 452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6047
timestamp 1713453518
transform 1 0 692 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_6048
timestamp 1713453518
transform 1 0 668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6049
timestamp 1713453518
transform 1 0 460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6050
timestamp 1713453518
transform 1 0 252 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_6051
timestamp 1713453518
transform 1 0 748 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6052
timestamp 1713453518
transform 1 0 452 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6053
timestamp 1713453518
transform 1 0 748 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_6054
timestamp 1713453518
transform 1 0 732 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6055
timestamp 1713453518
transform 1 0 500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6056
timestamp 1713453518
transform 1 0 420 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6057
timestamp 1713453518
transform 1 0 716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6058
timestamp 1713453518
transform 1 0 492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6059
timestamp 1713453518
transform 1 0 772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6060
timestamp 1713453518
transform 1 0 724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1713453518
transform 1 0 620 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_6062
timestamp 1713453518
transform 1 0 596 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6063
timestamp 1713453518
transform 1 0 572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6064
timestamp 1713453518
transform 1 0 788 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_6065
timestamp 1713453518
transform 1 0 604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6066
timestamp 1713453518
transform 1 0 524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6067
timestamp 1713453518
transform 1 0 500 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6068
timestamp 1713453518
transform 1 0 476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6069
timestamp 1713453518
transform 1 0 452 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1713453518
transform 1 0 452 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6071
timestamp 1713453518
transform 1 0 796 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6072
timestamp 1713453518
transform 1 0 788 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6073
timestamp 1713453518
transform 1 0 692 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6074
timestamp 1713453518
transform 1 0 692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6075
timestamp 1713453518
transform 1 0 684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6076
timestamp 1713453518
transform 1 0 636 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6077
timestamp 1713453518
transform 1 0 628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6078
timestamp 1713453518
transform 1 0 596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6079
timestamp 1713453518
transform 1 0 252 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1713453518
transform 1 0 604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1713453518
transform 1 0 588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6082
timestamp 1713453518
transform 1 0 628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6083
timestamp 1713453518
transform 1 0 604 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_6084
timestamp 1713453518
transform 1 0 780 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6085
timestamp 1713453518
transform 1 0 748 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6086
timestamp 1713453518
transform 1 0 676 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6087
timestamp 1713453518
transform 1 0 676 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6088
timestamp 1713453518
transform 1 0 612 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6089
timestamp 1713453518
transform 1 0 612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6090
timestamp 1713453518
transform 1 0 412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1713453518
transform 1 0 244 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6092
timestamp 1713453518
transform 1 0 660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6093
timestamp 1713453518
transform 1 0 396 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6094
timestamp 1713453518
transform 1 0 684 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6095
timestamp 1713453518
transform 1 0 660 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6096
timestamp 1713453518
transform 1 0 444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6097
timestamp 1713453518
transform 1 0 300 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6098
timestamp 1713453518
transform 1 0 772 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6099
timestamp 1713453518
transform 1 0 436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6100
timestamp 1713453518
transform 1 0 788 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6101
timestamp 1713453518
transform 1 0 764 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1713453518
transform 1 0 500 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6103
timestamp 1713453518
transform 1 0 292 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1713453518
transform 1 0 740 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6105
timestamp 1713453518
transform 1 0 492 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6106
timestamp 1713453518
transform 1 0 772 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6107
timestamp 1713453518
transform 1 0 740 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6108
timestamp 1713453518
transform 1 0 668 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6109
timestamp 1713453518
transform 1 0 652 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1713453518
transform 1 0 620 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6111
timestamp 1713453518
transform 1 0 604 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6112
timestamp 1713453518
transform 1 0 580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6113
timestamp 1713453518
transform 1 0 716 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_6114
timestamp 1713453518
transform 1 0 644 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6115
timestamp 1713453518
transform 1 0 524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6116
timestamp 1713453518
transform 1 0 508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6117
timestamp 1713453518
transform 1 0 508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6118
timestamp 1713453518
transform 1 0 508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6119
timestamp 1713453518
transform 1 0 676 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6120
timestamp 1713453518
transform 1 0 636 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1713453518
transform 1 0 812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6122
timestamp 1713453518
transform 1 0 804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6123
timestamp 1713453518
transform 1 0 780 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6124
timestamp 1713453518
transform 1 0 772 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6125
timestamp 1713453518
transform 1 0 692 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6126
timestamp 1713453518
transform 1 0 596 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6127
timestamp 1713453518
transform 1 0 564 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6128
timestamp 1713453518
transform 1 0 460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6129
timestamp 1713453518
transform 1 0 252 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6130
timestamp 1713453518
transform 1 0 716 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6131
timestamp 1713453518
transform 1 0 452 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1713453518
transform 1 0 716 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6133
timestamp 1713453518
transform 1 0 668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6134
timestamp 1713453518
transform 1 0 732 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6135
timestamp 1713453518
transform 1 0 732 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6136
timestamp 1713453518
transform 1 0 660 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6137
timestamp 1713453518
transform 1 0 636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6138
timestamp 1713453518
transform 1 0 628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6139
timestamp 1713453518
transform 1 0 620 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6140
timestamp 1713453518
transform 1 0 660 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1713453518
transform 1 0 636 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6142
timestamp 1713453518
transform 1 0 820 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6143
timestamp 1713453518
transform 1 0 652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6144
timestamp 1713453518
transform 1 0 804 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6145
timestamp 1713453518
transform 1 0 756 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6146
timestamp 1713453518
transform 1 0 660 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6147
timestamp 1713453518
transform 1 0 652 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6148
timestamp 1713453518
transform 1 0 836 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_6149
timestamp 1713453518
transform 1 0 628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6150
timestamp 1713453518
transform 1 0 836 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6151
timestamp 1713453518
transform 1 0 756 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6152
timestamp 1713453518
transform 1 0 540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1713453518
transform 1 0 508 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6154
timestamp 1713453518
transform 1 0 860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6155
timestamp 1713453518
transform 1 0 508 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6156
timestamp 1713453518
transform 1 0 868 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6157
timestamp 1713453518
transform 1 0 692 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6158
timestamp 1713453518
transform 1 0 636 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6159
timestamp 1713453518
transform 1 0 612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6160
timestamp 1713453518
transform 1 0 564 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6161
timestamp 1713453518
transform 1 0 548 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6162
timestamp 1713453518
transform 1 0 708 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6163
timestamp 1713453518
transform 1 0 660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6164
timestamp 1713453518
transform 1 0 596 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6165
timestamp 1713453518
transform 1 0 588 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6166
timestamp 1713453518
transform 1 0 532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6167
timestamp 1713453518
transform 1 0 532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6168
timestamp 1713453518
transform 1 0 740 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6169
timestamp 1713453518
transform 1 0 556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6170
timestamp 1713453518
transform 1 0 516 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1713453518
transform 1 0 516 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6172
timestamp 1713453518
transform 1 0 500 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6173
timestamp 1713453518
transform 1 0 668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6174
timestamp 1713453518
transform 1 0 604 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1713453518
transform 1 0 564 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6176
timestamp 1713453518
transform 1 0 540 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6177
timestamp 1713453518
transform 1 0 540 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6178
timestamp 1713453518
transform 1 0 500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6179
timestamp 1713453518
transform 1 0 420 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6180
timestamp 1713453518
transform 1 0 276 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6181
timestamp 1713453518
transform 1 0 556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6182
timestamp 1713453518
transform 1 0 412 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6183
timestamp 1713453518
transform 1 0 620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6184
timestamp 1713453518
transform 1 0 596 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6185
timestamp 1713453518
transform 1 0 564 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6186
timestamp 1713453518
transform 1 0 564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6187
timestamp 1713453518
transform 1 0 532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6188
timestamp 1713453518
transform 1 0 556 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6189
timestamp 1713453518
transform 1 0 516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6190
timestamp 1713453518
transform 1 0 540 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6191
timestamp 1713453518
transform 1 0 228 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_6192
timestamp 1713453518
transform 1 0 644 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6193
timestamp 1713453518
transform 1 0 532 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6194
timestamp 1713453518
transform 1 0 692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6195
timestamp 1713453518
transform 1 0 676 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6196
timestamp 1713453518
transform 1 0 468 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6197
timestamp 1713453518
transform 1 0 220 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6198
timestamp 1713453518
transform 1 0 604 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6199
timestamp 1713453518
transform 1 0 460 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6200
timestamp 1713453518
transform 1 0 644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6201
timestamp 1713453518
transform 1 0 628 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6202
timestamp 1713453518
transform 1 0 476 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6203
timestamp 1713453518
transform 1 0 236 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6204
timestamp 1713453518
transform 1 0 588 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6205
timestamp 1713453518
transform 1 0 468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6206
timestamp 1713453518
transform 1 0 588 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6207
timestamp 1713453518
transform 1 0 572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6208
timestamp 1713453518
transform 1 0 692 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6209
timestamp 1713453518
transform 1 0 596 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6210
timestamp 1713453518
transform 1 0 580 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6211
timestamp 1713453518
transform 1 0 532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6212
timestamp 1713453518
transform 1 0 524 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6213
timestamp 1713453518
transform 1 0 508 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6214
timestamp 1713453518
transform 1 0 772 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6215
timestamp 1713453518
transform 1 0 588 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6216
timestamp 1713453518
transform 1 0 524 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6217
timestamp 1713453518
transform 1 0 524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6218
timestamp 1713453518
transform 1 0 492 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6219
timestamp 1713453518
transform 1 0 484 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6220
timestamp 1713453518
transform 1 0 468 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6221
timestamp 1713453518
transform 1 0 532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6222
timestamp 1713453518
transform 1 0 524 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_6223
timestamp 1713453518
transform 1 0 500 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_6224
timestamp 1713453518
transform 1 0 484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6225
timestamp 1713453518
transform 1 0 476 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_6226
timestamp 1713453518
transform 1 0 476 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6227
timestamp 1713453518
transform 1 0 460 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6228
timestamp 1713453518
transform 1 0 444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6229
timestamp 1713453518
transform 1 0 532 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6230
timestamp 1713453518
transform 1 0 500 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6231
timestamp 1713453518
transform 1 0 412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6232
timestamp 1713453518
transform 1 0 412 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6233
timestamp 1713453518
transform 1 0 508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6234
timestamp 1713453518
transform 1 0 508 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6235
timestamp 1713453518
transform 1 0 604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6236
timestamp 1713453518
transform 1 0 540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6237
timestamp 1713453518
transform 1 0 572 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1713453518
transform 1 0 564 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_6239
timestamp 1713453518
transform 1 0 596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_6240
timestamp 1713453518
transform 1 0 564 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_6241
timestamp 1713453518
transform 1 0 596 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_6242
timestamp 1713453518
transform 1 0 588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6243
timestamp 1713453518
transform 1 0 580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_6244
timestamp 1713453518
transform 1 0 676 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6245
timestamp 1713453518
transform 1 0 596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6246
timestamp 1713453518
transform 1 0 612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6247
timestamp 1713453518
transform 1 0 524 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_6248
timestamp 1713453518
transform 1 0 532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6249
timestamp 1713453518
transform 1 0 484 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_6250
timestamp 1713453518
transform 1 0 492 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_6251
timestamp 1713453518
transform 1 0 404 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6252
timestamp 1713453518
transform 1 0 476 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6253
timestamp 1713453518
transform 1 0 380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_6254
timestamp 1713453518
transform 1 0 356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6255
timestamp 1713453518
transform 1 0 420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6256
timestamp 1713453518
transform 1 0 380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6257
timestamp 1713453518
transform 1 0 468 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6258
timestamp 1713453518
transform 1 0 452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6259
timestamp 1713453518
transform 1 0 516 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6260
timestamp 1713453518
transform 1 0 460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6261
timestamp 1713453518
transform 1 0 476 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6262
timestamp 1713453518
transform 1 0 468 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6263
timestamp 1713453518
transform 1 0 428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_6264
timestamp 1713453518
transform 1 0 548 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6265
timestamp 1713453518
transform 1 0 532 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6266
timestamp 1713453518
transform 1 0 460 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1713453518
transform 1 0 468 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6268
timestamp 1713453518
transform 1 0 460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6269
timestamp 1713453518
transform 1 0 508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6270
timestamp 1713453518
transform 1 0 436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6271
timestamp 1713453518
transform 1 0 660 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_6272
timestamp 1713453518
transform 1 0 540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6273
timestamp 1713453518
transform 1 0 484 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_6274
timestamp 1713453518
transform 1 0 676 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6275
timestamp 1713453518
transform 1 0 676 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6276
timestamp 1713453518
transform 1 0 668 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6277
timestamp 1713453518
transform 1 0 580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1713453518
transform 1 0 492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6279
timestamp 1713453518
transform 1 0 484 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6280
timestamp 1713453518
transform 1 0 452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6281
timestamp 1713453518
transform 1 0 316 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6282
timestamp 1713453518
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6283
timestamp 1713453518
transform 1 0 268 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6284
timestamp 1713453518
transform 1 0 260 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6285
timestamp 1713453518
transform 1 0 260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6286
timestamp 1713453518
transform 1 0 260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6287
timestamp 1713453518
transform 1 0 244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6288
timestamp 1713453518
transform 1 0 244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6289
timestamp 1713453518
transform 1 0 236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6290
timestamp 1713453518
transform 1 0 668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1713453518
transform 1 0 652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6292
timestamp 1713453518
transform 1 0 596 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_6293
timestamp 1713453518
transform 1 0 580 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_6294
timestamp 1713453518
transform 1 0 556 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_6295
timestamp 1713453518
transform 1 0 564 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_6296
timestamp 1713453518
transform 1 0 532 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_6297
timestamp 1713453518
transform 1 0 500 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_6298
timestamp 1713453518
transform 1 0 668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6299
timestamp 1713453518
transform 1 0 652 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_6300
timestamp 1713453518
transform 1 0 444 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_6301
timestamp 1713453518
transform 1 0 436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6302
timestamp 1713453518
transform 1 0 804 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6303
timestamp 1713453518
transform 1 0 764 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1713453518
transform 1 0 692 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1713453518
transform 1 0 684 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6306
timestamp 1713453518
transform 1 0 732 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6307
timestamp 1713453518
transform 1 0 716 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_6308
timestamp 1713453518
transform 1 0 708 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_6309
timestamp 1713453518
transform 1 0 708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6310
timestamp 1713453518
transform 1 0 724 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6311
timestamp 1713453518
transform 1 0 708 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_6312
timestamp 1713453518
transform 1 0 644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_6313
timestamp 1713453518
transform 1 0 604 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_6314
timestamp 1713453518
transform 1 0 348 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_6315
timestamp 1713453518
transform 1 0 340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6316
timestamp 1713453518
transform 1 0 324 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6317
timestamp 1713453518
transform 1 0 212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6318
timestamp 1713453518
transform 1 0 452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_6319
timestamp 1713453518
transform 1 0 356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6320
timestamp 1713453518
transform 1 0 164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6321
timestamp 1713453518
transform 1 0 140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1713453518
transform 1 0 124 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1713453518
transform 1 0 124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6324
timestamp 1713453518
transform 1 0 228 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1713453518
transform 1 0 156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1713453518
transform 1 0 276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6327
timestamp 1713453518
transform 1 0 260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6328
timestamp 1713453518
transform 1 0 236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6329
timestamp 1713453518
transform 1 0 116 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1713453518
transform 1 0 260 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1713453518
transform 1 0 148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6332
timestamp 1713453518
transform 1 0 236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6333
timestamp 1713453518
transform 1 0 116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6334
timestamp 1713453518
transform 1 0 172 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1713453518
transform 1 0 116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6336
timestamp 1713453518
transform 1 0 372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6337
timestamp 1713453518
transform 1 0 260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6338
timestamp 1713453518
transform 1 0 356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1713453518
transform 1 0 252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6340
timestamp 1713453518
transform 1 0 252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6341
timestamp 1713453518
transform 1 0 148 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6342
timestamp 1713453518
transform 1 0 252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6343
timestamp 1713453518
transform 1 0 140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6344
timestamp 1713453518
transform 1 0 260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6345
timestamp 1713453518
transform 1 0 148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6346
timestamp 1713453518
transform 1 0 260 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6347
timestamp 1713453518
transform 1 0 148 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6348
timestamp 1713453518
transform 1 0 252 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6349
timestamp 1713453518
transform 1 0 116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6350
timestamp 1713453518
transform 1 0 420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6351
timestamp 1713453518
transform 1 0 316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6352
timestamp 1713453518
transform 1 0 244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6353
timestamp 1713453518
transform 1 0 140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6354
timestamp 1713453518
transform 1 0 244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6355
timestamp 1713453518
transform 1 0 140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6356
timestamp 1713453518
transform 1 0 300 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6357
timestamp 1713453518
transform 1 0 148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6358
timestamp 1713453518
transform 1 0 292 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6359
timestamp 1713453518
transform 1 0 164 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6360
timestamp 1713453518
transform 1 0 252 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1713453518
transform 1 0 132 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6362
timestamp 1713453518
transform 1 0 620 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6363
timestamp 1713453518
transform 1 0 572 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1713453518
transform 1 0 660 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6365
timestamp 1713453518
transform 1 0 564 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6366
timestamp 1713453518
transform 1 0 468 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6367
timestamp 1713453518
transform 1 0 356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6368
timestamp 1713453518
transform 1 0 276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6369
timestamp 1713453518
transform 1 0 228 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6370
timestamp 1713453518
transform 1 0 228 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_6371
timestamp 1713453518
transform 1 0 132 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6372
timestamp 1713453518
transform 1 0 220 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6373
timestamp 1713453518
transform 1 0 132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6374
timestamp 1713453518
transform 1 0 236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6375
timestamp 1713453518
transform 1 0 132 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6376
timestamp 1713453518
transform 1 0 572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6377
timestamp 1713453518
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6378
timestamp 1713453518
transform 1 0 1244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6379
timestamp 1713453518
transform 1 0 1004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1713453518
transform 1 0 1140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6381
timestamp 1713453518
transform 1 0 1100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6382
timestamp 1713453518
transform 1 0 1132 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6383
timestamp 1713453518
transform 1 0 1092 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6384
timestamp 1713453518
transform 1 0 1260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6385
timestamp 1713453518
transform 1 0 1220 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1713453518
transform 1 0 1292 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1713453518
transform 1 0 1260 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_6388
timestamp 1713453518
transform 1 0 492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_6389
timestamp 1713453518
transform 1 0 492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6390
timestamp 1713453518
transform 1 0 876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6391
timestamp 1713453518
transform 1 0 844 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6392
timestamp 1713453518
transform 1 0 732 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_6393
timestamp 1713453518
transform 1 0 572 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6394
timestamp 1713453518
transform 1 0 420 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6395
timestamp 1713453518
transform 1 0 220 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1713453518
transform 1 0 460 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6397
timestamp 1713453518
transform 1 0 204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6398
timestamp 1713453518
transform 1 0 404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1713453518
transform 1 0 372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6400
timestamp 1713453518
transform 1 0 764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6401
timestamp 1713453518
transform 1 0 700 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_6402
timestamp 1713453518
transform 1 0 748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6403
timestamp 1713453518
transform 1 0 724 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_6404
timestamp 1713453518
transform 1 0 884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6405
timestamp 1713453518
transform 1 0 852 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_6406
timestamp 1713453518
transform 1 0 868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6407
timestamp 1713453518
transform 1 0 852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6408
timestamp 1713453518
transform 1 0 684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6409
timestamp 1713453518
transform 1 0 524 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6410
timestamp 1713453518
transform 1 0 804 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_6411
timestamp 1713453518
transform 1 0 724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6412
timestamp 1713453518
transform 1 0 844 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6413
timestamp 1713453518
transform 1 0 836 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_6414
timestamp 1713453518
transform 1 0 1604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6415
timestamp 1713453518
transform 1 0 1580 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6416
timestamp 1713453518
transform 1 0 1436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6417
timestamp 1713453518
transform 1 0 1420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_6418
timestamp 1713453518
transform 1 0 1412 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6419
timestamp 1713453518
transform 1 0 620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6420
timestamp 1713453518
transform 1 0 412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6421
timestamp 1713453518
transform 1 0 260 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6422
timestamp 1713453518
transform 1 0 1620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6423
timestamp 1713453518
transform 1 0 1548 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_6424
timestamp 1713453518
transform 1 0 1524 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6425
timestamp 1713453518
transform 1 0 1516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_6426
timestamp 1713453518
transform 1 0 1500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_6427
timestamp 1713453518
transform 1 0 1900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6428
timestamp 1713453518
transform 1 0 1836 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_6429
timestamp 1713453518
transform 1 0 1812 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6430
timestamp 1713453518
transform 1 0 1516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6431
timestamp 1713453518
transform 1 0 1420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6432
timestamp 1713453518
transform 1 0 1516 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6433
timestamp 1713453518
transform 1 0 1500 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6434
timestamp 1713453518
transform 1 0 1548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6435
timestamp 1713453518
transform 1 0 1516 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6436
timestamp 1713453518
transform 1 0 1556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6437
timestamp 1713453518
transform 1 0 1468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1713453518
transform 1 0 1428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6439
timestamp 1713453518
transform 1 0 1380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6440
timestamp 1713453518
transform 1 0 1532 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6441
timestamp 1713453518
transform 1 0 1492 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6442
timestamp 1713453518
transform 1 0 1468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6443
timestamp 1713453518
transform 1 0 1444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6444
timestamp 1713453518
transform 1 0 1388 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6445
timestamp 1713453518
transform 1 0 1420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6446
timestamp 1713453518
transform 1 0 1420 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6447
timestamp 1713453518
transform 1 0 1388 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6448
timestamp 1713453518
transform 1 0 1436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1713453518
transform 1 0 1396 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6450
timestamp 1713453518
transform 1 0 1372 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_6451
timestamp 1713453518
transform 1 0 1348 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_6452
timestamp 1713453518
transform 1 0 1340 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6453
timestamp 1713453518
transform 1 0 1492 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_6454
timestamp 1713453518
transform 1 0 1380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6455
timestamp 1713453518
transform 1 0 1412 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_6456
timestamp 1713453518
transform 1 0 1356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6457
timestamp 1713453518
transform 1 0 3044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6458
timestamp 1713453518
transform 1 0 2972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1713453518
transform 1 0 2604 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6460
timestamp 1713453518
transform 1 0 2404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6461
timestamp 1713453518
transform 1 0 2228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6462
timestamp 1713453518
transform 1 0 1644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6463
timestamp 1713453518
transform 1 0 1284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6464
timestamp 1713453518
transform 1 0 972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6465
timestamp 1713453518
transform 1 0 1316 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_6466
timestamp 1713453518
transform 1 0 1044 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_6467
timestamp 1713453518
transform 1 0 1708 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_6468
timestamp 1713453518
transform 1 0 1572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6469
timestamp 1713453518
transform 1 0 1580 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_6470
timestamp 1713453518
transform 1 0 948 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6471
timestamp 1713453518
transform 1 0 772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6472
timestamp 1713453518
transform 1 0 724 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6473
timestamp 1713453518
transform 1 0 652 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6474
timestamp 1713453518
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6475
timestamp 1713453518
transform 1 0 860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6476
timestamp 1713453518
transform 1 0 836 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6477
timestamp 1713453518
transform 1 0 836 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6478
timestamp 1713453518
transform 1 0 820 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6479
timestamp 1713453518
transform 1 0 820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6480
timestamp 1713453518
transform 1 0 812 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6481
timestamp 1713453518
transform 1 0 780 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6482
timestamp 1713453518
transform 1 0 756 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1713453518
transform 1 0 756 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_6484
timestamp 1713453518
transform 1 0 1412 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_6485
timestamp 1713453518
transform 1 0 1076 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6486
timestamp 1713453518
transform 1 0 756 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6487
timestamp 1713453518
transform 1 0 692 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_6488
timestamp 1713453518
transform 1 0 652 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6489
timestamp 1713453518
transform 1 0 628 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6490
timestamp 1713453518
transform 1 0 1372 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_6491
timestamp 1713453518
transform 1 0 996 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6492
timestamp 1713453518
transform 1 0 804 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_6493
timestamp 1713453518
transform 1 0 780 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6494
timestamp 1713453518
transform 1 0 676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6495
timestamp 1713453518
transform 1 0 652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6496
timestamp 1713453518
transform 1 0 1300 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_6497
timestamp 1713453518
transform 1 0 988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6498
timestamp 1713453518
transform 1 0 748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1713453518
transform 1 0 716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6500
timestamp 1713453518
transform 1 0 636 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_6501
timestamp 1713453518
transform 1 0 628 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6502
timestamp 1713453518
transform 1 0 1276 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_6503
timestamp 1713453518
transform 1 0 996 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6504
timestamp 1713453518
transform 1 0 932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6505
timestamp 1713453518
transform 1 0 740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6506
timestamp 1713453518
transform 1 0 724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6507
timestamp 1713453518
transform 1 0 940 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6508
timestamp 1713453518
transform 1 0 788 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6509
timestamp 1713453518
transform 1 0 772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6510
timestamp 1713453518
transform 1 0 580 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6511
timestamp 1713453518
transform 1 0 1476 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_6512
timestamp 1713453518
transform 1 0 1004 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6513
timestamp 1713453518
transform 1 0 788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6514
timestamp 1713453518
transform 1 0 724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6515
timestamp 1713453518
transform 1 0 724 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_6516
timestamp 1713453518
transform 1 0 684 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6517
timestamp 1713453518
transform 1 0 460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6518
timestamp 1713453518
transform 1 0 444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6519
timestamp 1713453518
transform 1 0 900 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6520
timestamp 1713453518
transform 1 0 748 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6521
timestamp 1713453518
transform 1 0 724 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6522
timestamp 1713453518
transform 1 0 572 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6523
timestamp 1713453518
transform 1 0 836 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6524
timestamp 1713453518
transform 1 0 772 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6525
timestamp 1713453518
transform 1 0 684 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6526
timestamp 1713453518
transform 1 0 588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6527
timestamp 1713453518
transform 1 0 1236 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_6528
timestamp 1713453518
transform 1 0 1068 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6529
timestamp 1713453518
transform 1 0 852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_6530
timestamp 1713453518
transform 1 0 748 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6531
timestamp 1713453518
transform 1 0 668 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_6532
timestamp 1713453518
transform 1 0 484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6533
timestamp 1713453518
transform 1 0 892 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6534
timestamp 1713453518
transform 1 0 844 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6535
timestamp 1713453518
transform 1 0 828 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6536
timestamp 1713453518
transform 1 0 700 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6537
timestamp 1713453518
transform 1 0 628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6538
timestamp 1713453518
transform 1 0 1412 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1713453518
transform 1 0 1324 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6540
timestamp 1713453518
transform 1 0 1052 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6541
timestamp 1713453518
transform 1 0 828 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6542
timestamp 1713453518
transform 1 0 684 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1713453518
transform 1 0 500 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6544
timestamp 1713453518
transform 1 0 444 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6545
timestamp 1713453518
transform 1 0 1236 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1713453518
transform 1 0 1052 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6547
timestamp 1713453518
transform 1 0 940 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6548
timestamp 1713453518
transform 1 0 924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1713453518
transform 1 0 1116 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_6550
timestamp 1713453518
transform 1 0 1108 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6551
timestamp 1713453518
transform 1 0 1004 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1713453518
transform 1 0 988 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6553
timestamp 1713453518
transform 1 0 1212 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6554
timestamp 1713453518
transform 1 0 1132 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1713453518
transform 1 0 1084 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6556
timestamp 1713453518
transform 1 0 916 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6557
timestamp 1713453518
transform 1 0 1484 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6558
timestamp 1713453518
transform 1 0 1044 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6559
timestamp 1713453518
transform 1 0 940 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6560
timestamp 1713453518
transform 1 0 908 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1713453518
transform 1 0 1260 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1713453518
transform 1 0 1052 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6563
timestamp 1713453518
transform 1 0 884 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1713453518
transform 1 0 868 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6565
timestamp 1713453518
transform 1 0 844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6566
timestamp 1713453518
transform 1 0 1124 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6567
timestamp 1713453518
transform 1 0 1004 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6568
timestamp 1713453518
transform 1 0 868 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6569
timestamp 1713453518
transform 1 0 844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6570
timestamp 1713453518
transform 1 0 812 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6571
timestamp 1713453518
transform 1 0 1092 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6572
timestamp 1713453518
transform 1 0 988 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1713453518
transform 1 0 836 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6574
timestamp 1713453518
transform 1 0 812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6575
timestamp 1713453518
transform 1 0 788 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6576
timestamp 1713453518
transform 1 0 780 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6577
timestamp 1713453518
transform 1 0 1540 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_6578
timestamp 1713453518
transform 1 0 1052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1713453518
transform 1 0 860 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6580
timestamp 1713453518
transform 1 0 844 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1713453518
transform 1 0 764 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1713453518
transform 1 0 732 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6583
timestamp 1713453518
transform 1 0 700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1713453518
transform 1 0 1052 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1713453518
transform 1 0 1004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6586
timestamp 1713453518
transform 1 0 900 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1713453518
transform 1 0 876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6588
timestamp 1713453518
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1713453518
transform 1 0 1468 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_6590
timestamp 1713453518
transform 1 0 1052 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6591
timestamp 1713453518
transform 1 0 1028 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6592
timestamp 1713453518
transform 1 0 860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6593
timestamp 1713453518
transform 1 0 844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6594
timestamp 1713453518
transform 1 0 724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6595
timestamp 1713453518
transform 1 0 692 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6596
timestamp 1713453518
transform 1 0 1628 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_6597
timestamp 1713453518
transform 1 0 956 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6598
timestamp 1713453518
transform 1 0 812 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6599
timestamp 1713453518
transform 1 0 788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6600
timestamp 1713453518
transform 1 0 748 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6601
timestamp 1713453518
transform 1 0 732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6602
timestamp 1713453518
transform 1 0 1012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6603
timestamp 1713453518
transform 1 0 820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6604
timestamp 1713453518
transform 1 0 820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1713453518
transform 1 0 740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6606
timestamp 1713453518
transform 1 0 660 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6607
timestamp 1713453518
transform 1 0 644 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6608
timestamp 1713453518
transform 1 0 1292 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_6609
timestamp 1713453518
transform 1 0 1004 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1713453518
transform 1 0 804 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6611
timestamp 1713453518
transform 1 0 724 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_6612
timestamp 1713453518
transform 1 0 588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6613
timestamp 1713453518
transform 1 0 564 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6614
timestamp 1713453518
transform 1 0 564 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6615
timestamp 1713453518
transform 1 0 1212 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_6616
timestamp 1713453518
transform 1 0 1068 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6617
timestamp 1713453518
transform 1 0 1044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6618
timestamp 1713453518
transform 1 0 860 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6619
timestamp 1713453518
transform 1 0 1444 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_6620
timestamp 1713453518
transform 1 0 1092 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6621
timestamp 1713453518
transform 1 0 1076 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6622
timestamp 1713453518
transform 1 0 1052 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6623
timestamp 1713453518
transform 1 0 908 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6624
timestamp 1713453518
transform 1 0 1412 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6625
timestamp 1713453518
transform 1 0 1052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6626
timestamp 1713453518
transform 1 0 1004 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6627
timestamp 1713453518
transform 1 0 884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6628
timestamp 1713453518
transform 1 0 1444 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6629
timestamp 1713453518
transform 1 0 996 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6630
timestamp 1713453518
transform 1 0 988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6631
timestamp 1713453518
transform 1 0 956 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6632
timestamp 1713453518
transform 1 0 940 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6633
timestamp 1713453518
transform 1 0 1476 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_6634
timestamp 1713453518
transform 1 0 964 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6635
timestamp 1713453518
transform 1 0 780 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6636
timestamp 1713453518
transform 1 0 732 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1713453518
transform 1 0 660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6638
timestamp 1713453518
transform 1 0 1524 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_6639
timestamp 1713453518
transform 1 0 1044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6640
timestamp 1713453518
transform 1 0 868 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6641
timestamp 1713453518
transform 1 0 692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6642
timestamp 1713453518
transform 1 0 564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6643
timestamp 1713453518
transform 1 0 836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6644
timestamp 1713453518
transform 1 0 788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6645
timestamp 1713453518
transform 1 0 692 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6646
timestamp 1713453518
transform 1 0 380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6647
timestamp 1713453518
transform 1 0 356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_6648
timestamp 1713453518
transform 1 0 700 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_6649
timestamp 1713453518
transform 1 0 460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6650
timestamp 1713453518
transform 1 0 420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6651
timestamp 1713453518
transform 1 0 348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_6652
timestamp 1713453518
transform 1 0 772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6653
timestamp 1713453518
transform 1 0 764 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6654
timestamp 1713453518
transform 1 0 732 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6655
timestamp 1713453518
transform 1 0 676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_6656
timestamp 1713453518
transform 1 0 884 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_6657
timestamp 1713453518
transform 1 0 828 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_6658
timestamp 1713453518
transform 1 0 1548 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_6659
timestamp 1713453518
transform 1 0 708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6660
timestamp 1713453518
transform 1 0 644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6661
timestamp 1713453518
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6662
timestamp 1713453518
transform 1 0 1020 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_6663
timestamp 1713453518
transform 1 0 940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6664
timestamp 1713453518
transform 1 0 916 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_6665
timestamp 1713453518
transform 1 0 700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6666
timestamp 1713453518
transform 1 0 612 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1713453518
transform 1 0 548 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6668
timestamp 1713453518
transform 1 0 508 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_6669
timestamp 1713453518
transform 1 0 388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1713453518
transform 1 0 1044 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_6671
timestamp 1713453518
transform 1 0 756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6672
timestamp 1713453518
transform 1 0 532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6673
timestamp 1713453518
transform 1 0 524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_6674
timestamp 1713453518
transform 1 0 428 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_6675
timestamp 1713453518
transform 1 0 1084 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_6676
timestamp 1713453518
transform 1 0 708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6677
timestamp 1713453518
transform 1 0 628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6678
timestamp 1713453518
transform 1 0 1292 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_6679
timestamp 1713453518
transform 1 0 1292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_6680
timestamp 1713453518
transform 1 0 804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6681
timestamp 1713453518
transform 1 0 620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6682
timestamp 1713453518
transform 1 0 612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6683
timestamp 1713453518
transform 1 0 340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6684
timestamp 1713453518
transform 1 0 1052 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_6685
timestamp 1713453518
transform 1 0 948 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6686
timestamp 1713453518
transform 1 0 684 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_6687
timestamp 1713453518
transform 1 0 612 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_6688
timestamp 1713453518
transform 1 0 444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_6689
timestamp 1713453518
transform 1 0 316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6690
timestamp 1713453518
transform 1 0 1116 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_6691
timestamp 1713453518
transform 1 0 748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6692
timestamp 1713453518
transform 1 0 564 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6693
timestamp 1713453518
transform 1 0 436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6694
timestamp 1713453518
transform 1 0 420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_6695
timestamp 1713453518
transform 1 0 1084 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_6696
timestamp 1713453518
transform 1 0 804 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6697
timestamp 1713453518
transform 1 0 660 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6698
timestamp 1713453518
transform 1 0 388 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_6699
timestamp 1713453518
transform 1 0 652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6700
timestamp 1713453518
transform 1 0 652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6701
timestamp 1713453518
transform 1 0 564 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6702
timestamp 1713453518
transform 1 0 436 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6703
timestamp 1713453518
transform 1 0 1060 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_6704
timestamp 1713453518
transform 1 0 724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6705
timestamp 1713453518
transform 1 0 708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6706
timestamp 1713453518
transform 1 0 652 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6707
timestamp 1713453518
transform 1 0 508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6708
timestamp 1713453518
transform 1 0 1044 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6709
timestamp 1713453518
transform 1 0 716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6710
timestamp 1713453518
transform 1 0 716 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6711
timestamp 1713453518
transform 1 0 708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6712
timestamp 1713453518
transform 1 0 700 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6713
timestamp 1713453518
transform 1 0 516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6714
timestamp 1713453518
transform 1 0 428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6715
timestamp 1713453518
transform 1 0 1108 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6716
timestamp 1713453518
transform 1 0 756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6717
timestamp 1713453518
transform 1 0 756 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1713453518
transform 1 0 740 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6719
timestamp 1713453518
transform 1 0 668 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6720
timestamp 1713453518
transform 1 0 420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6721
timestamp 1713453518
transform 1 0 1092 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6722
timestamp 1713453518
transform 1 0 988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6723
timestamp 1713453518
transform 1 0 708 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6724
timestamp 1713453518
transform 1 0 644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1713453518
transform 1 0 620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6726
timestamp 1713453518
transform 1 0 612 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6727
timestamp 1713453518
transform 1 0 428 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6728
timestamp 1713453518
transform 1 0 1108 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6729
timestamp 1713453518
transform 1 0 1068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6730
timestamp 1713453518
transform 1 0 724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6731
timestamp 1713453518
transform 1 0 708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6732
timestamp 1713453518
transform 1 0 700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6733
timestamp 1713453518
transform 1 0 684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6734
timestamp 1713453518
transform 1 0 668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6735
timestamp 1713453518
transform 1 0 396 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6736
timestamp 1713453518
transform 1 0 1204 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6737
timestamp 1713453518
transform 1 0 1108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6738
timestamp 1713453518
transform 1 0 804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6739
timestamp 1713453518
transform 1 0 772 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6740
timestamp 1713453518
transform 1 0 748 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6741
timestamp 1713453518
transform 1 0 652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6742
timestamp 1713453518
transform 1 0 380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6743
timestamp 1713453518
transform 1 0 1116 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_6744
timestamp 1713453518
transform 1 0 1020 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6745
timestamp 1713453518
transform 1 0 788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6746
timestamp 1713453518
transform 1 0 788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6747
timestamp 1713453518
transform 1 0 772 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_6748
timestamp 1713453518
transform 1 0 700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6749
timestamp 1713453518
transform 1 0 444 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6750
timestamp 1713453518
transform 1 0 684 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6751
timestamp 1713453518
transform 1 0 524 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6752
timestamp 1713453518
transform 1 0 476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6753
timestamp 1713453518
transform 1 0 1124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6754
timestamp 1713453518
transform 1 0 1108 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_6755
timestamp 1713453518
transform 1 0 836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6756
timestamp 1713453518
transform 1 0 780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6757
timestamp 1713453518
transform 1 0 468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6758
timestamp 1713453518
transform 1 0 1044 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_6759
timestamp 1713453518
transform 1 0 820 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6760
timestamp 1713453518
transform 1 0 772 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6761
timestamp 1713453518
transform 1 0 652 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_6762
timestamp 1713453518
transform 1 0 468 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6763
timestamp 1713453518
transform 1 0 1116 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_6764
timestamp 1713453518
transform 1 0 876 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6765
timestamp 1713453518
transform 1 0 708 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6766
timestamp 1713453518
transform 1 0 652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6767
timestamp 1713453518
transform 1 0 508 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6768
timestamp 1713453518
transform 1 0 1108 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_6769
timestamp 1713453518
transform 1 0 876 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6770
timestamp 1713453518
transform 1 0 612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6771
timestamp 1713453518
transform 1 0 604 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6772
timestamp 1713453518
transform 1 0 548 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6773
timestamp 1713453518
transform 1 0 1124 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6774
timestamp 1713453518
transform 1 0 844 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6775
timestamp 1713453518
transform 1 0 700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6776
timestamp 1713453518
transform 1 0 660 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6777
timestamp 1713453518
transform 1 0 420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6778
timestamp 1713453518
transform 1 0 1076 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6779
timestamp 1713453518
transform 1 0 876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6780
timestamp 1713453518
transform 1 0 764 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6781
timestamp 1713453518
transform 1 0 708 0 1 2555
box -2 -2 2 2
use M2_M1  M2_M1_6782
timestamp 1713453518
transform 1 0 660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6783
timestamp 1713453518
transform 1 0 452 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6784
timestamp 1713453518
transform 1 0 1092 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6785
timestamp 1713453518
transform 1 0 900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6786
timestamp 1713453518
transform 1 0 756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6787
timestamp 1713453518
transform 1 0 692 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6788
timestamp 1713453518
transform 1 0 580 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6789
timestamp 1713453518
transform 1 0 508 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6790
timestamp 1713453518
transform 1 0 884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6791
timestamp 1713453518
transform 1 0 780 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6792
timestamp 1713453518
transform 1 0 652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6793
timestamp 1713453518
transform 1 0 468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6794
timestamp 1713453518
transform 1 0 1140 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6795
timestamp 1713453518
transform 1 0 1140 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6796
timestamp 1713453518
transform 1 0 788 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6797
timestamp 1713453518
transform 1 0 740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6798
timestamp 1713453518
transform 1 0 684 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6799
timestamp 1713453518
transform 1 0 668 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6800
timestamp 1713453518
transform 1 0 1036 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6801
timestamp 1713453518
transform 1 0 1036 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6802
timestamp 1713453518
transform 1 0 756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6803
timestamp 1713453518
transform 1 0 716 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6804
timestamp 1713453518
transform 1 0 668 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6805
timestamp 1713453518
transform 1 0 636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6806
timestamp 1713453518
transform 1 0 1100 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6807
timestamp 1713453518
transform 1 0 980 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6808
timestamp 1713453518
transform 1 0 748 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6809
timestamp 1713453518
transform 1 0 676 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6810
timestamp 1713453518
transform 1 0 564 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6811
timestamp 1713453518
transform 1 0 548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6812
timestamp 1713453518
transform 1 0 444 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6813
timestamp 1713453518
transform 1 0 428 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6814
timestamp 1713453518
transform 1 0 1220 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6815
timestamp 1713453518
transform 1 0 1204 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6816
timestamp 1713453518
transform 1 0 860 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6817
timestamp 1713453518
transform 1 0 588 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6818
timestamp 1713453518
transform 1 0 1172 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6819
timestamp 1713453518
transform 1 0 1164 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6820
timestamp 1713453518
transform 1 0 732 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6821
timestamp 1713453518
transform 1 0 676 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6822
timestamp 1713453518
transform 1 0 500 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6823
timestamp 1713453518
transform 1 0 1180 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6824
timestamp 1713453518
transform 1 0 1052 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6825
timestamp 1713453518
transform 1 0 788 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6826
timestamp 1713453518
transform 1 0 668 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6827
timestamp 1713453518
transform 1 0 524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6828
timestamp 1713453518
transform 1 0 1732 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6829
timestamp 1713453518
transform 1 0 1716 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_6830
timestamp 1713453518
transform 1 0 1804 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_6831
timestamp 1713453518
transform 1 0 1772 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6832
timestamp 1713453518
transform 1 0 2820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6833
timestamp 1713453518
transform 1 0 2796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6834
timestamp 1713453518
transform 1 0 1380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6835
timestamp 1713453518
transform 1 0 1268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6836
timestamp 1713453518
transform 1 0 1260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_6837
timestamp 1713453518
transform 1 0 892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6838
timestamp 1713453518
transform 1 0 604 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6839
timestamp 1713453518
transform 1 0 508 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_6840
timestamp 1713453518
transform 1 0 484 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_6841
timestamp 1713453518
transform 1 0 468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_6842
timestamp 1713453518
transform 1 0 452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_6843
timestamp 1713453518
transform 1 0 452 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_6844
timestamp 1713453518
transform 1 0 436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6845
timestamp 1713453518
transform 1 0 716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6846
timestamp 1713453518
transform 1 0 700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6847
timestamp 1713453518
transform 1 0 668 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_6848
timestamp 1713453518
transform 1 0 76 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6849
timestamp 1713453518
transform 1 0 1268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6850
timestamp 1713453518
transform 1 0 1036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_6851
timestamp 1713453518
transform 1 0 388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_6852
timestamp 1713453518
transform 1 0 380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_6853
timestamp 1713453518
transform 1 0 324 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1713453518
transform 1 0 2540 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1713453518
transform 1 0 2508 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1713453518
transform 1 0 2772 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1713453518
transform 1 0 2620 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1713453518
transform 1 0 1204 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1713453518
transform 1 0 1140 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1713453518
transform 1 0 1412 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1713453518
transform 1 0 1292 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1713453518
transform 1 0 1212 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1713453518
transform 1 0 1180 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1713453518
transform 1 0 1668 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1713453518
transform 1 0 1228 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1713453518
transform 1 0 1148 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1713453518
transform 1 0 1676 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1713453518
transform 1 0 1596 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1713453518
transform 1 0 1580 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1713453518
transform 1 0 1244 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1713453518
transform 1 0 1228 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1713453518
transform 1 0 1220 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1713453518
transform 1 0 1156 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1713453518
transform 1 0 1124 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1713453518
transform 1 0 1756 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1713453518
transform 1 0 1244 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1713453518
transform 1 0 1244 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1713453518
transform 1 0 1228 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1713453518
transform 1 0 1220 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1713453518
transform 1 0 1140 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1713453518
transform 1 0 1884 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1713453518
transform 1 0 1668 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1713453518
transform 1 0 1652 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1713453518
transform 1 0 1588 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1713453518
transform 1 0 1548 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1713453518
transform 1 0 1548 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1713453518
transform 1 0 1484 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1713453518
transform 1 0 1460 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1713453518
transform 1 0 1764 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1713453518
transform 1 0 1580 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1713453518
transform 1 0 1556 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1713453518
transform 1 0 1516 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1713453518
transform 1 0 1364 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1713453518
transform 1 0 1324 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1713453518
transform 1 0 1324 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1713453518
transform 1 0 1284 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1713453518
transform 1 0 1284 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1713453518
transform 1 0 1252 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1713453518
transform 1 0 1252 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1713453518
transform 1 0 3412 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1713453518
transform 1 0 3396 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1713453518
transform 1 0 3356 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1713453518
transform 1 0 3348 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1713453518
transform 1 0 3276 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1713453518
transform 1 0 3444 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1713453518
transform 1 0 3308 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1713453518
transform 1 0 3340 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1713453518
transform 1 0 3252 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1713453518
transform 1 0 3220 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1713453518
transform 1 0 2276 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1713453518
transform 1 0 2172 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1713453518
transform 1 0 2140 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1713453518
transform 1 0 2380 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1713453518
transform 1 0 2244 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1713453518
transform 1 0 396 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1713453518
transform 1 0 316 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1713453518
transform 1 0 724 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1713453518
transform 1 0 668 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1713453518
transform 1 0 172 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1713453518
transform 1 0 100 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1713453518
transform 1 0 180 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1713453518
transform 1 0 84 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1713453518
transform 1 0 292 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1713453518
transform 1 0 212 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1713453518
transform 1 0 172 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1713453518
transform 1 0 124 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1713453518
transform 1 0 244 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1713453518
transform 1 0 204 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1713453518
transform 1 0 172 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1713453518
transform 1 0 140 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1713453518
transform 1 0 660 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1713453518
transform 1 0 540 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1713453518
transform 1 0 396 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1713453518
transform 1 0 932 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1713453518
transform 1 0 772 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1713453518
transform 1 0 444 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1713453518
transform 1 0 604 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1713453518
transform 1 0 404 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1713453518
transform 1 0 420 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1713453518
transform 1 0 356 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1713453518
transform 1 0 308 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1713453518
transform 1 0 476 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1713453518
transform 1 0 180 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1713453518
transform 1 0 428 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1713453518
transform 1 0 252 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1713453518
transform 1 0 220 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1713453518
transform 1 0 1348 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1713453518
transform 1 0 1244 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1713453518
transform 1 0 1308 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1713453518
transform 1 0 1268 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1713453518
transform 1 0 988 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1713453518
transform 1 0 900 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1713453518
transform 1 0 1028 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1713453518
transform 1 0 876 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1713453518
transform 1 0 996 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1713453518
transform 1 0 828 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1713453518
transform 1 0 932 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1713453518
transform 1 0 796 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1713453518
transform 1 0 988 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1713453518
transform 1 0 756 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1713453518
transform 1 0 980 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1713453518
transform 1 0 772 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1713453518
transform 1 0 932 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1713453518
transform 1 0 796 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1713453518
transform 1 0 1004 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1713453518
transform 1 0 772 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1713453518
transform 1 0 908 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1713453518
transform 1 0 804 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1713453518
transform 1 0 1028 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1713453518
transform 1 0 908 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1713453518
transform 1 0 948 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1713453518
transform 1 0 796 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1713453518
transform 1 0 1044 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1713453518
transform 1 0 908 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1713453518
transform 1 0 1044 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1713453518
transform 1 0 940 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1713453518
transform 1 0 1004 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1713453518
transform 1 0 900 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1713453518
transform 1 0 988 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1713453518
transform 1 0 820 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1713453518
transform 1 0 972 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1713453518
transform 1 0 844 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1713453518
transform 1 0 948 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1713453518
transform 1 0 812 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1713453518
transform 1 0 1004 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1713453518
transform 1 0 868 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1713453518
transform 1 0 1028 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1713453518
transform 1 0 868 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1713453518
transform 1 0 980 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1713453518
transform 1 0 836 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1713453518
transform 1 0 996 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1713453518
transform 1 0 860 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1713453518
transform 1 0 1044 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1713453518
transform 1 0 892 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1713453518
transform 1 0 1076 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1713453518
transform 1 0 932 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1713453518
transform 1 0 1100 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1713453518
transform 1 0 1020 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1713453518
transform 1 0 972 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1713453518
transform 1 0 876 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1713453518
transform 1 0 876 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1713453518
transform 1 0 852 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1713453518
transform 1 0 828 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1713453518
transform 1 0 804 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1713453518
transform 1 0 884 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1713453518
transform 1 0 740 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1713453518
transform 1 0 772 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1713453518
transform 1 0 524 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1713453518
transform 1 0 836 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1713453518
transform 1 0 524 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1713453518
transform 1 0 764 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1713453518
transform 1 0 708 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1713453518
transform 1 0 756 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1713453518
transform 1 0 196 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1713453518
transform 1 0 724 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1713453518
transform 1 0 356 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1713453518
transform 1 0 700 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1713453518
transform 1 0 284 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1713453518
transform 1 0 764 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1713453518
transform 1 0 316 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1713453518
transform 1 0 740 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1713453518
transform 1 0 396 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1713453518
transform 1 0 756 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1713453518
transform 1 0 452 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1713453518
transform 1 0 844 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1713453518
transform 1 0 396 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1713453518
transform 1 0 740 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1713453518
transform 1 0 380 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1713453518
transform 1 0 924 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1713453518
transform 1 0 868 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1713453518
transform 1 0 868 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1713453518
transform 1 0 820 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1713453518
transform 1 0 844 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1713453518
transform 1 0 404 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1713453518
transform 1 0 756 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1713453518
transform 1 0 436 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1713453518
transform 1 0 804 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1713453518
transform 1 0 436 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1713453518
transform 1 0 748 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1713453518
transform 1 0 436 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1713453518
transform 1 0 812 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1713453518
transform 1 0 564 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1713453518
transform 1 0 796 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1713453518
transform 1 0 388 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1713453518
transform 1 0 788 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1713453518
transform 1 0 420 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1713453518
transform 1 0 812 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1713453518
transform 1 0 476 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1713453518
transform 1 0 836 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1713453518
transform 1 0 484 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1713453518
transform 1 0 924 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1713453518
transform 1 0 436 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1713453518
transform 1 0 900 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1713453518
transform 1 0 804 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1713453518
transform 1 0 972 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1713453518
transform 1 0 780 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1713453518
transform 1 0 884 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1713453518
transform 1 0 468 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1713453518
transform 1 0 812 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1713453518
transform 1 0 500 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1713453518
transform 1 0 812 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1713453518
transform 1 0 364 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1713453518
transform 1 0 708 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1713453518
transform 1 0 444 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1713453518
transform 1 0 700 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1713453518
transform 1 0 380 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1713453518
transform 1 0 2484 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1713453518
transform 1 0 2388 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1713453518
transform 1 0 2340 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1713453518
transform 1 0 1868 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1713453518
transform 1 0 1868 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1713453518
transform 1 0 1108 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1713453518
transform 1 0 2620 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1713453518
transform 1 0 2532 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1713453518
transform 1 0 2524 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1713453518
transform 1 0 2500 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1713453518
transform 1 0 2436 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1713453518
transform 1 0 2204 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1713453518
transform 1 0 2204 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1713453518
transform 1 0 2036 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1713453518
transform 1 0 1900 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1713453518
transform 1 0 1900 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1713453518
transform 1 0 1804 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1713453518
transform 1 0 1380 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1713453518
transform 1 0 2644 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1713453518
transform 1 0 2556 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1713453518
transform 1 0 1700 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1713453518
transform 1 0 1636 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1713453518
transform 1 0 2980 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1713453518
transform 1 0 2924 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1713453518
transform 1 0 2772 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1713453518
transform 1 0 1628 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1713453518
transform 1 0 3068 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1713453518
transform 1 0 2932 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1713453518
transform 1 0 2932 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1713453518
transform 1 0 1748 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1713453518
transform 1 0 2252 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1713453518
transform 1 0 1892 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1713453518
transform 1 0 1892 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1713453518
transform 1 0 1852 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1713453518
transform 1 0 2412 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1713453518
transform 1 0 2364 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1713453518
transform 1 0 2092 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1713453518
transform 1 0 2060 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1713453518
transform 1 0 1740 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1713453518
transform 1 0 2356 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1713453518
transform 1 0 2220 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1713453518
transform 1 0 2572 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1713453518
transform 1 0 2500 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1713453518
transform 1 0 2396 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1713453518
transform 1 0 3332 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1713453518
transform 1 0 2900 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1713453518
transform 1 0 2900 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1713453518
transform 1 0 2324 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1713453518
transform 1 0 2764 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1713453518
transform 1 0 2644 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1713453518
transform 1 0 3196 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1713453518
transform 1 0 2716 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1713453518
transform 1 0 2452 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1713453518
transform 1 0 3316 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1713453518
transform 1 0 3012 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1713453518
transform 1 0 3140 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1713453518
transform 1 0 3092 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1713453518
transform 1 0 3092 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1713453518
transform 1 0 3044 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1713453518
transform 1 0 348 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1713453518
transform 1 0 204 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1713453518
transform 1 0 900 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1713453518
transform 1 0 828 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1713453518
transform 1 0 780 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1713453518
transform 1 0 740 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1713453518
transform 1 0 660 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1713453518
transform 1 0 564 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1713453518
transform 1 0 988 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1713453518
transform 1 0 908 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1713453518
transform 1 0 836 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1713453518
transform 1 0 756 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1713453518
transform 1 0 876 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1713453518
transform 1 0 772 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1713453518
transform 1 0 764 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1713453518
transform 1 0 668 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1713453518
transform 1 0 2948 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1713453518
transform 1 0 2852 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1713453518
transform 1 0 2748 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1713453518
transform 1 0 2700 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1713453518
transform 1 0 2532 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1713453518
transform 1 0 2516 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1713453518
transform 1 0 3036 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1713453518
transform 1 0 2156 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1713453518
transform 1 0 2052 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1713453518
transform 1 0 2044 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1713453518
transform 1 0 2004 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1713453518
transform 1 0 1972 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1713453518
transform 1 0 1972 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1713453518
transform 1 0 1956 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1713453518
transform 1 0 1956 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1713453518
transform 1 0 1932 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1713453518
transform 1 0 1892 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1713453518
transform 1 0 1852 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1713453518
transform 1 0 1804 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1713453518
transform 1 0 2364 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1713453518
transform 1 0 2284 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1713453518
transform 1 0 2284 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1713453518
transform 1 0 2196 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1713453518
transform 1 0 2148 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1713453518
transform 1 0 2412 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1713453518
transform 1 0 2356 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1713453518
transform 1 0 2348 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1713453518
transform 1 0 2300 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1713453518
transform 1 0 1564 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1713453518
transform 1 0 1532 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1713453518
transform 1 0 1644 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1713453518
transform 1 0 1644 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1713453518
transform 1 0 1636 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1713453518
transform 1 0 1628 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1713453518
transform 1 0 1620 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1713453518
transform 1 0 1620 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1713453518
transform 1 0 1596 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1713453518
transform 1 0 1588 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1713453518
transform 1 0 1588 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1713453518
transform 1 0 1524 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1713453518
transform 1 0 1524 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1713453518
transform 1 0 1500 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1713453518
transform 1 0 1500 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1713453518
transform 1 0 1476 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1713453518
transform 1 0 1444 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1713453518
transform 1 0 1436 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1713453518
transform 1 0 1340 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1713453518
transform 1 0 1284 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1713453518
transform 1 0 1284 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1713453518
transform 1 0 1268 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1713453518
transform 1 0 1260 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1713453518
transform 1 0 1244 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1713453518
transform 1 0 1236 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1713453518
transform 1 0 1236 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1713453518
transform 1 0 1148 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1713453518
transform 1 0 1116 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1713453518
transform 1 0 1116 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1713453518
transform 1 0 1092 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1713453518
transform 1 0 1092 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1713453518
transform 1 0 1404 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1713453518
transform 1 0 1348 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1713453518
transform 1 0 1364 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1713453518
transform 1 0 1316 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1713453518
transform 1 0 1316 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1713453518
transform 1 0 1276 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1713453518
transform 1 0 1540 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1713453518
transform 1 0 1516 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1713453518
transform 1 0 1492 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1713453518
transform 1 0 1484 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1713453518
transform 1 0 1484 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1713453518
transform 1 0 1484 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1713453518
transform 1 0 1460 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1713453518
transform 1 0 1428 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1713453518
transform 1 0 1428 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1713453518
transform 1 0 1420 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1713453518
transform 1 0 1412 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1713453518
transform 1 0 1404 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1713453518
transform 1 0 1380 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1713453518
transform 1 0 1372 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1713453518
transform 1 0 1292 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1713453518
transform 1 0 1276 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1713453518
transform 1 0 1268 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1713453518
transform 1 0 1244 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1713453518
transform 1 0 1236 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1713453518
transform 1 0 1188 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1713453518
transform 1 0 3276 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1713453518
transform 1 0 3260 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1713453518
transform 1 0 3220 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1713453518
transform 1 0 3212 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1713453518
transform 1 0 3396 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1713453518
transform 1 0 3364 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1713453518
transform 1 0 3172 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1713453518
transform 1 0 3100 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1713453518
transform 1 0 3100 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1713453518
transform 1 0 2596 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1713453518
transform 1 0 3348 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1713453518
transform 1 0 3284 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1713453518
transform 1 0 1276 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1713453518
transform 1 0 1236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1713453518
transform 1 0 1196 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1713453518
transform 1 0 1100 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1713453518
transform 1 0 1076 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1713453518
transform 1 0 1012 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1713453518
transform 1 0 2564 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1713453518
transform 1 0 2508 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1713453518
transform 1 0 2492 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1713453518
transform 1 0 2412 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1713453518
transform 1 0 2412 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1713453518
transform 1 0 2300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1713453518
transform 1 0 2300 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1713453518
transform 1 0 2156 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1713453518
transform 1 0 2140 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1713453518
transform 1 0 1340 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1713453518
transform 1 0 1340 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1713453518
transform 1 0 1164 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1713453518
transform 1 0 1164 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1713453518
transform 1 0 1092 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1713453518
transform 1 0 1084 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1713453518
transform 1 0 1068 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1713453518
transform 1 0 1028 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1713453518
transform 1 0 1204 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1713453518
transform 1 0 1180 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1713453518
transform 1 0 1260 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1713453518
transform 1 0 1156 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1713453518
transform 1 0 1100 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1713453518
transform 1 0 1188 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1713453518
transform 1 0 1188 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1713453518
transform 1 0 1180 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1713453518
transform 1 0 1132 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1713453518
transform 1 0 1116 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1713453518
transform 1 0 1108 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1713453518
transform 1 0 1076 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1713453518
transform 1 0 1332 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1713453518
transform 1 0 1244 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1713453518
transform 1 0 1396 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1713453518
transform 1 0 1396 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1713453518
transform 1 0 1388 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1713453518
transform 1 0 1388 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1713453518
transform 1 0 1356 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1713453518
transform 1 0 1300 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1713453518
transform 1 0 1292 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1713453518
transform 1 0 1284 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1713453518
transform 1 0 1284 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1713453518
transform 1 0 1236 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1713453518
transform 1 0 1236 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1713453518
transform 1 0 1188 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1713453518
transform 1 0 1172 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1713453518
transform 1 0 1172 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1713453518
transform 1 0 1164 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1713453518
transform 1 0 1148 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1713453518
transform 1 0 1148 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1713453518
transform 1 0 1108 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1713453518
transform 1 0 1108 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1713453518
transform 1 0 1436 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1713453518
transform 1 0 1212 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1713453518
transform 1 0 1188 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1713453518
transform 1 0 1156 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1713453518
transform 1 0 1572 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1713453518
transform 1 0 1524 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1713453518
transform 1 0 1492 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1713453518
transform 1 0 1532 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1713453518
transform 1 0 1516 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1713453518
transform 1 0 1484 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1713453518
transform 1 0 1436 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1713453518
transform 1 0 1340 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1713453518
transform 1 0 1340 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1713453518
transform 1 0 1316 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1713453518
transform 1 0 1292 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1713453518
transform 1 0 1220 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1713453518
transform 1 0 1404 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1713453518
transform 1 0 1380 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1713453518
transform 1 0 1204 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1713453518
transform 1 0 1172 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1713453518
transform 1 0 1172 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1713453518
transform 1 0 1148 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1713453518
transform 1 0 1148 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1713453518
transform 1 0 1148 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1713453518
transform 1 0 1108 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1713453518
transform 1 0 1620 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1713453518
transform 1 0 1524 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1713453518
transform 1 0 1252 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1713453518
transform 1 0 1244 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1713453518
transform 1 0 1212 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1713453518
transform 1 0 1140 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1713453518
transform 1 0 1644 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1713453518
transform 1 0 1612 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1713453518
transform 1 0 1460 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1713453518
transform 1 0 1260 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1713453518
transform 1 0 1260 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1713453518
transform 1 0 1212 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1713453518
transform 1 0 1204 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1713453518
transform 1 0 1172 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1713453518
transform 1 0 1404 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1713453518
transform 1 0 1396 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1713453518
transform 1 0 1396 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1713453518
transform 1 0 1396 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1713453518
transform 1 0 1380 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1713453518
transform 1 0 1380 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1713453518
transform 1 0 1364 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1713453518
transform 1 0 1356 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1713453518
transform 1 0 1340 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1713453518
transform 1 0 1332 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1713453518
transform 1 0 1332 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1713453518
transform 1 0 1324 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1713453518
transform 1 0 1292 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1713453518
transform 1 0 1260 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1713453518
transform 1 0 1228 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1713453518
transform 1 0 1132 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1713453518
transform 1 0 1132 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1713453518
transform 1 0 1108 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1713453518
transform 1 0 1436 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1713453518
transform 1 0 1388 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1713453518
transform 1 0 1340 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1713453518
transform 1 0 1332 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1713453518
transform 1 0 1276 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1713453518
transform 1 0 1180 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1713453518
transform 1 0 1700 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1713453518
transform 1 0 1636 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1713453518
transform 1 0 1332 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1713453518
transform 1 0 1324 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1713453518
transform 1 0 1300 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1713453518
transform 1 0 1276 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1713453518
transform 1 0 1212 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1713453518
transform 1 0 1644 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1713453518
transform 1 0 1596 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1713453518
transform 1 0 1468 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1713453518
transform 1 0 1420 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1713453518
transform 1 0 1412 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1713453518
transform 1 0 1396 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1713453518
transform 1 0 1388 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1713453518
transform 1 0 1236 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1713453518
transform 1 0 1188 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1713453518
transform 1 0 1724 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1713453518
transform 1 0 1684 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1713453518
transform 1 0 1420 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1713453518
transform 1 0 1388 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1713453518
transform 1 0 1356 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1713453518
transform 1 0 1316 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1713453518
transform 1 0 1164 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1713453518
transform 1 0 1156 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1713453518
transform 1 0 1156 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1713453518
transform 1 0 1124 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1713453518
transform 1 0 1124 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1713453518
transform 1 0 1124 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1713453518
transform 1 0 1116 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1713453518
transform 1 0 1380 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1713453518
transform 1 0 1284 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1713453518
transform 1 0 1172 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1713453518
transform 1 0 1684 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1713453518
transform 1 0 1556 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1713453518
transform 1 0 1556 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1713453518
transform 1 0 1460 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1713453518
transform 1 0 1636 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1713453518
transform 1 0 1612 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1713453518
transform 1 0 1572 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1713453518
transform 1 0 1508 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1713453518
transform 1 0 1508 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1713453518
transform 1 0 1436 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1713453518
transform 1 0 1108 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1713453518
transform 1 0 1100 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1713453518
transform 1 0 1100 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1713453518
transform 1 0 1052 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1713453518
transform 1 0 1012 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1713453518
transform 1 0 1012 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1713453518
transform 1 0 1444 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1713453518
transform 1 0 1396 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1713453518
transform 1 0 1388 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1713453518
transform 1 0 1380 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1713453518
transform 1 0 1364 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1713453518
transform 1 0 1180 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1713453518
transform 1 0 1164 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1713453518
transform 1 0 1156 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1713453518
transform 1 0 1148 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1713453518
transform 1 0 1364 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1713453518
transform 1 0 1204 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1713453518
transform 1 0 1172 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1713453518
transform 1 0 1628 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1713453518
transform 1 0 1492 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1713453518
transform 1 0 1492 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1713453518
transform 1 0 1476 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1713453518
transform 1 0 1452 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1713453518
transform 1 0 1532 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1713453518
transform 1 0 1484 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1713453518
transform 1 0 1476 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1713453518
transform 1 0 1444 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1713453518
transform 1 0 1444 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1713453518
transform 1 0 1396 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1713453518
transform 1 0 1348 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1713453518
transform 1 0 1340 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1713453518
transform 1 0 1324 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1713453518
transform 1 0 1324 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1713453518
transform 1 0 1308 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1713453518
transform 1 0 1308 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1713453518
transform 1 0 1308 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1713453518
transform 1 0 1292 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1713453518
transform 1 0 1284 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1713453518
transform 1 0 1180 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1713453518
transform 1 0 1180 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1713453518
transform 1 0 1164 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1713453518
transform 1 0 1140 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1713453518
transform 1 0 1140 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1713453518
transform 1 0 1108 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1713453518
transform 1 0 1100 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1713453518
transform 1 0 1708 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1713453518
transform 1 0 1708 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1713453518
transform 1 0 1652 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1713453518
transform 1 0 1580 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1713453518
transform 1 0 1500 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1713453518
transform 1 0 1492 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1713453518
transform 1 0 1684 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1713453518
transform 1 0 1628 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1713453518
transform 1 0 1612 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1713453518
transform 1 0 1524 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1713453518
transform 1 0 1492 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1713453518
transform 1 0 1492 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1713453518
transform 1 0 1460 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1713453518
transform 1 0 1548 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1713453518
transform 1 0 1524 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1713453518
transform 1 0 1460 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1713453518
transform 1 0 1428 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1713453518
transform 1 0 1428 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1713453518
transform 1 0 1412 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1713453518
transform 1 0 1412 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1713453518
transform 1 0 1396 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1713453518
transform 1 0 1396 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1713453518
transform 1 0 1388 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1713453518
transform 1 0 1620 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1713453518
transform 1 0 1492 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1713453518
transform 1 0 1244 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1713453518
transform 1 0 1204 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1713453518
transform 1 0 1676 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1713453518
transform 1 0 1604 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1713453518
transform 1 0 1492 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1713453518
transform 1 0 1316 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1713453518
transform 1 0 1268 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1713453518
transform 1 0 1252 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1713453518
transform 1 0 1212 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1713453518
transform 1 0 1132 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1713453518
transform 1 0 1612 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1713453518
transform 1 0 1548 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1713453518
transform 1 0 1452 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1713453518
transform 1 0 1436 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1713453518
transform 1 0 1540 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1713453518
transform 1 0 1412 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1713453518
transform 1 0 1372 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1713453518
transform 1 0 1340 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1713453518
transform 1 0 2460 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1713453518
transform 1 0 1692 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1713453518
transform 1 0 3084 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1713453518
transform 1 0 2996 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1713453518
transform 1 0 3124 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1713453518
transform 1 0 3060 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1713453518
transform 1 0 3020 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1713453518
transform 1 0 2908 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1713453518
transform 1 0 3316 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1713453518
transform 1 0 3276 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1713453518
transform 1 0 3420 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1713453518
transform 1 0 3380 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1713453518
transform 1 0 3308 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1713453518
transform 1 0 3268 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1713453518
transform 1 0 2796 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1713453518
transform 1 0 3396 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1713453518
transform 1 0 3388 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1713453518
transform 1 0 3332 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1713453518
transform 1 0 3316 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1713453518
transform 1 0 3316 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1713453518
transform 1 0 3268 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1713453518
transform 1 0 3260 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1713453518
transform 1 0 3204 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1713453518
transform 1 0 3076 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1713453518
transform 1 0 3428 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1713453518
transform 1 0 3428 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1713453518
transform 1 0 3388 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1713453518
transform 1 0 3388 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1713453518
transform 1 0 3380 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1713453518
transform 1 0 3020 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1713453518
transform 1 0 3020 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1713453518
transform 1 0 2820 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1713453518
transform 1 0 2244 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1713453518
transform 1 0 2244 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1713453518
transform 1 0 2164 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1713453518
transform 1 0 3412 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1713453518
transform 1 0 2812 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1713453518
transform 1 0 2740 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1713453518
transform 1 0 2708 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1713453518
transform 1 0 2676 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1713453518
transform 1 0 2148 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1713453518
transform 1 0 2900 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1713453518
transform 1 0 2772 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1713453518
transform 1 0 2772 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1713453518
transform 1 0 2628 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1713453518
transform 1 0 2612 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1713453518
transform 1 0 2124 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1713453518
transform 1 0 1900 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1713453518
transform 1 0 1900 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1713453518
transform 1 0 1796 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1713453518
transform 1 0 3428 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1713453518
transform 1 0 3292 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1713453518
transform 1 0 3244 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1713453518
transform 1 0 3244 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1713453518
transform 1 0 3220 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1713453518
transform 1 0 3052 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1713453518
transform 1 0 2988 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1713453518
transform 1 0 2444 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1713453518
transform 1 0 1860 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1713453518
transform 1 0 1852 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1713453518
transform 1 0 1724 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1713453518
transform 1 0 3364 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1713453518
transform 1 0 3356 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1713453518
transform 1 0 3340 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1713453518
transform 1 0 3340 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1713453518
transform 1 0 3316 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1713453518
transform 1 0 3316 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1713453518
transform 1 0 3100 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1713453518
transform 1 0 2924 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1713453518
transform 1 0 3372 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1713453518
transform 1 0 3348 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1713453518
transform 1 0 3348 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1713453518
transform 1 0 3044 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1713453518
transform 1 0 2980 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1713453518
transform 1 0 2764 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1713453518
transform 1 0 2684 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1713453518
transform 1 0 2684 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1713453518
transform 1 0 1980 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1713453518
transform 1 0 1980 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1713453518
transform 1 0 1964 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1713453518
transform 1 0 1948 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1713453518
transform 1 0 1948 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1713453518
transform 1 0 3252 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1713453518
transform 1 0 3228 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1713453518
transform 1 0 3164 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1713453518
transform 1 0 3156 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1713453518
transform 1 0 3124 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1713453518
transform 1 0 3116 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1713453518
transform 1 0 2588 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1713453518
transform 1 0 2412 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1713453518
transform 1 0 2412 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1713453518
transform 1 0 2372 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1713453518
transform 1 0 2092 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1713453518
transform 1 0 1428 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1713453518
transform 1 0 2956 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1713453518
transform 1 0 2924 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1713453518
transform 1 0 2852 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1713453518
transform 1 0 2548 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1713453518
transform 1 0 1924 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1713453518
transform 1 0 1924 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1713453518
transform 1 0 1836 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1713453518
transform 1 0 3180 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1713453518
transform 1 0 3116 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1713453518
transform 1 0 3020 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1713453518
transform 1 0 2964 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1713453518
transform 1 0 2964 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1713453518
transform 1 0 2868 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1713453518
transform 1 0 2860 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1713453518
transform 1 0 2812 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1713453518
transform 1 0 3308 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1713453518
transform 1 0 3092 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1713453518
transform 1 0 3060 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1713453518
transform 1 0 3036 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1713453518
transform 1 0 3036 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1713453518
transform 1 0 2980 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1713453518
transform 1 0 2876 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1713453518
transform 1 0 2300 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1713453518
transform 1 0 3340 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1713453518
transform 1 0 3292 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1713453518
transform 1 0 3372 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1713453518
transform 1 0 3340 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1713453518
transform 1 0 3308 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1713453518
transform 1 0 3292 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1713453518
transform 1 0 3196 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1713453518
transform 1 0 3300 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1713453518
transform 1 0 1804 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1713453518
transform 1 0 3372 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1713453518
transform 1 0 2972 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1713453518
transform 1 0 1916 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1713453518
transform 1 0 1836 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1713453518
transform 1 0 1828 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1713453518
transform 1 0 1764 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1713453518
transform 1 0 2884 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1713453518
transform 1 0 2788 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1713453518
transform 1 0 2652 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1713453518
transform 1 0 2652 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1713453518
transform 1 0 1980 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1713453518
transform 1 0 1508 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1713453518
transform 1 0 2748 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1713453518
transform 1 0 2364 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1713453518
transform 1 0 2284 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1713453518
transform 1 0 2284 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1713453518
transform 1 0 2188 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1713453518
transform 1 0 2188 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1713453518
transform 1 0 1948 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1713453518
transform 1 0 2916 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1713453518
transform 1 0 2836 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1713453518
transform 1 0 2788 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1713453518
transform 1 0 2764 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1713453518
transform 1 0 2652 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1713453518
transform 1 0 2644 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1713453518
transform 1 0 2548 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1713453518
transform 1 0 3380 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1713453518
transform 1 0 3340 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1713453518
transform 1 0 3308 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1713453518
transform 1 0 2796 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1713453518
transform 1 0 2652 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1713453518
transform 1 0 2212 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1713453518
transform 1 0 2252 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1713453518
transform 1 0 2036 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1713453518
transform 1 0 2036 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1713453518
transform 1 0 1900 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1713453518
transform 1 0 2196 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1713453518
transform 1 0 2084 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1713453518
transform 1 0 1748 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1713453518
transform 1 0 2884 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1713453518
transform 1 0 2836 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1713453518
transform 1 0 2612 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1713453518
transform 1 0 2612 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1713453518
transform 1 0 2588 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1713453518
transform 1 0 2580 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1713453518
transform 1 0 1908 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1713453518
transform 1 0 3444 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1713453518
transform 1 0 3436 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1713453518
transform 1 0 3380 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1713453518
transform 1 0 3348 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1713453518
transform 1 0 3348 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1713453518
transform 1 0 3220 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1713453518
transform 1 0 3212 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1713453518
transform 1 0 3148 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1713453518
transform 1 0 3044 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1713453518
transform 1 0 1820 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1713453518
transform 1 0 1812 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1713453518
transform 1 0 1684 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1713453518
transform 1 0 3052 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1713453518
transform 1 0 2820 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1713453518
transform 1 0 2820 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1713453518
transform 1 0 2676 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1713453518
transform 1 0 2668 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1713453518
transform 1 0 2124 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1713453518
transform 1 0 3180 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1713453518
transform 1 0 3036 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1713453518
transform 1 0 3036 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1713453518
transform 1 0 2732 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1713453518
transform 1 0 2732 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1713453518
transform 1 0 2692 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1713453518
transform 1 0 2692 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1713453518
transform 1 0 2644 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1713453518
transform 1 0 2644 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1713453518
transform 1 0 2476 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1713453518
transform 1 0 2468 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1713453518
transform 1 0 2436 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1713453518
transform 1 0 2436 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1713453518
transform 1 0 2308 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1713453518
transform 1 0 2308 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1713453518
transform 1 0 2220 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1713453518
transform 1 0 3396 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1713453518
transform 1 0 3348 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1713453518
transform 1 0 3276 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1713453518
transform 1 0 3228 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1713453518
transform 1 0 2476 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1713453518
transform 1 0 2476 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1713453518
transform 1 0 2436 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1713453518
transform 1 0 2340 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1713453518
transform 1 0 3108 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1713453518
transform 1 0 3036 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1713453518
transform 1 0 3036 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1713453518
transform 1 0 2724 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1713453518
transform 1 0 2716 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1713453518
transform 1 0 2508 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1713453518
transform 1 0 2364 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1713453518
transform 1 0 2364 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1713453518
transform 1 0 2252 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1713453518
transform 1 0 2252 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1713453518
transform 1 0 1972 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1713453518
transform 1 0 3244 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1713453518
transform 1 0 3212 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1713453518
transform 1 0 3148 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1713453518
transform 1 0 3108 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1713453518
transform 1 0 3084 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1713453518
transform 1 0 2812 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1713453518
transform 1 0 2156 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1713453518
transform 1 0 2052 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1713453518
transform 1 0 2052 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1713453518
transform 1 0 1980 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1713453518
transform 1 0 1900 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1713453518
transform 1 0 3028 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1713453518
transform 1 0 2932 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1713453518
transform 1 0 3148 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1713453518
transform 1 0 2972 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1713453518
transform 1 0 2964 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1713453518
transform 1 0 2836 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1713453518
transform 1 0 2836 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1713453518
transform 1 0 2604 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1713453518
transform 1 0 2484 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1713453518
transform 1 0 2484 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1713453518
transform 1 0 2380 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1713453518
transform 1 0 1948 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1713453518
transform 1 0 2812 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1713453518
transform 1 0 2628 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1713453518
transform 1 0 2628 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1713453518
transform 1 0 2428 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1713453518
transform 1 0 2428 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1713453518
transform 1 0 1996 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1713453518
transform 1 0 3140 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1713453518
transform 1 0 2964 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1713453518
transform 1 0 2908 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1713453518
transform 1 0 2756 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1713453518
transform 1 0 2748 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1713453518
transform 1 0 2732 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1713453518
transform 1 0 2708 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1713453518
transform 1 0 2708 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1713453518
transform 1 0 2700 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1713453518
transform 1 0 2300 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1713453518
transform 1 0 3012 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1713453518
transform 1 0 2940 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1713453518
transform 1 0 2996 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1713453518
transform 1 0 2932 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1713453518
transform 1 0 2900 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1713453518
transform 1 0 2828 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1713453518
transform 1 0 2780 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1713453518
transform 1 0 2188 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1713453518
transform 1 0 2236 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1713453518
transform 1 0 2004 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1713453518
transform 1 0 1828 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1713453518
transform 1 0 3004 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1713453518
transform 1 0 2988 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1713453518
transform 1 0 2940 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1713453518
transform 1 0 2932 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1713453518
transform 1 0 2932 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1713453518
transform 1 0 2884 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1713453518
transform 1 0 2884 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1713453518
transform 1 0 2844 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1713453518
transform 1 0 2028 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1713453518
transform 1 0 3444 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1713453518
transform 1 0 3404 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1713453518
transform 1 0 3308 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1713453518
transform 1 0 3228 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1713453518
transform 1 0 3180 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1713453518
transform 1 0 3172 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1713453518
transform 1 0 3156 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1713453518
transform 1 0 3156 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1713453518
transform 1 0 3100 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1713453518
transform 1 0 2484 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1713453518
transform 1 0 2444 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1713453518
transform 1 0 2380 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1713453518
transform 1 0 2196 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1713453518
transform 1 0 3276 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1713453518
transform 1 0 3244 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1713453518
transform 1 0 3324 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1713453518
transform 1 0 3292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1713453518
transform 1 0 3292 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1713453518
transform 1 0 3044 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1713453518
transform 1 0 3044 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1713453518
transform 1 0 2668 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1713453518
transform 1 0 2460 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1713453518
transform 1 0 2868 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1713453518
transform 1 0 2620 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1713453518
transform 1 0 2788 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1713453518
transform 1 0 2724 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1713453518
transform 1 0 2196 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1713453518
transform 1 0 2500 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1713453518
transform 1 0 2244 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1713453518
transform 1 0 2244 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1713453518
transform 1 0 2084 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1713453518
transform 1 0 2084 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1713453518
transform 1 0 2004 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1713453518
transform 1 0 3052 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1713453518
transform 1 0 2996 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1713453518
transform 1 0 2988 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1713453518
transform 1 0 2820 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1713453518
transform 1 0 2812 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1713453518
transform 1 0 2644 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1713453518
transform 1 0 2628 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1713453518
transform 1 0 2564 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1713453518
transform 1 0 2532 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1713453518
transform 1 0 2532 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1713453518
transform 1 0 1996 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1713453518
transform 1 0 1996 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1713453518
transform 1 0 1900 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1713453518
transform 1 0 1900 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1713453518
transform 1 0 1844 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1713453518
transform 1 0 244 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1713453518
transform 1 0 220 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1713453518
transform 1 0 300 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1713453518
transform 1 0 284 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1713453518
transform 1 0 252 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1713453518
transform 1 0 212 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1713453518
transform 1 0 428 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1713453518
transform 1 0 388 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1713453518
transform 1 0 260 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1713453518
transform 1 0 220 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1713453518
transform 1 0 260 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1713453518
transform 1 0 220 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1713453518
transform 1 0 220 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1713453518
transform 1 0 148 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1713453518
transform 1 0 324 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1713453518
transform 1 0 284 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1713453518
transform 1 0 476 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1713453518
transform 1 0 356 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1713453518
transform 1 0 260 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1713453518
transform 1 0 228 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1713453518
transform 1 0 196 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1713453518
transform 1 0 92 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1713453518
transform 1 0 220 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1713453518
transform 1 0 116 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1713453518
transform 1 0 148 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1713453518
transform 1 0 116 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1713453518
transform 1 0 380 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1713453518
transform 1 0 308 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1713453518
transform 1 0 324 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1713453518
transform 1 0 292 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1713453518
transform 1 0 932 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1713453518
transform 1 0 860 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1713453518
transform 1 0 812 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1713453518
transform 1 0 676 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1713453518
transform 1 0 676 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1713453518
transform 1 0 588 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1713453518
transform 1 0 468 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1713453518
transform 1 0 1372 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1713453518
transform 1 0 1292 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1713453518
transform 1 0 1292 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1713453518
transform 1 0 996 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1713453518
transform 1 0 884 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1713453518
transform 1 0 820 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1713453518
transform 1 0 740 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1713453518
transform 1 0 700 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1713453518
transform 1 0 636 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1713453518
transform 1 0 580 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1713453518
transform 1 0 556 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1713453518
transform 1 0 2396 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1713453518
transform 1 0 1308 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1713453518
transform 1 0 1308 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1713453518
transform 1 0 1020 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1713453518
transform 1 0 980 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1713453518
transform 1 0 924 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1713453518
transform 1 0 892 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1713453518
transform 1 0 692 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1713453518
transform 1 0 692 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1713453518
transform 1 0 572 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1713453518
transform 1 0 2428 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1713453518
transform 1 0 2364 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1713453518
transform 1 0 2260 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1713453518
transform 1 0 2212 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1713453518
transform 1 0 2076 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1713453518
transform 1 0 2132 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1713453518
transform 1 0 2012 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1713453518
transform 1 0 3100 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1713453518
transform 1 0 2940 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1713453518
transform 1 0 2748 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1713453518
transform 1 0 2636 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1713453518
transform 1 0 2436 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1713453518
transform 1 0 2436 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1713453518
transform 1 0 2012 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1713453518
transform 1 0 2012 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1713453518
transform 1 0 1948 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1713453518
transform 1 0 2276 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1713453518
transform 1 0 1676 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1713453518
transform 1 0 1652 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1713453518
transform 1 0 1540 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1713453518
transform 1 0 1356 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1713453518
transform 1 0 1460 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1713453518
transform 1 0 1396 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1713453518
transform 1 0 3108 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1713453518
transform 1 0 3052 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1713453518
transform 1 0 2932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1713453518
transform 1 0 2932 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1713453518
transform 1 0 2868 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1713453518
transform 1 0 2428 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1713453518
transform 1 0 1956 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1713453518
transform 1 0 412 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1713453518
transform 1 0 380 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1713453518
transform 1 0 3332 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1713453518
transform 1 0 2692 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1713453518
transform 1 0 3148 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1713453518
transform 1 0 2652 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1713453518
transform 1 0 2748 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1713453518
transform 1 0 2516 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1713453518
transform 1 0 3164 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1713453518
transform 1 0 3124 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1713453518
transform 1 0 2700 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1713453518
transform 1 0 2620 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1713453518
transform 1 0 2500 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1713453518
transform 1 0 3012 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1713453518
transform 1 0 2964 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1713453518
transform 1 0 2116 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1713453518
transform 1 0 2076 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1713453518
transform 1 0 2596 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1713453518
transform 1 0 2564 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1713453518
transform 1 0 1324 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1713453518
transform 1 0 1300 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1713453518
transform 1 0 2044 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1713453518
transform 1 0 1908 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1713453518
transform 1 0 1764 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1713453518
transform 1 0 1452 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1713453518
transform 1 0 1396 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1713453518
transform 1 0 1396 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1713453518
transform 1 0 1372 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1713453518
transform 1 0 1740 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1713453518
transform 1 0 1604 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1713453518
transform 1 0 1572 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1713453518
transform 1 0 1516 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1713453518
transform 1 0 2260 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1713453518
transform 1 0 1844 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1713453518
transform 1 0 2020 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1713453518
transform 1 0 1900 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1713453518
transform 1 0 1724 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1713453518
transform 1 0 2260 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1713453518
transform 1 0 2100 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1713453518
transform 1 0 3044 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1713453518
transform 1 0 3004 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1713453518
transform 1 0 1364 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1713453518
transform 1 0 1196 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1713453518
transform 1 0 2428 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1713453518
transform 1 0 1244 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1713453518
transform 1 0 3060 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1713453518
transform 1 0 2908 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1713453518
transform 1 0 2276 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1713453518
transform 1 0 1308 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1713453518
transform 1 0 3412 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1713453518
transform 1 0 3388 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1713453518
transform 1 0 548 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1713453518
transform 1 0 508 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1713453518
transform 1 0 2772 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1713453518
transform 1 0 2684 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1713453518
transform 1 0 2684 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1713453518
transform 1 0 2604 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1713453518
transform 1 0 3076 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1713453518
transform 1 0 3052 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1713453518
transform 1 0 3412 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1713453518
transform 1 0 3388 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1713453518
transform 1 0 2388 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1713453518
transform 1 0 2340 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1713453518
transform 1 0 524 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1713453518
transform 1 0 468 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1713453518
transform 1 0 460 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1713453518
transform 1 0 420 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1713453518
transform 1 0 764 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1713453518
transform 1 0 764 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1713453518
transform 1 0 724 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1713453518
transform 1 0 724 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1713453518
transform 1 0 676 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1713453518
transform 1 0 644 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1713453518
transform 1 0 2788 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1713453518
transform 1 0 2644 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1713453518
transform 1 0 2596 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1713453518
transform 1 0 3412 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1713453518
transform 1 0 3364 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1713453518
transform 1 0 2836 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1713453518
transform 1 0 2772 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1713453518
transform 1 0 2380 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1713453518
transform 1 0 2380 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1713453518
transform 1 0 2156 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1713453518
transform 1 0 3036 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1713453518
transform 1 0 2996 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1713453518
transform 1 0 2956 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1713453518
transform 1 0 2716 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1713453518
transform 1 0 2660 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1713453518
transform 1 0 3012 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1713453518
transform 1 0 2900 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1713453518
transform 1 0 540 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1713453518
transform 1 0 508 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1713453518
transform 1 0 700 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1713453518
transform 1 0 636 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1713453518
transform 1 0 636 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1713453518
transform 1 0 580 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1713453518
transform 1 0 2188 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1713453518
transform 1 0 2060 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1713453518
transform 1 0 2996 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1713453518
transform 1 0 2956 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1713453518
transform 1 0 3412 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1713453518
transform 1 0 3380 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1713453518
transform 1 0 2524 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1713453518
transform 1 0 2492 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1713453518
transform 1 0 3132 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1713453518
transform 1 0 2780 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1713453518
transform 1 0 3076 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1713453518
transform 1 0 2932 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1713453518
transform 1 0 2804 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1713453518
transform 1 0 2660 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1713453518
transform 1 0 2724 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1713453518
transform 1 0 2660 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1713453518
transform 1 0 3156 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1713453518
transform 1 0 3060 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1713453518
transform 1 0 532 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1713453518
transform 1 0 500 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1713453518
transform 1 0 644 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1713453518
transform 1 0 596 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1713453518
transform 1 0 556 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1713453518
transform 1 0 3292 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1713453518
transform 1 0 2724 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1713453518
transform 1 0 2628 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1713453518
transform 1 0 2628 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1713453518
transform 1 0 732 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1713453518
transform 1 0 692 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1713453518
transform 1 0 668 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1713453518
transform 1 0 612 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1713453518
transform 1 0 604 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1713453518
transform 1 0 548 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1713453518
transform 1 0 548 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1713453518
transform 1 0 492 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1713453518
transform 1 0 580 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1713453518
transform 1 0 532 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1713453518
transform 1 0 452 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1713453518
transform 1 0 452 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1713453518
transform 1 0 564 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1713453518
transform 1 0 548 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1713453518
transform 1 0 484 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1713453518
transform 1 0 484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1713453518
transform 1 0 388 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1713453518
transform 1 0 1796 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1713453518
transform 1 0 1780 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1713453518
transform 1 0 2132 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1713453518
transform 1 0 1988 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1713453518
transform 1 0 1956 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1713453518
transform 1 0 1916 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1713453518
transform 1 0 1860 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1713453518
transform 1 0 2052 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1713453518
transform 1 0 2012 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1713453518
transform 1 0 2148 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1713453518
transform 1 0 2052 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1713453518
transform 1 0 2348 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1713453518
transform 1 0 2220 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1713453518
transform 1 0 1300 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1713453518
transform 1 0 1276 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1713453518
transform 1 0 1228 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1713453518
transform 1 0 1012 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1713453518
transform 1 0 1068 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1713453518
transform 1 0 900 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1713453518
transform 1 0 876 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1713453518
transform 1 0 876 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1713453518
transform 1 0 716 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1713453518
transform 1 0 716 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1713453518
transform 1 0 668 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1713453518
transform 1 0 540 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1713453518
transform 1 0 540 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1713453518
transform 1 0 436 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1713453518
transform 1 0 436 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1713453518
transform 1 0 412 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1713453518
transform 1 0 516 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1713453518
transform 1 0 492 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1713453518
transform 1 0 484 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1713453518
transform 1 0 468 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1713453518
transform 1 0 444 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1713453518
transform 1 0 420 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1713453518
transform 1 0 396 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1713453518
transform 1 0 268 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1713453518
transform 1 0 140 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1713453518
transform 1 0 964 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1713453518
transform 1 0 852 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1713453518
transform 1 0 636 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1713453518
transform 1 0 524 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1713453518
transform 1 0 468 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1713453518
transform 1 0 468 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1713453518
transform 1 0 404 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1713453518
transform 1 0 404 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1713453518
transform 1 0 316 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1713453518
transform 1 0 316 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1713453518
transform 1 0 316 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1713453518
transform 1 0 212 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1713453518
transform 1 0 164 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1713453518
transform 1 0 100 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1713453518
transform 1 0 92 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1713453518
transform 1 0 340 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1713453518
transform 1 0 268 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1713453518
transform 1 0 220 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1713453518
transform 1 0 204 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1713453518
transform 1 0 100 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1713453518
transform 1 0 92 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1713453518
transform 1 0 92 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1713453518
transform 1 0 92 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1713453518
transform 1 0 1076 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1713453518
transform 1 0 524 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1713453518
transform 1 0 492 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1713453518
transform 1 0 492 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1713453518
transform 1 0 308 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1713453518
transform 1 0 180 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1713453518
transform 1 0 92 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1713453518
transform 1 0 68 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1713453518
transform 1 0 3364 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1713453518
transform 1 0 3268 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1713453518
transform 1 0 3164 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1713453518
transform 1 0 3164 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1713453518
transform 1 0 3052 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1713453518
transform 1 0 2356 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1713453518
transform 1 0 2356 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1713453518
transform 1 0 2244 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1713453518
transform 1 0 1804 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1713453518
transform 1 0 1692 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1713453518
transform 1 0 1692 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1713453518
transform 1 0 1580 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1713453518
transform 1 0 1332 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1713453518
transform 1 0 260 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1713453518
transform 1 0 220 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1713453518
transform 1 0 116 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1713453518
transform 1 0 1108 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1713453518
transform 1 0 788 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1713453518
transform 1 0 748 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1713453518
transform 1 0 740 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1713453518
transform 1 0 636 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1713453518
transform 1 0 612 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1713453518
transform 1 0 588 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1713453518
transform 1 0 420 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1713453518
transform 1 0 412 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1713453518
transform 1 0 412 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1713453518
transform 1 0 396 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1713453518
transform 1 0 276 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1713453518
transform 1 0 212 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1713453518
transform 1 0 180 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1713453518
transform 1 0 172 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1713453518
transform 1 0 100 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1713453518
transform 1 0 788 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1713453518
transform 1 0 748 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1713453518
transform 1 0 732 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1713453518
transform 1 0 484 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1713453518
transform 1 0 332 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1713453518
transform 1 0 332 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1713453518
transform 1 0 332 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1713453518
transform 1 0 316 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1713453518
transform 1 0 308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1713453518
transform 1 0 284 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1713453518
transform 1 0 260 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1713453518
transform 1 0 820 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1713453518
transform 1 0 820 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1713453518
transform 1 0 804 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1713453518
transform 1 0 724 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1713453518
transform 1 0 700 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1713453518
transform 1 0 692 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1713453518
transform 1 0 396 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1713453518
transform 1 0 380 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1713453518
transform 1 0 372 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1713453518
transform 1 0 372 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1713453518
transform 1 0 324 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1713453518
transform 1 0 324 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1713453518
transform 1 0 308 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1713453518
transform 1 0 284 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1713453518
transform 1 0 196 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1713453518
transform 1 0 188 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1713453518
transform 1 0 948 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1713453518
transform 1 0 948 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1713453518
transform 1 0 948 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1713453518
transform 1 0 924 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1713453518
transform 1 0 908 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1713453518
transform 1 0 908 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1713453518
transform 1 0 868 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1713453518
transform 1 0 852 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1713453518
transform 1 0 844 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1713453518
transform 1 0 836 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1713453518
transform 1 0 836 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1713453518
transform 1 0 828 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1713453518
transform 1 0 748 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1713453518
transform 1 0 996 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1713453518
transform 1 0 956 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1713453518
transform 1 0 956 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1713453518
transform 1 0 948 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1713453518
transform 1 0 924 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1713453518
transform 1 0 916 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1713453518
transform 1 0 916 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1713453518
transform 1 0 868 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1713453518
transform 1 0 3012 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1713453518
transform 1 0 2988 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1713453518
transform 1 0 2932 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1713453518
transform 1 0 2820 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1713453518
transform 1 0 2644 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1713453518
transform 1 0 2492 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1713453518
transform 1 0 2124 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1713453518
transform 1 0 1020 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1713453518
transform 1 0 1004 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1713453518
transform 1 0 996 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1713453518
transform 1 0 940 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1713453518
transform 1 0 932 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1713453518
transform 1 0 924 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1713453518
transform 1 0 892 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1713453518
transform 1 0 884 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1713453518
transform 1 0 876 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1713453518
transform 1 0 844 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1713453518
transform 1 0 836 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1713453518
transform 1 0 804 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1713453518
transform 1 0 796 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1713453518
transform 1 0 796 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1713453518
transform 1 0 796 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1713453518
transform 1 0 748 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1713453518
transform 1 0 748 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1713453518
transform 1 0 308 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1713453518
transform 1 0 292 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1713453518
transform 1 0 900 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1713453518
transform 1 0 804 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1713453518
transform 1 0 804 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1713453518
transform 1 0 732 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1713453518
transform 1 0 796 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1713453518
transform 1 0 748 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1713453518
transform 1 0 980 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1713453518
transform 1 0 948 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1713453518
transform 1 0 812 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1713453518
transform 1 0 804 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1713453518
transform 1 0 780 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1713453518
transform 1 0 780 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1713453518
transform 1 0 780 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1713453518
transform 1 0 772 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1713453518
transform 1 0 772 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1713453518
transform 1 0 772 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1713453518
transform 1 0 764 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1713453518
transform 1 0 764 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1713453518
transform 1 0 708 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1713453518
transform 1 0 708 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1713453518
transform 1 0 964 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1713453518
transform 1 0 948 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1713453518
transform 1 0 940 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1713453518
transform 1 0 932 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1713453518
transform 1 0 924 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1713453518
transform 1 0 908 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1713453518
transform 1 0 908 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1713453518
transform 1 0 908 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1713453518
transform 1 0 876 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1713453518
transform 1 0 876 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1713453518
transform 1 0 836 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1713453518
transform 1 0 812 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1713453518
transform 1 0 700 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1713453518
transform 1 0 668 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1713453518
transform 1 0 900 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1713453518
transform 1 0 900 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1713453518
transform 1 0 884 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1713453518
transform 1 0 884 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1713453518
transform 1 0 884 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1713453518
transform 1 0 852 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1713453518
transform 1 0 852 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1713453518
transform 1 0 852 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1713453518
transform 1 0 836 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1713453518
transform 1 0 836 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1713453518
transform 1 0 836 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1713453518
transform 1 0 804 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1713453518
transform 1 0 780 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1713453518
transform 1 0 836 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1713453518
transform 1 0 796 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1713453518
transform 1 0 900 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1713453518
transform 1 0 876 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1713453518
transform 1 0 876 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1713453518
transform 1 0 844 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1713453518
transform 1 0 772 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1713453518
transform 1 0 772 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1713453518
transform 1 0 996 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1713453518
transform 1 0 948 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1713453518
transform 1 0 948 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1713453518
transform 1 0 940 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1713453518
transform 1 0 924 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1713453518
transform 1 0 916 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1713453518
transform 1 0 916 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1713453518
transform 1 0 916 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1713453518
transform 1 0 900 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1713453518
transform 1 0 900 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1713453518
transform 1 0 892 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1713453518
transform 1 0 884 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1713453518
transform 1 0 876 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1713453518
transform 1 0 868 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1713453518
transform 1 0 868 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1713453518
transform 1 0 852 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1713453518
transform 1 0 852 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1713453518
transform 1 0 828 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1713453518
transform 1 0 820 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1713453518
transform 1 0 812 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1713453518
transform 1 0 796 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1713453518
transform 1 0 940 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1713453518
transform 1 0 932 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1713453518
transform 1 0 932 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1713453518
transform 1 0 908 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1713453518
transform 1 0 892 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1713453518
transform 1 0 860 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1713453518
transform 1 0 836 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1713453518
transform 1 0 836 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1713453518
transform 1 0 828 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1713453518
transform 1 0 796 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1713453518
transform 1 0 788 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1713453518
transform 1 0 788 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1713453518
transform 1 0 780 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1713453518
transform 1 0 780 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1713453518
transform 1 0 748 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1713453518
transform 1 0 748 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1713453518
transform 1 0 748 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1713453518
transform 1 0 732 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1713453518
transform 1 0 716 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1713453518
transform 1 0 572 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1713453518
transform 1 0 444 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1713453518
transform 1 0 396 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1713453518
transform 1 0 324 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1713453518
transform 1 0 324 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1713453518
transform 1 0 308 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1713453518
transform 1 0 300 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1713453518
transform 1 0 300 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1713453518
transform 1 0 300 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1713453518
transform 1 0 284 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1713453518
transform 1 0 276 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1713453518
transform 1 0 276 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1713453518
transform 1 0 268 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1713453518
transform 1 0 204 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1713453518
transform 1 0 124 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1713453518
transform 1 0 124 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1713453518
transform 1 0 676 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1713453518
transform 1 0 620 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1713453518
transform 1 0 612 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1713453518
transform 1 0 556 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1713453518
transform 1 0 532 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1713453518
transform 1 0 532 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1713453518
transform 1 0 524 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1713453518
transform 1 0 524 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1713453518
transform 1 0 516 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1713453518
transform 1 0 516 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1713453518
transform 1 0 492 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1713453518
transform 1 0 484 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1713453518
transform 1 0 484 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1713453518
transform 1 0 476 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1713453518
transform 1 0 476 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1713453518
transform 1 0 476 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1713453518
transform 1 0 476 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1713453518
transform 1 0 468 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1713453518
transform 1 0 460 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1713453518
transform 1 0 452 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1713453518
transform 1 0 452 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1713453518
transform 1 0 452 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1713453518
transform 1 0 444 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1713453518
transform 1 0 444 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1713453518
transform 1 0 436 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1713453518
transform 1 0 420 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1713453518
transform 1 0 404 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1713453518
transform 1 0 236 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1713453518
transform 1 0 220 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1713453518
transform 1 0 404 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1713453518
transform 1 0 396 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1713453518
transform 1 0 348 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1713453518
transform 1 0 332 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1713453518
transform 1 0 324 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1713453518
transform 1 0 252 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1713453518
transform 1 0 252 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1713453518
transform 1 0 244 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1713453518
transform 1 0 236 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1713453518
transform 1 0 228 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1713453518
transform 1 0 212 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1713453518
transform 1 0 204 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1713453518
transform 1 0 148 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1713453518
transform 1 0 140 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1713453518
transform 1 0 2228 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1713453518
transform 1 0 2228 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1713453518
transform 1 0 2188 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1713453518
transform 1 0 2188 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1713453518
transform 1 0 2172 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1713453518
transform 1 0 2140 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1713453518
transform 1 0 2004 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1713453518
transform 1 0 2004 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1713453518
transform 1 0 1932 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1713453518
transform 1 0 1636 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1713453518
transform 1 0 1548 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1713453518
transform 1 0 1508 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1713453518
transform 1 0 2388 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1713453518
transform 1 0 2308 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1713453518
transform 1 0 2276 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1713453518
transform 1 0 2196 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1713453518
transform 1 0 2180 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1713453518
transform 1 0 2180 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1713453518
transform 1 0 2140 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1713453518
transform 1 0 2132 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1713453518
transform 1 0 3372 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1713453518
transform 1 0 3372 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1713453518
transform 1 0 3316 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1713453518
transform 1 0 3236 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1713453518
transform 1 0 3196 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1713453518
transform 1 0 3188 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1713453518
transform 1 0 3188 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1713453518
transform 1 0 3124 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1713453518
transform 1 0 3108 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1713453518
transform 1 0 3108 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1713453518
transform 1 0 3084 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1713453518
transform 1 0 3084 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1713453518
transform 1 0 3084 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1713453518
transform 1 0 3076 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1713453518
transform 1 0 3076 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1713453518
transform 1 0 3068 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1713453518
transform 1 0 2892 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1713453518
transform 1 0 2884 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1713453518
transform 1 0 2868 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1713453518
transform 1 0 2812 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1713453518
transform 1 0 2796 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1713453518
transform 1 0 2796 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1713453518
transform 1 0 2780 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1713453518
transform 1 0 2756 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1713453518
transform 1 0 2732 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1713453518
transform 1 0 2716 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1713453518
transform 1 0 2700 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1713453518
transform 1 0 2684 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1713453518
transform 1 0 2684 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1713453518
transform 1 0 2660 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1713453518
transform 1 0 2660 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1713453518
transform 1 0 2620 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1713453518
transform 1 0 2620 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1713453518
transform 1 0 2260 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1713453518
transform 1 0 2220 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1713453518
transform 1 0 2948 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1713453518
transform 1 0 2932 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1713453518
transform 1 0 2924 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1713453518
transform 1 0 2852 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1713453518
transform 1 0 2780 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1713453518
transform 1 0 2660 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1713453518
transform 1 0 2660 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1713453518
transform 1 0 2604 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1713453518
transform 1 0 2524 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1713453518
transform 1 0 2500 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1713453518
transform 1 0 2500 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1713453518
transform 1 0 2484 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1713453518
transform 1 0 2476 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1713453518
transform 1 0 2468 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1713453518
transform 1 0 2460 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1713453518
transform 1 0 2460 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1713453518
transform 1 0 2452 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1713453518
transform 1 0 2436 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1713453518
transform 1 0 2420 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1713453518
transform 1 0 2420 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1713453518
transform 1 0 2412 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1713453518
transform 1 0 2404 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1713453518
transform 1 0 2356 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1713453518
transform 1 0 2348 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1713453518
transform 1 0 2324 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1713453518
transform 1 0 2300 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1713453518
transform 1 0 2284 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1713453518
transform 1 0 3404 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1713453518
transform 1 0 3396 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1713453518
transform 1 0 3372 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1713453518
transform 1 0 3332 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1713453518
transform 1 0 3332 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1713453518
transform 1 0 3308 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1713453518
transform 1 0 3308 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1713453518
transform 1 0 3300 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1713453518
transform 1 0 3292 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1713453518
transform 1 0 3268 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1713453518
transform 1 0 3084 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1713453518
transform 1 0 2996 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1713453518
transform 1 0 2988 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1713453518
transform 1 0 2988 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1713453518
transform 1 0 2956 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1713453518
transform 1 0 2948 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1713453518
transform 1 0 2892 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1713453518
transform 1 0 2884 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1713453518
transform 1 0 2860 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1713453518
transform 1 0 2828 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1713453518
transform 1 0 3436 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1713453518
transform 1 0 3436 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1713453518
transform 1 0 3428 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1713453518
transform 1 0 3404 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1713453518
transform 1 0 3380 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1713453518
transform 1 0 3372 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1713453518
transform 1 0 3356 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1713453518
transform 1 0 3356 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1713453518
transform 1 0 3324 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1713453518
transform 1 0 3268 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1713453518
transform 1 0 3268 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1713453518
transform 1 0 3164 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1713453518
transform 1 0 3164 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1713453518
transform 1 0 3028 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1713453518
transform 1 0 3428 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1713453518
transform 1 0 3428 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1713453518
transform 1 0 3404 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1713453518
transform 1 0 3404 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1713453518
transform 1 0 3396 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1713453518
transform 1 0 3388 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1713453518
transform 1 0 3388 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1713453518
transform 1 0 3388 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1713453518
transform 1 0 3388 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1713453518
transform 1 0 3372 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1713453518
transform 1 0 3348 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1713453518
transform 1 0 3348 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1713453518
transform 1 0 3348 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1713453518
transform 1 0 3332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1713453518
transform 1 0 3316 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1713453518
transform 1 0 3308 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1713453518
transform 1 0 3308 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1713453518
transform 1 0 3300 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1713453518
transform 1 0 3244 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1713453518
transform 1 0 3244 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1713453518
transform 1 0 3236 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1713453518
transform 1 0 3236 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1713453518
transform 1 0 3100 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1713453518
transform 1 0 3100 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1713453518
transform 1 0 3092 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1713453518
transform 1 0 3092 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1713453518
transform 1 0 3084 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1713453518
transform 1 0 3084 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1713453518
transform 1 0 3044 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1713453518
transform 1 0 3044 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1713453518
transform 1 0 2980 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1713453518
transform 1 0 2940 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1713453518
transform 1 0 2932 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1713453518
transform 1 0 2932 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1713453518
transform 1 0 2916 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1713453518
transform 1 0 2900 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1713453518
transform 1 0 2900 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1713453518
transform 1 0 2804 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1713453518
transform 1 0 2804 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1713453518
transform 1 0 3260 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1713453518
transform 1 0 3252 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1713453518
transform 1 0 3236 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1713453518
transform 1 0 3236 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1713453518
transform 1 0 3236 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1713453518
transform 1 0 3196 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1713453518
transform 1 0 3188 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1713453518
transform 1 0 3172 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1713453518
transform 1 0 3132 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1713453518
transform 1 0 3116 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1713453518
transform 1 0 3108 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1713453518
transform 1 0 3108 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1713453518
transform 1 0 3084 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1713453518
transform 1 0 3084 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1713453518
transform 1 0 3068 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1713453518
transform 1 0 3068 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1713453518
transform 1 0 3068 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1713453518
transform 1 0 3036 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1713453518
transform 1 0 2988 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1713453518
transform 1 0 2980 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1713453518
transform 1 0 2956 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1713453518
transform 1 0 2852 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1713453518
transform 1 0 2820 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1713453518
transform 1 0 2788 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1713453518
transform 1 0 2788 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1713453518
transform 1 0 2740 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1713453518
transform 1 0 2740 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1713453518
transform 1 0 2732 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1713453518
transform 1 0 2732 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1713453518
transform 1 0 2716 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1713453518
transform 1 0 2684 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1713453518
transform 1 0 2676 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1713453518
transform 1 0 2676 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1713453518
transform 1 0 2636 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1713453518
transform 1 0 2636 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1713453518
transform 1 0 2876 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1713453518
transform 1 0 2780 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1713453518
transform 1 0 2580 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1713453518
transform 1 0 2956 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1713453518
transform 1 0 2588 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1713453518
transform 1 0 2580 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1713453518
transform 1 0 2452 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1713453518
transform 1 0 2276 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1713453518
transform 1 0 2596 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1713453518
transform 1 0 2540 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1713453518
transform 1 0 2516 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1713453518
transform 1 0 2420 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1713453518
transform 1 0 2412 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1713453518
transform 1 0 2412 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1713453518
transform 1 0 2380 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1713453518
transform 1 0 2348 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1713453518
transform 1 0 2316 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1713453518
transform 1 0 2308 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1713453518
transform 1 0 2268 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1713453518
transform 1 0 2228 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1713453518
transform 1 0 2212 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1713453518
transform 1 0 2212 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1713453518
transform 1 0 2212 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1713453518
transform 1 0 2204 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1713453518
transform 1 0 2180 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1713453518
transform 1 0 2180 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1713453518
transform 1 0 2180 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1713453518
transform 1 0 2092 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1713453518
transform 1 0 2076 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1713453518
transform 1 0 2076 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1713453518
transform 1 0 2076 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1713453518
transform 1 0 2076 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1713453518
transform 1 0 2020 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1713453518
transform 1 0 2012 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1713453518
transform 1 0 1980 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1713453518
transform 1 0 1964 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1713453518
transform 1 0 1932 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1713453518
transform 1 0 1916 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1713453518
transform 1 0 1892 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1713453518
transform 1 0 1892 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1713453518
transform 1 0 1884 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1713453518
transform 1 0 1884 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1713453518
transform 1 0 1884 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1713453518
transform 1 0 1884 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1713453518
transform 1 0 1860 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1713453518
transform 1 0 1852 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1713453518
transform 1 0 1844 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1713453518
transform 1 0 1828 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1713453518
transform 1 0 1820 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1713453518
transform 1 0 1516 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1713453518
transform 1 0 1508 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1713453518
transform 1 0 1476 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1713453518
transform 1 0 2388 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1713453518
transform 1 0 2308 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1713453518
transform 1 0 2164 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1713453518
transform 1 0 2156 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1713453518
transform 1 0 2140 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1713453518
transform 1 0 2116 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1713453518
transform 1 0 2116 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1713453518
transform 1 0 2060 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1713453518
transform 1 0 2060 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1713453518
transform 1 0 2012 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1713453518
transform 1 0 1972 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1713453518
transform 1 0 1940 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1713453518
transform 1 0 1868 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1713453518
transform 1 0 2188 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1713453518
transform 1 0 2164 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1713453518
transform 1 0 2140 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1713453518
transform 1 0 2132 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1713453518
transform 1 0 2132 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1713453518
transform 1 0 2132 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1713453518
transform 1 0 2100 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1713453518
transform 1 0 2100 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1713453518
transform 1 0 2036 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1713453518
transform 1 0 2036 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1713453518
transform 1 0 2028 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1713453518
transform 1 0 2004 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1713453518
transform 1 0 1932 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1713453518
transform 1 0 1932 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1713453518
transform 1 0 1900 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1713453518
transform 1 0 1892 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1713453518
transform 1 0 1868 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1713453518
transform 1 0 2340 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1713453518
transform 1 0 2252 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1713453518
transform 1 0 2196 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1713453518
transform 1 0 2196 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1713453518
transform 1 0 2124 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1713453518
transform 1 0 2124 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1713453518
transform 1 0 2116 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1713453518
transform 1 0 2084 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1713453518
transform 1 0 2084 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1713453518
transform 1 0 2084 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1713453518
transform 1 0 2076 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1713453518
transform 1 0 1988 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1713453518
transform 1 0 1988 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1713453518
transform 1 0 1988 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1713453518
transform 1 0 1980 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1713453518
transform 1 0 1924 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1713453518
transform 1 0 1908 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1713453518
transform 1 0 2132 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1713453518
transform 1 0 2124 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1713453518
transform 1 0 2116 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1713453518
transform 1 0 2084 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1713453518
transform 1 0 2052 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1713453518
transform 1 0 2052 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1713453518
transform 1 0 2036 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1713453518
transform 1 0 2028 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1713453518
transform 1 0 2012 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1713453518
transform 1 0 2012 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1713453518
transform 1 0 1996 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1713453518
transform 1 0 1964 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1713453518
transform 1 0 1964 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1713453518
transform 1 0 1964 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1713453518
transform 1 0 1964 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1713453518
transform 1 0 1932 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1713453518
transform 1 0 1932 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1713453518
transform 1 0 1892 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1713453518
transform 1 0 1868 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1713453518
transform 1 0 1868 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1713453518
transform 1 0 1868 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1713453518
transform 1 0 1804 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1713453518
transform 1 0 1764 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1713453518
transform 1 0 1764 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1713453518
transform 1 0 1732 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1713453518
transform 1 0 1644 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1713453518
transform 1 0 1540 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1713453518
transform 1 0 2508 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1713453518
transform 1 0 2468 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1713453518
transform 1 0 2404 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1713453518
transform 1 0 2404 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1713453518
transform 1 0 2364 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1713453518
transform 1 0 2228 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1713453518
transform 1 0 2620 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1713453518
transform 1 0 2588 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1713453518
transform 1 0 2540 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1713453518
transform 1 0 2540 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1713453518
transform 1 0 2476 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1713453518
transform 1 0 2476 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1713453518
transform 1 0 2388 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1713453518
transform 1 0 2324 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1713453518
transform 1 0 2324 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1713453518
transform 1 0 2228 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1713453518
transform 1 0 1708 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1713453518
transform 1 0 1660 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1713453518
transform 1 0 1660 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1713453518
transform 1 0 1604 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1713453518
transform 1 0 1604 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1713453518
transform 1 0 1580 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1713453518
transform 1 0 1572 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1713453518
transform 1 0 1572 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1713453518
transform 1 0 1564 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1713453518
transform 1 0 1548 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1713453518
transform 1 0 1524 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1713453518
transform 1 0 1524 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1713453518
transform 1 0 1404 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1713453518
transform 1 0 1372 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1713453518
transform 1 0 1676 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1713453518
transform 1 0 1668 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1713453518
transform 1 0 1524 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1713453518
transform 1 0 1524 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1713453518
transform 1 0 1508 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1713453518
transform 1 0 1500 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1713453518
transform 1 0 1492 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1713453518
transform 1 0 1492 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1713453518
transform 1 0 1372 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1713453518
transform 1 0 1372 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1713453518
transform 1 0 1348 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1713453518
transform 1 0 1348 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1713453518
transform 1 0 1292 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1713453518
transform 1 0 1292 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1713453518
transform 1 0 1716 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1713453518
transform 1 0 1692 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1713453518
transform 1 0 1652 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1713453518
transform 1 0 1588 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1713453518
transform 1 0 1572 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1713453518
transform 1 0 1564 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1713453518
transform 1 0 1556 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1713453518
transform 1 0 1556 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1713453518
transform 1 0 1476 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1713453518
transform 1 0 1468 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1713453518
transform 1 0 1468 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1713453518
transform 1 0 1452 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1713453518
transform 1 0 1420 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1713453518
transform 1 0 1420 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1713453518
transform 1 0 1420 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1713453518
transform 1 0 1420 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1713453518
transform 1 0 1380 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1713453518
transform 1 0 1380 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1713453518
transform 1 0 1692 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1713453518
transform 1 0 1684 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1713453518
transform 1 0 1668 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1713453518
transform 1 0 1652 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1713453518
transform 1 0 1644 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1713453518
transform 1 0 1628 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1713453518
transform 1 0 1628 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1713453518
transform 1 0 1596 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1713453518
transform 1 0 1596 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1713453518
transform 1 0 1572 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1713453518
transform 1 0 1564 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1713453518
transform 1 0 1540 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1713453518
transform 1 0 1540 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1713453518
transform 1 0 1540 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1713453518
transform 1 0 1524 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1713453518
transform 1 0 1500 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1713453518
transform 1 0 1492 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1713453518
transform 1 0 1452 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1713453518
transform 1 0 1444 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1713453518
transform 1 0 1444 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1713453518
transform 1 0 1428 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1713453518
transform 1 0 1412 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1713453518
transform 1 0 1404 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1713453518
transform 1 0 1396 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1713453518
transform 1 0 1388 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1713453518
transform 1 0 1364 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1713453518
transform 1 0 1356 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1713453518
transform 1 0 1316 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1713453518
transform 1 0 1300 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1713453518
transform 1 0 2812 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1713453518
transform 1 0 2412 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1713453518
transform 1 0 1052 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1713453518
transform 1 0 1044 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1713453518
transform 1 0 1044 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1713453518
transform 1 0 1028 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1713453518
transform 1 0 1020 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1713453518
transform 1 0 1004 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1713453518
transform 1 0 988 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1713453518
transform 1 0 900 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1713453518
transform 1 0 1068 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1713453518
transform 1 0 1060 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1713453518
transform 1 0 1060 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1713453518
transform 1 0 1060 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1713453518
transform 1 0 1044 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1713453518
transform 1 0 1012 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1713453518
transform 1 0 1012 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1713453518
transform 1 0 1012 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1713453518
transform 1 0 1004 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1713453518
transform 1 0 1004 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1713453518
transform 1 0 972 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1713453518
transform 1 0 972 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1713453518
transform 1 0 964 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1713453518
transform 1 0 2884 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1713453518
transform 1 0 2820 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1713453518
transform 1 0 2764 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1713453518
transform 1 0 2732 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1713453518
transform 1 0 2428 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1713453518
transform 1 0 2252 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1713453518
transform 1 0 1356 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1713453518
transform 1 0 1060 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1713453518
transform 1 0 1052 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1713453518
transform 1 0 1012 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1713453518
transform 1 0 996 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1713453518
transform 1 0 964 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1713453518
transform 1 0 892 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1713453518
transform 1 0 852 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1713453518
transform 1 0 836 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1713453518
transform 1 0 836 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1713453518
transform 1 0 828 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1713453518
transform 1 0 828 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1713453518
transform 1 0 828 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1713453518
transform 1 0 820 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1713453518
transform 1 0 812 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1713453518
transform 1 0 812 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1713453518
transform 1 0 612 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1713453518
transform 1 0 572 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1713453518
transform 1 0 516 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1713453518
transform 1 0 484 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1713453518
transform 1 0 484 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1713453518
transform 1 0 444 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1713453518
transform 1 0 428 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1713453518
transform 1 0 428 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1713453518
transform 1 0 412 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1713453518
transform 1 0 404 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1713453518
transform 1 0 404 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1713453518
transform 1 0 396 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1713453518
transform 1 0 500 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1713453518
transform 1 0 468 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1713453518
transform 1 0 468 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1713453518
transform 1 0 460 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1713453518
transform 1 0 444 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1713453518
transform 1 0 444 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1713453518
transform 1 0 436 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1713453518
transform 1 0 436 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1713453518
transform 1 0 436 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1713453518
transform 1 0 420 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1713453518
transform 1 0 404 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1713453518
transform 1 0 404 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1713453518
transform 1 0 388 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1713453518
transform 1 0 356 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1713453518
transform 1 0 340 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1713453518
transform 1 0 300 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1713453518
transform 1 0 2732 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1713453518
transform 1 0 2724 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1713453518
transform 1 0 2668 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1713453518
transform 1 0 2636 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1713453518
transform 1 0 2636 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1713453518
transform 1 0 2444 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1713453518
transform 1 0 2300 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1713453518
transform 1 0 2268 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1713453518
transform 1 0 2268 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1713453518
transform 1 0 2260 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1713453518
transform 1 0 2260 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1713453518
transform 1 0 2180 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1713453518
transform 1 0 2172 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1713453518
transform 1 0 2116 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1713453518
transform 1 0 1892 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1713453518
transform 1 0 1644 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1713453518
transform 1 0 3428 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1713453518
transform 1 0 3388 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1713453518
transform 1 0 3364 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1713453518
transform 1 0 3364 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1713453518
transform 1 0 3324 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1713453518
transform 1 0 3324 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1713453518
transform 1 0 3268 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1713453518
transform 1 0 3220 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1713453518
transform 1 0 3148 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1713453518
transform 1 0 1788 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1713453518
transform 1 0 1788 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1713453518
transform 1 0 1780 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1713453518
transform 1 0 1780 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1713453518
transform 1 0 1764 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1713453518
transform 1 0 1764 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1713453518
transform 1 0 1732 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1713453518
transform 1 0 1724 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1713453518
transform 1 0 1716 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1713453518
transform 1 0 1716 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1713453518
transform 1 0 1700 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1713453518
transform 1 0 1556 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1713453518
transform 1 0 1548 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1713453518
transform 1 0 1444 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1713453518
transform 1 0 1492 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1713453518
transform 1 0 1444 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1713453518
transform 1 0 1436 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1713453518
transform 1 0 1428 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1713453518
transform 1 0 1412 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1713453518
transform 1 0 1388 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1713453518
transform 1 0 1356 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1713453518
transform 1 0 1332 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1713453518
transform 1 0 1332 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1713453518
transform 1 0 1316 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1713453518
transform 1 0 1316 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1713453518
transform 1 0 1316 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1713453518
transform 1 0 1316 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1713453518
transform 1 0 1268 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1713453518
transform 1 0 1268 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1713453518
transform 1 0 1228 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1713453518
transform 1 0 1228 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1713453518
transform 1 0 1228 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1713453518
transform 1 0 1212 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1713453518
transform 1 0 1188 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1713453518
transform 1 0 1188 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1713453518
transform 1 0 1172 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1713453518
transform 1 0 1172 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1713453518
transform 1 0 1156 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1713453518
transform 1 0 1156 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1713453518
transform 1 0 1124 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1713453518
transform 1 0 1516 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1713453518
transform 1 0 1508 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1713453518
transform 1 0 1500 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1713453518
transform 1 0 1484 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1713453518
transform 1 0 1484 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1713453518
transform 1 0 1468 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1713453518
transform 1 0 1460 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1713453518
transform 1 0 1452 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1713453518
transform 1 0 1452 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1713453518
transform 1 0 1436 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1713453518
transform 1 0 1428 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1713453518
transform 1 0 1428 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1713453518
transform 1 0 1388 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1713453518
transform 1 0 1348 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1713453518
transform 1 0 1348 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1713453518
transform 1 0 1348 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1713453518
transform 1 0 1300 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1713453518
transform 1 0 1244 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1713453518
transform 1 0 1196 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1713453518
transform 1 0 2892 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1713453518
transform 1 0 2828 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1713453518
transform 1 0 2764 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1713453518
transform 1 0 2668 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1713453518
transform 1 0 2492 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1713453518
transform 1 0 2492 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1713453518
transform 1 0 2420 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1713453518
transform 1 0 2404 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1713453518
transform 1 0 2404 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1713453518
transform 1 0 2388 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1713453518
transform 1 0 2300 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1713453518
transform 1 0 2228 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1713453518
transform 1 0 1404 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1713453518
transform 1 0 1404 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1713453518
transform 1 0 1356 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1713453518
transform 1 0 1332 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1713453518
transform 1 0 1324 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1713453518
transform 1 0 1268 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1713453518
transform 1 0 1220 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1713453518
transform 1 0 1108 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1713453518
transform 1 0 3356 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1713453518
transform 1 0 3324 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1713453518
transform 1 0 3300 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1713453518
transform 1 0 3284 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1713453518
transform 1 0 3244 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1713453518
transform 1 0 3244 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1713453518
transform 1 0 2780 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1713453518
transform 1 0 2716 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1713453518
transform 1 0 2668 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1713453518
transform 1 0 2668 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1713453518
transform 1 0 2668 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1713453518
transform 1 0 2580 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1713453518
transform 1 0 2548 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1713453518
transform 1 0 2540 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1713453518
transform 1 0 2460 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1713453518
transform 1 0 2420 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1713453518
transform 1 0 1812 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1713453518
transform 1 0 3420 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1713453518
transform 1 0 3412 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1713453518
transform 1 0 3196 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1713453518
transform 1 0 3188 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1713453518
transform 1 0 3012 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1713453518
transform 1 0 2748 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1713453518
transform 1 0 2740 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1713453518
transform 1 0 2588 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1713453518
transform 1 0 2588 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1713453518
transform 1 0 2508 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1713453518
transform 1 0 2508 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1713453518
transform 1 0 2484 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1713453518
transform 1 0 2484 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1713453518
transform 1 0 2388 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1713453518
transform 1 0 2388 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1713453518
transform 1 0 1868 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1713453518
transform 1 0 3404 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1713453518
transform 1 0 3180 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1713453518
transform 1 0 3172 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1713453518
transform 1 0 2900 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1713453518
transform 1 0 2900 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1713453518
transform 1 0 2796 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1713453518
transform 1 0 2756 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1713453518
transform 1 0 2716 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1713453518
transform 1 0 2612 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1713453518
transform 1 0 2604 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1713453518
transform 1 0 2604 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1713453518
transform 1 0 2572 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1713453518
transform 1 0 2476 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1713453518
transform 1 0 2452 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1713453518
transform 1 0 2740 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1713453518
transform 1 0 2628 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1713453518
transform 1 0 2572 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1713453518
transform 1 0 2228 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1713453518
transform 1 0 1988 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1713453518
transform 1 0 1988 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1713453518
transform 1 0 1132 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1713453518
transform 1 0 1124 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1713453518
transform 1 0 1108 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1713453518
transform 1 0 1076 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1713453518
transform 1 0 1068 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1713453518
transform 1 0 1052 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1713453518
transform 1 0 1020 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1713453518
transform 1 0 2956 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1713453518
transform 1 0 2956 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1713453518
transform 1 0 2916 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1713453518
transform 1 0 2916 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1713453518
transform 1 0 2860 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1713453518
transform 1 0 2852 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1713453518
transform 1 0 2852 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1713453518
transform 1 0 2652 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1713453518
transform 1 0 2492 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1713453518
transform 1 0 2492 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1713453518
transform 1 0 2492 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1713453518
transform 1 0 2212 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1713453518
transform 1 0 3332 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1713453518
transform 1 0 3220 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1713453518
transform 1 0 3220 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1713453518
transform 1 0 3204 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1713453518
transform 1 0 3084 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1713453518
transform 1 0 2916 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1713453518
transform 1 0 2916 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1713453518
transform 1 0 2828 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1713453518
transform 1 0 2644 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1713453518
transform 1 0 2612 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1713453518
transform 1 0 2612 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1713453518
transform 1 0 2612 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1713453518
transform 1 0 2572 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1713453518
transform 1 0 2540 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1713453518
transform 1 0 2444 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1713453518
transform 1 0 1700 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1713453518
transform 1 0 3404 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1713453518
transform 1 0 3332 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1713453518
transform 1 0 3332 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1713453518
transform 1 0 3292 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1713453518
transform 1 0 3180 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1713453518
transform 1 0 2996 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1713453518
transform 1 0 2996 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1713453518
transform 1 0 2980 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1713453518
transform 1 0 2980 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1713453518
transform 1 0 2948 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1713453518
transform 1 0 2948 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1713453518
transform 1 0 2932 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1713453518
transform 1 0 2700 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1713453518
transform 1 0 2684 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1713453518
transform 1 0 2660 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1713453518
transform 1 0 2652 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1713453518
transform 1 0 2468 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1713453518
transform 1 0 1836 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1713453518
transform 1 0 3276 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1713453518
transform 1 0 3140 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1713453518
transform 1 0 3044 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1713453518
transform 1 0 3012 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1713453518
transform 1 0 2948 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1713453518
transform 1 0 2764 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1713453518
transform 1 0 2764 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1713453518
transform 1 0 2572 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1713453518
transform 1 0 2572 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1713453518
transform 1 0 2572 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1713453518
transform 1 0 2524 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1713453518
transform 1 0 2380 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1713453518
transform 1 0 2380 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1713453518
transform 1 0 1652 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1713453518
transform 1 0 3140 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1713453518
transform 1 0 3076 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1713453518
transform 1 0 2956 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1713453518
transform 1 0 2956 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1713453518
transform 1 0 2892 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1713453518
transform 1 0 2796 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1713453518
transform 1 0 2692 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1713453518
transform 1 0 2580 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1713453518
transform 1 0 2580 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1713453518
transform 1 0 2420 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1713453518
transform 1 0 2412 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1713453518
transform 1 0 2140 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1713453518
transform 1 0 2140 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1713453518
transform 1 0 1876 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1713453518
transform 1 0 1300 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1713453518
transform 1 0 2836 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1713453518
transform 1 0 2772 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1713453518
transform 1 0 2684 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1713453518
transform 1 0 2556 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1713453518
transform 1 0 2260 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1713453518
transform 1 0 2260 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1713453518
transform 1 0 2172 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1713453518
transform 1 0 2172 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1713453518
transform 1 0 1588 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1713453518
transform 1 0 1588 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1713453518
transform 1 0 1236 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1713453518
transform 1 0 1236 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1713453518
transform 1 0 1188 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1713453518
transform 1 0 1148 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1713453518
transform 1 0 1076 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1713453518
transform 1 0 1020 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1713453518
transform 1 0 3124 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1713453518
transform 1 0 3076 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1713453518
transform 1 0 3044 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1713453518
transform 1 0 3004 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1713453518
transform 1 0 3004 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1713453518
transform 1 0 2724 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1713453518
transform 1 0 2436 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1713453518
transform 1 0 2292 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1713453518
transform 1 0 2292 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1713453518
transform 1 0 1948 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1713453518
transform 1 0 1948 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1713453518
transform 1 0 1732 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1713453518
transform 1 0 1644 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1713453518
transform 1 0 1524 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1713453518
transform 1 0 2556 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1713453518
transform 1 0 2308 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1713453518
transform 1 0 2308 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1713453518
transform 1 0 2020 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1713453518
transform 1 0 2020 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1713453518
transform 1 0 1428 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1713453518
transform 1 0 1580 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1713453518
transform 1 0 1532 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1713453518
transform 1 0 1516 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1713453518
transform 1 0 1500 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1713453518
transform 1 0 1500 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1713453518
transform 1 0 1324 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1713453518
transform 1 0 1292 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1713453518
transform 1 0 2796 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1713453518
transform 1 0 2716 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1713453518
transform 1 0 3100 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1713453518
transform 1 0 3068 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1713453518
transform 1 0 2980 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1713453518
transform 1 0 2980 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1713453518
transform 1 0 2436 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1713453518
transform 1 0 2084 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1713453518
transform 1 0 3148 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1713453518
transform 1 0 3036 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1713453518
transform 1 0 2828 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1713453518
transform 1 0 2828 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1713453518
transform 1 0 2828 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1713453518
transform 1 0 2740 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1713453518
transform 1 0 2676 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1713453518
transform 1 0 2676 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1713453518
transform 1 0 2300 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1713453518
transform 1 0 3100 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1713453518
transform 1 0 3036 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1713453518
transform 1 0 3036 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1713453518
transform 1 0 2940 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1713453518
transform 1 0 2892 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1713453518
transform 1 0 2892 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1713453518
transform 1 0 2860 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1713453518
transform 1 0 2860 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1713453518
transform 1 0 2860 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1713453518
transform 1 0 2668 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1713453518
transform 1 0 2380 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1713453518
transform 1 0 2380 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1713453518
transform 1 0 2324 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1713453518
transform 1 0 3212 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1713453518
transform 1 0 3156 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1713453518
transform 1 0 2876 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1713453518
transform 1 0 2484 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1713453518
transform 1 0 2356 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1713453518
transform 1 0 2356 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1713453518
transform 1 0 2204 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1713453518
transform 1 0 2156 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1713453518
transform 1 0 3372 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1713453518
transform 1 0 3348 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1713453518
transform 1 0 3332 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1713453518
transform 1 0 3324 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1713453518
transform 1 0 3324 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1713453518
transform 1 0 3076 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1713453518
transform 1 0 2228 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1713453518
transform 1 0 2196 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1713453518
transform 1 0 2188 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1713453518
transform 1 0 3284 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1713453518
transform 1 0 3284 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1713453518
transform 1 0 3276 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1713453518
transform 1 0 3220 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1713453518
transform 1 0 3220 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1713453518
transform 1 0 2804 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1713453518
transform 1 0 2644 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1713453518
transform 1 0 2180 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1713453518
transform 1 0 3452 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1713453518
transform 1 0 3452 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1713453518
transform 1 0 3420 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1713453518
transform 1 0 3412 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1713453518
transform 1 0 3300 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1713453518
transform 1 0 3188 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1713453518
transform 1 0 2908 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1713453518
transform 1 0 2196 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1713453518
transform 1 0 3364 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1713453518
transform 1 0 3364 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1713453518
transform 1 0 3324 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1713453518
transform 1 0 3260 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1713453518
transform 1 0 3252 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1713453518
transform 1 0 3020 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1713453518
transform 1 0 2236 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1713453518
transform 1 0 2172 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1713453518
transform 1 0 2164 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1713453518
transform 1 0 2156 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1713453518
transform 1 0 2068 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1713453518
transform 1 0 2044 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1713453518
transform 1 0 2020 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1713453518
transform 1 0 1644 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1713453518
transform 1 0 1380 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1713453518
transform 1 0 1316 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1713453518
transform 1 0 1284 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1713453518
transform 1 0 1284 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1713453518
transform 1 0 1284 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1713453518
transform 1 0 1276 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1713453518
transform 1 0 1276 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1713453518
transform 1 0 1236 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1713453518
transform 1 0 1236 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1713453518
transform 1 0 1220 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1713453518
transform 1 0 1220 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1713453518
transform 1 0 1220 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1713453518
transform 1 0 1204 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1713453518
transform 1 0 1204 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1713453518
transform 1 0 1180 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1713453518
transform 1 0 1124 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1713453518
transform 1 0 1076 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1713453518
transform 1 0 1404 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1713453518
transform 1 0 1380 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1713453518
transform 1 0 1372 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1713453518
transform 1 0 1372 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1713453518
transform 1 0 1356 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1713453518
transform 1 0 1284 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1713453518
transform 1 0 1268 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1713453518
transform 1 0 1228 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1713453518
transform 1 0 1180 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1713453518
transform 1 0 1172 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1713453518
transform 1 0 1140 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1713453518
transform 1 0 1124 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1713453518
transform 1 0 1916 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1713453518
transform 1 0 1916 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1713453518
transform 1 0 1884 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1713453518
transform 1 0 1876 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1713453518
transform 1 0 1844 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1713453518
transform 1 0 1820 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1713453518
transform 1 0 1492 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1713453518
transform 1 0 3356 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1713453518
transform 1 0 3356 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1713453518
transform 1 0 3188 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1713453518
transform 1 0 3188 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1713453518
transform 1 0 2676 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1713453518
transform 1 0 2180 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1713453518
transform 1 0 1556 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1713453518
transform 1 0 1516 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1713453518
transform 1 0 1452 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1713453518
transform 1 0 1452 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1713453518
transform 1 0 1388 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1713453518
transform 1 0 1388 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1713453518
transform 1 0 1332 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1713453518
transform 1 0 1308 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1713453518
transform 1 0 1276 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1713453518
transform 1 0 1212 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1713453518
transform 1 0 1204 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1713453518
transform 1 0 1204 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1713453518
transform 1 0 1196 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1713453518
transform 1 0 1188 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1713453518
transform 1 0 1172 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1713453518
transform 1 0 1140 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1713453518
transform 1 0 1116 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1713453518
transform 1 0 1108 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1713453518
transform 1 0 2044 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1713453518
transform 1 0 1948 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1713453518
transform 1 0 1844 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1713453518
transform 1 0 1972 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1713453518
transform 1 0 1852 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1713453518
transform 1 0 1724 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1713453518
transform 1 0 2740 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1713453518
transform 1 0 2700 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1713453518
transform 1 0 2724 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1713453518
transform 1 0 2660 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1713453518
transform 1 0 3044 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1713453518
transform 1 0 2948 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1713453518
transform 1 0 3388 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1713453518
transform 1 0 3140 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1713453518
transform 1 0 3076 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1713453518
transform 1 0 2708 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1713453518
transform 1 0 3292 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1713453518
transform 1 0 2788 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1713453518
transform 1 0 3316 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1713453518
transform 1 0 3020 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1713453518
transform 1 0 3420 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1713453518
transform 1 0 3252 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1713453518
transform 1 0 3452 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1713453518
transform 1 0 3452 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1713453518
transform 1 0 3412 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1713453518
transform 1 0 3388 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1713453518
transform 1 0 3324 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1713453518
transform 1 0 3284 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1713453518
transform 1 0 3204 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1713453518
transform 1 0 2836 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1713453518
transform 1 0 3316 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1713453518
transform 1 0 3300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1713453518
transform 1 0 3300 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1713453518
transform 1 0 3212 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1713453518
transform 1 0 3412 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1713453518
transform 1 0 3412 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1713453518
transform 1 0 3372 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1713453518
transform 1 0 3316 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1713453518
transform 1 0 3196 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1713453518
transform 1 0 3148 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1713453518
transform 1 0 3148 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1713453518
transform 1 0 3028 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1713453518
transform 1 0 3028 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1713453518
transform 1 0 2804 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1713453518
transform 1 0 3244 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1713453518
transform 1 0 3172 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1713453518
transform 1 0 3132 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1713453518
transform 1 0 3020 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1713453518
transform 1 0 3348 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1713453518
transform 1 0 3188 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1713453518
transform 1 0 3084 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1713453518
transform 1 0 3012 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1713453518
transform 1 0 2924 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1713453518
transform 1 0 2868 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1713453518
transform 1 0 2780 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1713453518
transform 1 0 2692 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1713453518
transform 1 0 2956 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1713453518
transform 1 0 2868 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1713453518
transform 1 0 3036 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1713453518
transform 1 0 2948 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1713453518
transform 1 0 2268 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1713453518
transform 1 0 2172 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1713453518
transform 1 0 2516 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1713453518
transform 1 0 2444 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1713453518
transform 1 0 884 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1713453518
transform 1 0 796 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1713453518
transform 1 0 1028 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1713453518
transform 1 0 956 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1713453518
transform 1 0 1084 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1713453518
transform 1 0 988 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1713453518
transform 1 0 1044 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1713453518
transform 1 0 964 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1713453518
transform 1 0 980 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1713453518
transform 1 0 900 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1713453518
transform 1 0 1036 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1713453518
transform 1 0 956 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1713453518
transform 1 0 1044 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1713453518
transform 1 0 940 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1713453518
transform 1 0 1020 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1713453518
transform 1 0 900 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1713453518
transform 1 0 1092 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1713453518
transform 1 0 964 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1713453518
transform 1 0 988 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1713453518
transform 1 0 876 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1713453518
transform 1 0 1084 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1713453518
transform 1 0 988 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1713453518
transform 1 0 1012 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1713453518
transform 1 0 916 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1713453518
transform 1 0 1052 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1713453518
transform 1 0 956 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1713453518
transform 1 0 1028 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1713453518
transform 1 0 1004 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1713453518
transform 1 0 1084 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1713453518
transform 1 0 1004 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1713453518
transform 1 0 1084 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1713453518
transform 1 0 964 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1713453518
transform 1 0 1044 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1713453518
transform 1 0 956 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1713453518
transform 1 0 1028 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1713453518
transform 1 0 940 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1713453518
transform 1 0 1012 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1713453518
transform 1 0 916 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1713453518
transform 1 0 1068 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1713453518
transform 1 0 972 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1713453518
transform 1 0 1092 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1713453518
transform 1 0 996 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1713453518
transform 1 0 1044 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1713453518
transform 1 0 948 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1713453518
transform 1 0 1052 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1713453518
transform 1 0 964 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1713453518
transform 1 0 1092 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1713453518
transform 1 0 1004 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1713453518
transform 1 0 1068 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1713453518
transform 1 0 996 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1713453518
transform 1 0 1124 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1713453518
transform 1 0 1036 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1713453518
transform 1 0 1140 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1713453518
transform 1 0 1068 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1713453518
transform 1 0 1100 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1713453518
transform 1 0 956 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1713453518
transform 1 0 1068 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1713453518
transform 1 0 940 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1713453518
transform 1 0 908 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1713453518
transform 1 0 844 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1713453518
transform 1 0 892 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1713453518
transform 1 0 796 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1713453518
transform 1 0 916 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1713453518
transform 1 0 852 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1713453518
transform 1 0 1052 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1713453518
transform 1 0 852 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1713453518
transform 1 0 3068 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1713453518
transform 1 0 3020 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1713453518
transform 1 0 2220 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1713453518
transform 1 0 2172 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1713453518
transform 1 0 2172 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1713453518
transform 1 0 2156 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1713453518
transform 1 0 3100 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1713453518
transform 1 0 3004 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1713453518
transform 1 0 2732 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1713453518
transform 1 0 2636 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1713453518
transform 1 0 2468 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1713453518
transform 1 0 2068 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1713453518
transform 1 0 1924 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1713453518
transform 1 0 1804 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1713453518
transform 1 0 1796 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1713453518
transform 1 0 1740 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1713453518
transform 1 0 1620 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1713453518
transform 1 0 1532 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1713453518
transform 1 0 1524 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1713453518
transform 1 0 1468 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1713453518
transform 1 0 636 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1713453518
transform 1 0 420 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1713453518
transform 1 0 404 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1713453518
transform 1 0 348 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1713453518
transform 1 0 212 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1713453518
transform 1 0 196 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1713453518
transform 1 0 2028 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1713453518
transform 1 0 1748 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1713453518
transform 1 0 1708 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1713453518
transform 1 0 1068 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1713453518
transform 1 0 1068 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1713453518
transform 1 0 1044 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2584
timestamp 1713453518
transform 1 0 2988 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1713453518
transform 1 0 1988 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1713453518
transform 1 0 2084 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1713453518
transform 1 0 1996 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1713453518
transform 1 0 2012 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1713453518
transform 1 0 1964 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1713453518
transform 1 0 2252 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1713453518
transform 1 0 2052 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1713453518
transform 1 0 2316 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1713453518
transform 1 0 2244 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1713453518
transform 1 0 2692 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1713453518
transform 1 0 2340 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1713453518
transform 1 0 2716 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1713453518
transform 1 0 2652 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1713453518
transform 1 0 2660 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2599
timestamp 1713453518
transform 1 0 2452 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1713453518
transform 1 0 2452 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1713453518
transform 1 0 2332 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1713453518
transform 1 0 3028 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1713453518
transform 1 0 2740 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1713453518
transform 1 0 2652 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1713453518
transform 1 0 1988 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1713453518
transform 1 0 2060 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1713453518
transform 1 0 1956 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1713453518
transform 1 0 1916 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1713453518
transform 1 0 1940 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1713453518
transform 1 0 1692 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1713453518
transform 1 0 1636 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1713453518
transform 1 0 1332 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1713453518
transform 1 0 3244 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1713453518
transform 1 0 3204 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1713453518
transform 1 0 3204 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1713453518
transform 1 0 3196 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1713453518
transform 1 0 3188 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1713453518
transform 1 0 3188 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1713453518
transform 1 0 3164 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1713453518
transform 1 0 3164 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1713453518
transform 1 0 2772 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1713453518
transform 1 0 2684 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1713453518
transform 1 0 2684 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1713453518
transform 1 0 2588 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1713453518
transform 1 0 2476 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1713453518
transform 1 0 1748 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1713453518
transform 1 0 1692 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1713453518
transform 1 0 1564 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1713453518
transform 1 0 1564 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1713453518
transform 1 0 1404 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1713453518
transform 1 0 2348 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1713453518
transform 1 0 2236 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1713453518
transform 1 0 1724 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1713453518
transform 1 0 1684 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1713453518
transform 1 0 1412 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1713453518
transform 1 0 2932 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1713453518
transform 1 0 2724 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1713453518
transform 1 0 2692 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1713453518
transform 1 0 2684 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1713453518
transform 1 0 2956 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1713453518
transform 1 0 2932 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1713453518
transform 1 0 3076 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1713453518
transform 1 0 2948 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1713453518
transform 1 0 2948 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1713453518
transform 1 0 2660 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1713453518
transform 1 0 1580 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1713453518
transform 1 0 3260 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1713453518
transform 1 0 3204 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1713453518
transform 1 0 3148 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1713453518
transform 1 0 3148 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1713453518
transform 1 0 3012 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1713453518
transform 1 0 3012 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1713453518
transform 1 0 2972 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1713453518
transform 1 0 2948 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1713453518
transform 1 0 2900 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1713453518
transform 1 0 2900 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1713453518
transform 1 0 2836 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1713453518
transform 1 0 2836 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1713453518
transform 1 0 2812 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1713453518
transform 1 0 2812 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1713453518
transform 1 0 2580 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1713453518
transform 1 0 2356 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1713453518
transform 1 0 1748 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1713453518
transform 1 0 2988 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1713453518
transform 1 0 2612 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1713453518
transform 1 0 2588 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1713453518
transform 1 0 1692 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1713453518
transform 1 0 2716 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1713453518
transform 1 0 2628 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1713453518
transform 1 0 2308 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1713453518
transform 1 0 1812 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1713453518
transform 1 0 2652 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1713453518
transform 1 0 2572 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1713453518
transform 1 0 2276 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1713453518
transform 1 0 2276 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1713453518
transform 1 0 1884 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1713453518
transform 1 0 2676 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1713453518
transform 1 0 2660 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1713453518
transform 1 0 2660 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1713453518
transform 1 0 2572 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1713453518
transform 1 0 2276 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1713453518
transform 1 0 2204 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1713453518
transform 1 0 2636 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1713453518
transform 1 0 2604 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1713453518
transform 1 0 2612 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1713453518
transform 1 0 2572 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1713453518
transform 1 0 2884 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1713453518
transform 1 0 2796 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1713453518
transform 1 0 3396 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1713453518
transform 1 0 3380 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1713453518
transform 1 0 3244 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1713453518
transform 1 0 3204 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1713453518
transform 1 0 2852 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1713453518
transform 1 0 2844 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1713453518
transform 1 0 2836 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1713453518
transform 1 0 2788 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1713453518
transform 1 0 2780 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1713453518
transform 1 0 2780 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1713453518
transform 1 0 2676 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1713453518
transform 1 0 2580 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1713453518
transform 1 0 2564 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1713453518
transform 1 0 2548 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1713453518
transform 1 0 1908 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1713453518
transform 1 0 2972 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1713453518
transform 1 0 2860 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1713453518
transform 1 0 2716 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1713453518
transform 1 0 2684 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1713453518
transform 1 0 2972 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1713453518
transform 1 0 2892 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1713453518
transform 1 0 2804 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1713453518
transform 1 0 2764 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1713453518
transform 1 0 2780 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1713453518
transform 1 0 2428 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1713453518
transform 1 0 1836 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1713453518
transform 1 0 2356 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1713453518
transform 1 0 2276 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1713453518
transform 1 0 2532 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2718
timestamp 1713453518
transform 1 0 2388 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1713453518
transform 1 0 2476 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1713453518
transform 1 0 2436 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1713453518
transform 1 0 2668 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1713453518
transform 1 0 2388 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1713453518
transform 1 0 2524 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1713453518
transform 1 0 2412 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1713453518
transform 1 0 2388 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1713453518
transform 1 0 2188 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1713453518
transform 1 0 2164 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1713453518
transform 1 0 2116 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1713453518
transform 1 0 2220 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1713453518
transform 1 0 2124 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1713453518
transform 1 0 2164 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1713453518
transform 1 0 2052 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1713453518
transform 1 0 2892 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1713453518
transform 1 0 2188 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1713453518
transform 1 0 2148 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1713453518
transform 1 0 2036 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1713453518
transform 1 0 2036 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1713453518
transform 1 0 1820 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1713453518
transform 1 0 2644 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1713453518
transform 1 0 2484 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1713453518
transform 1 0 2252 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1713453518
transform 1 0 3244 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2743
timestamp 1713453518
transform 1 0 3228 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1713453518
transform 1 0 3180 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1713453518
transform 1 0 3172 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1713453518
transform 1 0 3172 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1713453518
transform 1 0 3036 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1713453518
transform 1 0 2812 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1713453518
transform 1 0 2748 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1713453518
transform 1 0 2748 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1713453518
transform 1 0 2228 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1713453518
transform 1 0 1996 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1713453518
transform 1 0 3044 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1713453518
transform 1 0 3012 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1713453518
transform 1 0 2508 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1713453518
transform 1 0 2028 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2757
timestamp 1713453518
transform 1 0 2012 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1713453518
transform 1 0 1924 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1713453518
transform 1 0 1916 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1713453518
transform 1 0 1868 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1713453518
transform 1 0 1852 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1713453518
transform 1 0 1828 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2763
timestamp 1713453518
transform 1 0 1924 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1713453518
transform 1 0 1788 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1713453518
transform 1 0 1596 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1713453518
transform 1 0 3260 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2767
timestamp 1713453518
transform 1 0 3236 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1713453518
transform 1 0 3180 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1713453518
transform 1 0 3108 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1713453518
transform 1 0 2532 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1713453518
transform 1 0 2500 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1713453518
transform 1 0 2308 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1713453518
transform 1 0 2292 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1713453518
transform 1 0 2292 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1713453518
transform 1 0 1932 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1713453518
transform 1 0 2972 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1713453518
transform 1 0 2556 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1713453518
transform 1 0 2540 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1713453518
transform 1 0 2404 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1713453518
transform 1 0 2604 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1713453518
transform 1 0 2564 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1713453518
transform 1 0 3276 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1713453518
transform 1 0 3236 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1713453518
transform 1 0 2884 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1713453518
transform 1 0 2604 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1713453518
transform 1 0 2372 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1713453518
transform 1 0 2348 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1713453518
transform 1 0 2340 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1713453518
transform 1 0 2740 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1713453518
transform 1 0 2676 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1713453518
transform 1 0 3316 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1713453518
transform 1 0 3284 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1713453518
transform 1 0 3284 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1713453518
transform 1 0 3284 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1713453518
transform 1 0 3268 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1713453518
transform 1 0 3236 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1713453518
transform 1 0 2828 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1713453518
transform 1 0 2828 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1713453518
transform 1 0 2684 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1713453518
transform 1 0 2364 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1713453518
transform 1 0 2356 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1713453518
transform 1 0 2132 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1713453518
transform 1 0 2116 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1713453518
transform 1 0 2036 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1713453518
transform 1 0 2548 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1713453518
transform 1 0 2508 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2807
timestamp 1713453518
transform 1 0 3260 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1713453518
transform 1 0 3132 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1713453518
transform 1 0 3004 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1713453518
transform 1 0 3004 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1713453518
transform 1 0 3004 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1713453518
transform 1 0 2948 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1713453518
transform 1 0 2948 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1713453518
transform 1 0 2692 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1713453518
transform 1 0 2692 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2816
timestamp 1713453518
transform 1 0 2516 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1713453518
transform 1 0 2516 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1713453518
transform 1 0 1924 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1713453518
transform 1 0 2540 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1713453518
transform 1 0 2412 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1713453518
transform 1 0 2364 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1713453518
transform 1 0 2308 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1713453518
transform 1 0 2452 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1713453518
transform 1 0 2316 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1713453518
transform 1 0 2860 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1713453518
transform 1 0 2860 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2827
timestamp 1713453518
transform 1 0 2788 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2828
timestamp 1713453518
transform 1 0 2652 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1713453518
transform 1 0 2484 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1713453518
transform 1 0 2484 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1713453518
transform 1 0 2436 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1713453518
transform 1 0 2620 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1713453518
transform 1 0 2548 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1713453518
transform 1 0 2548 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1713453518
transform 1 0 2332 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2836
timestamp 1713453518
transform 1 0 2332 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1713453518
transform 1 0 2308 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1713453518
transform 1 0 2196 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1713453518
transform 1 0 2172 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2840
timestamp 1713453518
transform 1 0 2156 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1713453518
transform 1 0 2684 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1713453518
transform 1 0 2596 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1713453518
transform 1 0 2884 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1713453518
transform 1 0 2692 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1713453518
transform 1 0 2492 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2846
timestamp 1713453518
transform 1 0 2132 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1713453518
transform 1 0 2676 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1713453518
transform 1 0 2532 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1713453518
transform 1 0 2892 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1713453518
transform 1 0 2756 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1713453518
transform 1 0 2676 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1713453518
transform 1 0 2620 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1713453518
transform 1 0 2620 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1713453518
transform 1 0 1796 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1713453518
transform 1 0 2564 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1713453518
transform 1 0 2420 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1713453518
transform 1 0 2340 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1713453518
transform 1 0 2252 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1713453518
transform 1 0 2220 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1713453518
transform 1 0 2196 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1713453518
transform 1 0 2188 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1713453518
transform 1 0 2084 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1713453518
transform 1 0 2308 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1713453518
transform 1 0 2300 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1713453518
transform 1 0 2292 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1713453518
transform 1 0 2252 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1713453518
transform 1 0 2428 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1713453518
transform 1 0 2204 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1713453518
transform 1 0 2148 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1713453518
transform 1 0 2148 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2871
timestamp 1713453518
transform 1 0 2148 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1713453518
transform 1 0 2100 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2873
timestamp 1713453518
transform 1 0 2100 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1713453518
transform 1 0 2444 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1713453518
transform 1 0 2332 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2876
timestamp 1713453518
transform 1 0 2252 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1713453518
transform 1 0 2500 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1713453518
transform 1 0 2492 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1713453518
transform 1 0 2412 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1713453518
transform 1 0 2388 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1713453518
transform 1 0 2276 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1713453518
transform 1 0 1916 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1713453518
transform 1 0 1892 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1713453518
transform 1 0 1860 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1713453518
transform 1 0 1852 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1713453518
transform 1 0 1836 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1713453518
transform 1 0 2332 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1713453518
transform 1 0 2260 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1713453518
transform 1 0 2340 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1713453518
transform 1 0 2300 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1713453518
transform 1 0 2548 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1713453518
transform 1 0 2500 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1713453518
transform 1 0 2444 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1713453518
transform 1 0 2252 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1713453518
transform 1 0 2364 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1713453518
transform 1 0 2300 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1713453518
transform 1 0 2564 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1713453518
transform 1 0 2452 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1713453518
transform 1 0 2404 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1713453518
transform 1 0 2308 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1713453518
transform 1 0 2308 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1713453518
transform 1 0 2204 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1713453518
transform 1 0 2372 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1713453518
transform 1 0 2340 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1713453518
transform 1 0 2548 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1713453518
transform 1 0 2524 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1713453518
transform 1 0 2444 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1713453518
transform 1 0 2324 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1713453518
transform 1 0 2268 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1713453518
transform 1 0 2316 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1713453518
transform 1 0 2276 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1713453518
transform 1 0 2588 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1713453518
transform 1 0 2484 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1713453518
transform 1 0 2356 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1713453518
transform 1 0 2140 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1713453518
transform 1 0 1932 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1713453518
transform 1 0 2404 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1713453518
transform 1 0 2356 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1713453518
transform 1 0 2948 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1713453518
transform 1 0 2948 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1713453518
transform 1 0 2916 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1713453518
transform 1 0 2796 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1713453518
transform 1 0 2796 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1713453518
transform 1 0 2524 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1713453518
transform 1 0 2380 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1713453518
transform 1 0 2060 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1713453518
transform 1 0 2036 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1713453518
transform 1 0 2444 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1713453518
transform 1 0 2404 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1713453518
transform 1 0 2572 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1713453518
transform 1 0 2468 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1713453518
transform 1 0 2428 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1713453518
transform 1 0 2116 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1713453518
transform 1 0 2116 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1713453518
transform 1 0 2084 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1713453518
transform 1 0 2076 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1713453518
transform 1 0 2540 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1713453518
transform 1 0 2508 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1713453518
transform 1 0 2484 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1713453518
transform 1 0 1732 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1713453518
transform 1 0 1612 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1713453518
transform 1 0 1788 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1713453518
transform 1 0 1652 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1713453518
transform 1 0 2340 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1713453518
transform 1 0 2244 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1713453518
transform 1 0 2188 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1713453518
transform 1 0 2012 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1713453518
transform 1 0 2340 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1713453518
transform 1 0 2284 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1713453518
transform 1 0 2284 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1713453518
transform 1 0 2252 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1713453518
transform 1 0 2900 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1713453518
transform 1 0 2860 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1713453518
transform 1 0 2836 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1713453518
transform 1 0 2828 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2956
timestamp 1713453518
transform 1 0 2476 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1713453518
transform 1 0 2276 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1713453518
transform 1 0 2116 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1713453518
transform 1 0 2116 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1713453518
transform 1 0 2060 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2961
timestamp 1713453518
transform 1 0 2060 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1713453518
transform 1 0 2020 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2963
timestamp 1713453518
transform 1 0 2388 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1713453518
transform 1 0 2356 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1713453518
transform 1 0 2012 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1713453518
transform 1 0 1972 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1713453518
transform 1 0 2028 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1713453518
transform 1 0 1948 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1713453518
transform 1 0 1988 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1713453518
transform 1 0 1948 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1713453518
transform 1 0 2252 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1713453518
transform 1 0 2028 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2973
timestamp 1713453518
transform 1 0 2068 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1713453518
transform 1 0 2044 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1713453518
transform 1 0 2020 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1713453518
transform 1 0 1980 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1713453518
transform 1 0 2068 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1713453518
transform 1 0 2060 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1713453518
transform 1 0 2044 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1713453518
transform 1 0 2028 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1713453518
transform 1 0 1948 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1713453518
transform 1 0 1852 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1713453518
transform 1 0 2052 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1713453518
transform 1 0 1852 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1713453518
transform 1 0 1484 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1713453518
transform 1 0 2348 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1713453518
transform 1 0 2244 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1713453518
transform 1 0 2340 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1713453518
transform 1 0 2284 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1713453518
transform 1 0 2260 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1713453518
transform 1 0 1924 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1713453518
transform 1 0 1716 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1713453518
transform 1 0 2372 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1713453518
transform 1 0 2116 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2995
timestamp 1713453518
transform 1 0 2092 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2996
timestamp 1713453518
transform 1 0 2052 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2997
timestamp 1713453518
transform 1 0 2156 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1713453518
transform 1 0 2012 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1713453518
transform 1 0 1884 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1713453518
transform 1 0 2356 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1713453518
transform 1 0 2172 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1713453518
transform 1 0 2388 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1713453518
transform 1 0 2348 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1713453518
transform 1 0 2468 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1713453518
transform 1 0 2364 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1713453518
transform 1 0 2132 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1713453518
transform 1 0 1852 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1713453518
transform 1 0 1812 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3009
timestamp 1713453518
transform 1 0 2004 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1713453518
transform 1 0 1972 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1713453518
transform 1 0 1852 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1713453518
transform 1 0 2028 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3013
timestamp 1713453518
transform 1 0 1988 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1713453518
transform 1 0 1996 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1713453518
transform 1 0 1948 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1713453518
transform 1 0 2084 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1713453518
transform 1 0 2012 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1713453518
transform 1 0 2252 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3019
timestamp 1713453518
transform 1 0 2100 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1713453518
transform 1 0 2060 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1713453518
transform 1 0 2100 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1713453518
transform 1 0 1964 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1713453518
transform 1 0 2060 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3024
timestamp 1713453518
transform 1 0 1876 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1713453518
transform 1 0 1900 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1713453518
transform 1 0 1740 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1713453518
transform 1 0 1748 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1713453518
transform 1 0 1668 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1713453518
transform 1 0 1740 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1713453518
transform 1 0 1660 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3031
timestamp 1713453518
transform 1 0 2212 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1713453518
transform 1 0 1988 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1713453518
transform 1 0 1820 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1713453518
transform 1 0 2084 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1713453518
transform 1 0 2076 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1713453518
transform 1 0 1988 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1713453518
transform 1 0 1988 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1713453518
transform 1 0 2116 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1713453518
transform 1 0 2092 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3040
timestamp 1713453518
transform 1 0 2092 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1713453518
transform 1 0 1924 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1713453518
transform 1 0 1948 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1713453518
transform 1 0 1876 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1713453518
transform 1 0 1868 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1713453518
transform 1 0 1828 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1713453518
transform 1 0 1820 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1713453518
transform 1 0 1796 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1713453518
transform 1 0 2124 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3049
timestamp 1713453518
transform 1 0 2076 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1713453518
transform 1 0 1988 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3051
timestamp 1713453518
transform 1 0 2196 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1713453518
transform 1 0 2132 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1713453518
transform 1 0 2100 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1713453518
transform 1 0 1940 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1713453518
transform 1 0 1892 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1713453518
transform 1 0 2148 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1713453518
transform 1 0 1908 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1713453518
transform 1 0 2228 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1713453518
transform 1 0 2132 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1713453518
transform 1 0 2412 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1713453518
transform 1 0 2060 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1713453518
transform 1 0 2076 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1713453518
transform 1 0 1556 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1713453518
transform 1 0 1540 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1713453518
transform 1 0 1500 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1713453518
transform 1 0 1252 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1713453518
transform 1 0 1548 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1713453518
transform 1 0 1444 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1713453518
transform 1 0 2396 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1713453518
transform 1 0 2316 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1713453518
transform 1 0 2940 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1713453518
transform 1 0 2444 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1713453518
transform 1 0 2932 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1713453518
transform 1 0 2860 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1713453518
transform 1 0 2796 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1713453518
transform 1 0 2324 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1713453518
transform 1 0 1228 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1713453518
transform 1 0 2948 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1713453518
transform 1 0 2708 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1713453518
transform 1 0 2644 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1713453518
transform 1 0 2644 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1713453518
transform 1 0 2396 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1713453518
transform 1 0 2396 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1713453518
transform 1 0 1196 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1713453518
transform 1 0 2220 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1713453518
transform 1 0 2100 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1713453518
transform 1 0 2100 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1713453518
transform 1 0 1308 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1713453518
transform 1 0 1260 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1713453518
transform 1 0 2324 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1713453518
transform 1 0 1932 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1713453518
transform 1 0 1932 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1713453518
transform 1 0 1540 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1713453518
transform 1 0 1540 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1713453518
transform 1 0 1356 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1713453518
transform 1 0 2316 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1713453518
transform 1 0 2132 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1713453518
transform 1 0 2212 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1713453518
transform 1 0 2140 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1713453518
transform 1 0 2172 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1713453518
transform 1 0 2012 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1713453518
transform 1 0 1820 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1713453518
transform 1 0 1788 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1713453518
transform 1 0 1660 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1713453518
transform 1 0 1148 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1713453518
transform 1 0 2276 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1713453518
transform 1 0 2100 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1713453518
transform 1 0 1740 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1713453518
transform 1 0 1660 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1713453518
transform 1 0 1660 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1713453518
transform 1 0 1612 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1713453518
transform 1 0 2252 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1713453518
transform 1 0 2220 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1713453518
transform 1 0 2156 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1713453518
transform 1 0 1460 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1713453518
transform 1 0 2788 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1713453518
transform 1 0 2660 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1713453518
transform 1 0 2420 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1713453518
transform 1 0 2420 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1713453518
transform 1 0 2332 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1713453518
transform 1 0 1964 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1713453518
transform 1 0 1964 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1713453518
transform 1 0 1692 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1713453518
transform 1 0 2188 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1713453518
transform 1 0 2148 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1713453518
transform 1 0 1532 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1713453518
transform 1 0 2100 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1713453518
transform 1 0 2004 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1713453518
transform 1 0 1548 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1713453518
transform 1 0 1292 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1713453518
transform 1 0 2180 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1713453518
transform 1 0 2076 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1713453518
transform 1 0 2076 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1713453518
transform 1 0 1932 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1713453518
transform 1 0 1524 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1713453518
transform 1 0 1404 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1713453518
transform 1 0 1132 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1713453518
transform 1 0 2084 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1713453518
transform 1 0 1980 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3140
timestamp 1713453518
transform 1 0 2092 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1713453518
transform 1 0 2036 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1713453518
transform 1 0 1196 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1713453518
transform 1 0 3364 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1713453518
transform 1 0 3332 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1713453518
transform 1 0 3332 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1713453518
transform 1 0 3180 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1713453518
transform 1 0 3172 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1713453518
transform 1 0 3116 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1713453518
transform 1 0 2892 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1713453518
transform 1 0 2884 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1713453518
transform 1 0 2572 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1713453518
transform 1 0 2556 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1713453518
transform 1 0 2556 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1713453518
transform 1 0 2532 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1713453518
transform 1 0 2532 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1713453518
transform 1 0 2484 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1713453518
transform 1 0 2476 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1713453518
transform 1 0 2436 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1713453518
transform 1 0 2028 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1713453518
transform 1 0 1908 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1713453518
transform 1 0 2172 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1713453518
transform 1 0 2140 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1713453518
transform 1 0 2052 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1713453518
transform 1 0 1708 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1713453518
transform 1 0 1596 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3166
timestamp 1713453518
transform 1 0 1260 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1713453518
transform 1 0 2156 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1713453518
transform 1 0 1788 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1713453518
transform 1 0 1788 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1713453518
transform 1 0 1724 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1713453518
transform 1 0 1428 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1713453518
transform 1 0 1428 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3173
timestamp 1713453518
transform 1 0 1340 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1713453518
transform 1 0 2196 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1713453518
transform 1 0 2124 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1713453518
transform 1 0 2180 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1713453518
transform 1 0 2156 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1713453518
transform 1 0 2236 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1713453518
transform 1 0 2196 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3180
timestamp 1713453518
transform 1 0 2188 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1713453518
transform 1 0 2132 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1713453518
transform 1 0 1924 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1713453518
transform 1 0 1924 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1713453518
transform 1 0 1524 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1713453518
transform 1 0 2228 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3186
timestamp 1713453518
transform 1 0 2020 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1713453518
transform 1 0 1684 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1713453518
transform 1 0 1644 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1713453518
transform 1 0 1564 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1713453518
transform 1 0 1516 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1713453518
transform 1 0 2124 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1713453518
transform 1 0 1708 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1713453518
transform 1 0 1708 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3194
timestamp 1713453518
transform 1 0 1684 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1713453518
transform 1 0 1452 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1713453518
transform 1 0 2204 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3197
timestamp 1713453518
transform 1 0 1708 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1713453518
transform 1 0 1500 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1713453518
transform 1 0 2156 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1713453518
transform 1 0 1884 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1713453518
transform 1 0 1732 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1713453518
transform 1 0 1340 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1713453518
transform 1 0 2140 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1713453518
transform 1 0 1932 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1713453518
transform 1 0 1924 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3206
timestamp 1713453518
transform 1 0 1748 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1713453518
transform 1 0 1684 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1713453518
transform 1 0 1300 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1713453518
transform 1 0 1868 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1713453518
transform 1 0 1764 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1713453518
transform 1 0 1532 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1713453518
transform 1 0 1340 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1713453518
transform 1 0 1964 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1713453518
transform 1 0 1900 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1713453518
transform 1 0 2604 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1713453518
transform 1 0 2532 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1713453518
transform 1 0 2012 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1713453518
transform 1 0 1948 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3219
timestamp 1713453518
transform 1 0 1924 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3220
timestamp 1713453518
transform 1 0 1580 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3221
timestamp 1713453518
transform 1 0 2540 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1713453518
transform 1 0 2508 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3223
timestamp 1713453518
transform 1 0 2348 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1713453518
transform 1 0 2348 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1713453518
transform 1 0 2156 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1713453518
transform 1 0 2116 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1713453518
transform 1 0 1972 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3228
timestamp 1713453518
transform 1 0 1628 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1713453518
transform 1 0 1836 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1713453518
transform 1 0 1812 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1713453518
transform 1 0 1604 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1713453518
transform 1 0 1460 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1713453518
transform 1 0 2092 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3234
timestamp 1713453518
transform 1 0 1892 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3235
timestamp 1713453518
transform 1 0 1892 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1713453518
transform 1 0 1740 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1713453518
transform 1 0 1676 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3238
timestamp 1713453518
transform 1 0 1428 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1713453518
transform 1 0 2932 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3240
timestamp 1713453518
transform 1 0 2836 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3241
timestamp 1713453518
transform 1 0 3092 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1713453518
transform 1 0 2972 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1713453518
transform 1 0 3052 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3244
timestamp 1713453518
transform 1 0 2980 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1713453518
transform 1 0 3436 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1713453518
transform 1 0 3100 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3247
timestamp 1713453518
transform 1 0 3444 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3248
timestamp 1713453518
transform 1 0 3356 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1713453518
transform 1 0 3412 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1713453518
transform 1 0 3396 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1713453518
transform 1 0 3404 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1713453518
transform 1 0 3068 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1713453518
transform 1 0 3364 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1713453518
transform 1 0 3244 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1713453518
transform 1 0 3404 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1713453518
transform 1 0 3388 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1713453518
transform 1 0 3364 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1713453518
transform 1 0 3348 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1713453518
transform 1 0 3324 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1713453518
transform 1 0 3324 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1713453518
transform 1 0 2852 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1713453518
transform 1 0 2780 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1713453518
transform 1 0 2764 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1713453518
transform 1 0 2684 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3265
timestamp 1713453518
transform 1 0 2420 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1713453518
transform 1 0 2372 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1713453518
transform 1 0 2308 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1713453518
transform 1 0 2060 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1713453518
transform 1 0 2060 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1713453518
transform 1 0 1844 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1713453518
transform 1 0 3404 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1713453518
transform 1 0 3340 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1713453518
transform 1 0 3412 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1713453518
transform 1 0 3356 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1713453518
transform 1 0 3316 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1713453518
transform 1 0 3292 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1713453518
transform 1 0 3292 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1713453518
transform 1 0 3212 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1713453518
transform 1 0 3188 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1713453518
transform 1 0 3188 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1713453518
transform 1 0 3164 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1713453518
transform 1 0 3100 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1713453518
transform 1 0 3100 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1713453518
transform 1 0 2860 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1713453518
transform 1 0 2812 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1713453518
transform 1 0 2796 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1713453518
transform 1 0 2604 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1713453518
transform 1 0 2420 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1713453518
transform 1 0 2380 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3290
timestamp 1713453518
transform 1 0 2380 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1713453518
transform 1 0 2356 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3292
timestamp 1713453518
transform 1 0 2356 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1713453518
transform 1 0 2292 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1713453518
transform 1 0 2292 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1713453518
transform 1 0 2268 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1713453518
transform 1 0 1796 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1713453518
transform 1 0 3196 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1713453518
transform 1 0 3164 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1713453518
transform 1 0 3188 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1713453518
transform 1 0 3156 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1713453518
transform 1 0 3180 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3302
timestamp 1713453518
transform 1 0 2892 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1713453518
transform 1 0 2860 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1713453518
transform 1 0 2980 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3305
timestamp 1713453518
transform 1 0 2876 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3306
timestamp 1713453518
transform 1 0 2916 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1713453518
transform 1 0 2892 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1713453518
transform 1 0 2940 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3309
timestamp 1713453518
transform 1 0 2876 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1713453518
transform 1 0 2916 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1713453518
transform 1 0 2804 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1713453518
transform 1 0 3164 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3313
timestamp 1713453518
transform 1 0 3068 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3314
timestamp 1713453518
transform 1 0 3068 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3315
timestamp 1713453518
transform 1 0 3052 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3316
timestamp 1713453518
transform 1 0 2996 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1713453518
transform 1 0 2876 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3318
timestamp 1713453518
transform 1 0 2876 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1713453518
transform 1 0 3044 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3320
timestamp 1713453518
transform 1 0 3020 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3321
timestamp 1713453518
transform 1 0 2988 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3322
timestamp 1713453518
transform 1 0 2876 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3323
timestamp 1713453518
transform 1 0 2772 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3324
timestamp 1713453518
transform 1 0 3420 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1713453518
transform 1 0 3204 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1713453518
transform 1 0 3228 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3327
timestamp 1713453518
transform 1 0 3156 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1713453518
transform 1 0 3140 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1713453518
transform 1 0 3140 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3330
timestamp 1713453518
transform 1 0 3132 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3331
timestamp 1713453518
transform 1 0 3092 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3332
timestamp 1713453518
transform 1 0 2812 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3333
timestamp 1713453518
transform 1 0 2756 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3334
timestamp 1713453518
transform 1 0 2692 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1713453518
transform 1 0 2500 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3336
timestamp 1713453518
transform 1 0 2404 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3337
timestamp 1713453518
transform 1 0 2404 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_3338
timestamp 1713453518
transform 1 0 1772 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3339
timestamp 1713453518
transform 1 0 3172 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1713453518
transform 1 0 3068 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3341
timestamp 1713453518
transform 1 0 3084 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1713453518
transform 1 0 2948 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3343
timestamp 1713453518
transform 1 0 2908 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1713453518
transform 1 0 3028 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3345
timestamp 1713453518
transform 1 0 2988 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3346
timestamp 1713453518
transform 1 0 3396 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1713453518
transform 1 0 3316 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1713453518
transform 1 0 3340 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1713453518
transform 1 0 3300 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1713453518
transform 1 0 3340 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3351
timestamp 1713453518
transform 1 0 3316 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_3352
timestamp 1713453518
transform 1 0 3420 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1713453518
transform 1 0 3356 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3354
timestamp 1713453518
transform 1 0 3436 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3355
timestamp 1713453518
transform 1 0 3396 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1713453518
transform 1 0 2404 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1713453518
transform 1 0 3364 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1713453518
transform 1 0 3292 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1713453518
transform 1 0 3292 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_3360
timestamp 1713453518
transform 1 0 3212 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1713453518
transform 1 0 3420 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1713453518
transform 1 0 3372 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3363
timestamp 1713453518
transform 1 0 3380 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1713453518
transform 1 0 3340 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1713453518
transform 1 0 3332 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3366
timestamp 1713453518
transform 1 0 3316 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1713453518
transform 1 0 3404 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3368
timestamp 1713453518
transform 1 0 3316 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3369
timestamp 1713453518
transform 1 0 2964 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1713453518
transform 1 0 2540 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3371
timestamp 1713453518
transform 1 0 2940 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1713453518
transform 1 0 2916 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1713453518
transform 1 0 2940 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1713453518
transform 1 0 2796 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3375
timestamp 1713453518
transform 1 0 2500 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1713453518
transform 1 0 2500 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3377
timestamp 1713453518
transform 1 0 2004 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3378
timestamp 1713453518
transform 1 0 3292 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3379
timestamp 1713453518
transform 1 0 2980 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3380
timestamp 1713453518
transform 1 0 3244 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3381
timestamp 1713453518
transform 1 0 3236 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3382
timestamp 1713453518
transform 1 0 3220 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3383
timestamp 1713453518
transform 1 0 3220 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3384
timestamp 1713453518
transform 1 0 3292 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_3385
timestamp 1713453518
transform 1 0 3220 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_3386
timestamp 1713453518
transform 1 0 3252 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3387
timestamp 1713453518
transform 1 0 3140 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1713453518
transform 1 0 3028 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3389
timestamp 1713453518
transform 1 0 2924 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1713453518
transform 1 0 2924 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3391
timestamp 1713453518
transform 1 0 2916 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1713453518
transform 1 0 2908 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1713453518
transform 1 0 2876 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3394
timestamp 1713453518
transform 1 0 2876 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_3395
timestamp 1713453518
transform 1 0 2908 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3396
timestamp 1713453518
transform 1 0 2852 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3397
timestamp 1713453518
transform 1 0 2852 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3398
timestamp 1713453518
transform 1 0 2772 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3399
timestamp 1713453518
transform 1 0 3052 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3400
timestamp 1713453518
transform 1 0 2932 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3401
timestamp 1713453518
transform 1 0 3196 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3402
timestamp 1713453518
transform 1 0 3068 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1713453518
transform 1 0 3116 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3404
timestamp 1713453518
transform 1 0 3060 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3405
timestamp 1713453518
transform 1 0 3196 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3406
timestamp 1713453518
transform 1 0 3108 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3407
timestamp 1713453518
transform 1 0 3180 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3408
timestamp 1713453518
transform 1 0 3148 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3409
timestamp 1713453518
transform 1 0 3164 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3410
timestamp 1713453518
transform 1 0 2868 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_3411
timestamp 1713453518
transform 1 0 2836 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3412
timestamp 1713453518
transform 1 0 2772 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3413
timestamp 1713453518
transform 1 0 2748 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1713453518
transform 1 0 2716 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3415
timestamp 1713453518
transform 1 0 2684 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3416
timestamp 1713453518
transform 1 0 2636 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1713453518
transform 1 0 2636 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3418
timestamp 1713453518
transform 1 0 2548 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3419
timestamp 1713453518
transform 1 0 2548 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_3420
timestamp 1713453518
transform 1 0 2436 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3421
timestamp 1713453518
transform 1 0 2436 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1713453518
transform 1 0 2020 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1713453518
transform 1 0 2812 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3424
timestamp 1713453518
transform 1 0 2788 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3425
timestamp 1713453518
transform 1 0 2748 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3426
timestamp 1713453518
transform 1 0 2772 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3427
timestamp 1713453518
transform 1 0 2684 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3428
timestamp 1713453518
transform 1 0 2604 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3429
timestamp 1713453518
transform 1 0 2596 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1713453518
transform 1 0 2580 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3431
timestamp 1713453518
transform 1 0 2556 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3432
timestamp 1713453518
transform 1 0 2212 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3433
timestamp 1713453518
transform 1 0 3372 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1713453518
transform 1 0 3220 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3435
timestamp 1713453518
transform 1 0 2492 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1713453518
transform 1 0 2692 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3437
timestamp 1713453518
transform 1 0 2556 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3438
timestamp 1713453518
transform 1 0 3044 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1713453518
transform 1 0 2868 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1713453518
transform 1 0 2780 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3441
timestamp 1713453518
transform 1 0 2692 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1713453518
transform 1 0 2604 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3443
timestamp 1713453518
transform 1 0 2732 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1713453518
transform 1 0 2652 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3445
timestamp 1713453518
transform 1 0 2572 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3446
timestamp 1713453518
transform 1 0 2636 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1713453518
transform 1 0 2564 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3448
timestamp 1713453518
transform 1 0 3220 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1713453518
transform 1 0 2604 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3450
timestamp 1713453518
transform 1 0 2948 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3451
timestamp 1713453518
transform 1 0 2916 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1713453518
transform 1 0 2916 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3453
timestamp 1713453518
transform 1 0 2860 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1713453518
transform 1 0 3036 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1713453518
transform 1 0 2852 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1713453518
transform 1 0 2836 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3457
timestamp 1713453518
transform 1 0 2852 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3458
timestamp 1713453518
transform 1 0 2780 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1713453518
transform 1 0 2716 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1713453518
transform 1 0 2620 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1713453518
transform 1 0 2612 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3462
timestamp 1713453518
transform 1 0 2100 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1713453518
transform 1 0 3092 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1713453518
transform 1 0 2972 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3465
timestamp 1713453518
transform 1 0 2892 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1713453518
transform 1 0 3196 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1713453518
transform 1 0 2996 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1713453518
transform 1 0 2956 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3469
timestamp 1713453518
transform 1 0 2884 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1713453518
transform 1 0 2852 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3471
timestamp 1713453518
transform 1 0 2820 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3472
timestamp 1713453518
transform 1 0 2724 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1713453518
transform 1 0 3036 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3474
timestamp 1713453518
transform 1 0 2964 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1713453518
transform 1 0 3148 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3476
timestamp 1713453518
transform 1 0 3100 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3477
timestamp 1713453518
transform 1 0 3396 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1713453518
transform 1 0 3052 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3479
timestamp 1713453518
transform 1 0 3116 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3480
timestamp 1713453518
transform 1 0 3116 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3481
timestamp 1713453518
transform 1 0 3084 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3482
timestamp 1713453518
transform 1 0 2964 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3483
timestamp 1713453518
transform 1 0 2956 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1713453518
transform 1 0 2748 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3485
timestamp 1713453518
transform 1 0 3412 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1713453518
transform 1 0 3388 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3487
timestamp 1713453518
transform 1 0 3452 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3488
timestamp 1713453518
transform 1 0 3420 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3489
timestamp 1713453518
transform 1 0 3452 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1713453518
transform 1 0 3420 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3491
timestamp 1713453518
transform 1 0 3412 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3492
timestamp 1713453518
transform 1 0 2932 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3493
timestamp 1713453518
transform 1 0 3020 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_3494
timestamp 1713453518
transform 1 0 2916 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_3495
timestamp 1713453518
transform 1 0 2996 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3496
timestamp 1713453518
transform 1 0 2932 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3497
timestamp 1713453518
transform 1 0 2892 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3498
timestamp 1713453518
transform 1 0 3428 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1713453518
transform 1 0 3372 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1713453518
transform 1 0 3420 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3501
timestamp 1713453518
transform 1 0 3324 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3502
timestamp 1713453518
transform 1 0 3420 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_3503
timestamp 1713453518
transform 1 0 3388 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_3504
timestamp 1713453518
transform 1 0 3364 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_3505
timestamp 1713453518
transform 1 0 3292 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_3506
timestamp 1713453518
transform 1 0 3196 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_3507
timestamp 1713453518
transform 1 0 3396 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_3508
timestamp 1713453518
transform 1 0 3356 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1713453518
transform 1 0 3332 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3510
timestamp 1713453518
transform 1 0 3300 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3511
timestamp 1713453518
transform 1 0 3404 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3512
timestamp 1713453518
transform 1 0 3364 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1713453518
transform 1 0 3340 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1713453518
transform 1 0 3396 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3515
timestamp 1713453518
transform 1 0 3316 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3516
timestamp 1713453518
transform 1 0 3292 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1713453518
transform 1 0 3260 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3518
timestamp 1713453518
transform 1 0 2180 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3519
timestamp 1713453518
transform 1 0 2060 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3520
timestamp 1713453518
transform 1 0 2756 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_3521
timestamp 1713453518
transform 1 0 2100 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_3522
timestamp 1713453518
transform 1 0 1340 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_3523
timestamp 1713453518
transform 1 0 3164 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3524
timestamp 1713453518
transform 1 0 3044 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3525
timestamp 1713453518
transform 1 0 3332 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1713453518
transform 1 0 3060 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3527
timestamp 1713453518
transform 1 0 3436 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3528
timestamp 1713453518
transform 1 0 3364 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1713453518
transform 1 0 3436 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3530
timestamp 1713453518
transform 1 0 3380 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1713453518
transform 1 0 3372 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3532
timestamp 1713453518
transform 1 0 3300 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3533
timestamp 1713453518
transform 1 0 3388 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3534
timestamp 1713453518
transform 1 0 3356 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3535
timestamp 1713453518
transform 1 0 3324 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3536
timestamp 1713453518
transform 1 0 3420 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3537
timestamp 1713453518
transform 1 0 3324 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3538
timestamp 1713453518
transform 1 0 3292 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3539
timestamp 1713453518
transform 1 0 2884 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3540
timestamp 1713453518
transform 1 0 2956 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3541
timestamp 1713453518
transform 1 0 2876 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1713453518
transform 1 0 2972 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3543
timestamp 1713453518
transform 1 0 2892 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3544
timestamp 1713453518
transform 1 0 2836 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1713453518
transform 1 0 3268 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1713453518
transform 1 0 3236 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3547
timestamp 1713453518
transform 1 0 3044 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3548
timestamp 1713453518
transform 1 0 2980 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3549
timestamp 1713453518
transform 1 0 3052 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3550
timestamp 1713453518
transform 1 0 2828 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3551
timestamp 1713453518
transform 1 0 2828 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3552
timestamp 1713453518
transform 1 0 2812 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1713453518
transform 1 0 2788 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3554
timestamp 1713453518
transform 1 0 2972 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3555
timestamp 1713453518
transform 1 0 2916 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3556
timestamp 1713453518
transform 1 0 3068 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1713453518
transform 1 0 2988 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3558
timestamp 1713453518
transform 1 0 3084 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3559
timestamp 1713453518
transform 1 0 2932 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3560
timestamp 1713453518
transform 1 0 3012 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1713453518
transform 1 0 2964 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1713453518
transform 1 0 2860 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3563
timestamp 1713453518
transform 1 0 2756 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3564
timestamp 1713453518
transform 1 0 2564 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3565
timestamp 1713453518
transform 1 0 2788 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3566
timestamp 1713453518
transform 1 0 2772 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1713453518
transform 1 0 2772 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1713453518
transform 1 0 2764 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3569
timestamp 1713453518
transform 1 0 2740 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1713453518
transform 1 0 2740 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1713453518
transform 1 0 2740 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_3572
timestamp 1713453518
transform 1 0 2724 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3573
timestamp 1713453518
transform 1 0 2820 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3574
timestamp 1713453518
transform 1 0 2764 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3575
timestamp 1713453518
transform 1 0 2868 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3576
timestamp 1713453518
transform 1 0 2772 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3577
timestamp 1713453518
transform 1 0 2772 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1713453518
transform 1 0 2756 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3579
timestamp 1713453518
transform 1 0 2708 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3580
timestamp 1713453518
transform 1 0 2684 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3581
timestamp 1713453518
transform 1 0 2692 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3582
timestamp 1713453518
transform 1 0 2564 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3583
timestamp 1713453518
transform 1 0 2604 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3584
timestamp 1713453518
transform 1 0 2468 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3585
timestamp 1713453518
transform 1 0 2564 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3586
timestamp 1713453518
transform 1 0 2452 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3587
timestamp 1713453518
transform 1 0 2716 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3588
timestamp 1713453518
transform 1 0 2676 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3589
timestamp 1713453518
transform 1 0 2612 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1713453518
transform 1 0 2604 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3591
timestamp 1713453518
transform 1 0 2580 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3592
timestamp 1713453518
transform 1 0 2660 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3593
timestamp 1713453518
transform 1 0 2620 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1713453518
transform 1 0 2788 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3595
timestamp 1713453518
transform 1 0 2604 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3596
timestamp 1713453518
transform 1 0 2452 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_3597
timestamp 1713453518
transform 1 0 2596 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3598
timestamp 1713453518
transform 1 0 2300 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3599
timestamp 1713453518
transform 1 0 2572 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1713453518
transform 1 0 2420 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1713453518
transform 1 0 2308 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3602
timestamp 1713453518
transform 1 0 2612 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3603
timestamp 1713453518
transform 1 0 2484 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3604
timestamp 1713453518
transform 1 0 2356 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3605
timestamp 1713453518
transform 1 0 2900 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3606
timestamp 1713453518
transform 1 0 2788 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3607
timestamp 1713453518
transform 1 0 2612 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1713453518
transform 1 0 2980 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1713453518
transform 1 0 2820 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1713453518
transform 1 0 2740 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_3611
timestamp 1713453518
transform 1 0 2932 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1713453518
transform 1 0 2876 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1713453518
transform 1 0 2708 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1713453518
transform 1 0 2852 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3615
timestamp 1713453518
transform 1 0 2812 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1713453518
transform 1 0 2924 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3617
timestamp 1713453518
transform 1 0 2868 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1713453518
transform 1 0 2844 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1713453518
transform 1 0 2844 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1713453518
transform 1 0 2772 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1713453518
transform 1 0 2772 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3622
timestamp 1713453518
transform 1 0 2836 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1713453518
transform 1 0 2772 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1713453518
transform 1 0 2012 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3625
timestamp 1713453518
transform 1 0 1916 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1713453518
transform 1 0 1804 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3627
timestamp 1713453518
transform 1 0 1772 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3628
timestamp 1713453518
transform 1 0 2180 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3629
timestamp 1713453518
transform 1 0 1988 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3630
timestamp 1713453518
transform 1 0 2484 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3631
timestamp 1713453518
transform 1 0 2420 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1713453518
transform 1 0 2548 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1713453518
transform 1 0 2468 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1713453518
transform 1 0 2588 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1713453518
transform 1 0 2556 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1713453518
transform 1 0 2676 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3637
timestamp 1713453518
transform 1 0 2636 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3638
timestamp 1713453518
transform 1 0 2684 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3639
timestamp 1713453518
transform 1 0 2652 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3640
timestamp 1713453518
transform 1 0 2572 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1713453518
transform 1 0 2508 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3642
timestamp 1713453518
transform 1 0 2660 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1713453518
transform 1 0 2516 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1713453518
transform 1 0 2900 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1713453518
transform 1 0 2732 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3646
timestamp 1713453518
transform 1 0 2732 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3647
timestamp 1713453518
transform 1 0 2700 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_3648
timestamp 1713453518
transform 1 0 2572 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1713453518
transform 1 0 2572 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3650
timestamp 1713453518
transform 1 0 2516 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1713453518
transform 1 0 2468 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3652
timestamp 1713453518
transform 1 0 2372 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1713453518
transform 1 0 2516 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1713453518
transform 1 0 2428 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1713453518
transform 1 0 2596 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1713453518
transform 1 0 2540 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1713453518
transform 1 0 2452 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3658
timestamp 1713453518
transform 1 0 2412 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3659
timestamp 1713453518
transform 1 0 2452 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3660
timestamp 1713453518
transform 1 0 2452 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1713453518
transform 1 0 2404 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1713453518
transform 1 0 2340 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3663
timestamp 1713453518
transform 1 0 2428 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1713453518
transform 1 0 2380 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3665
timestamp 1713453518
transform 1 0 2284 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1713453518
transform 1 0 2484 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3667
timestamp 1713453518
transform 1 0 2380 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1713453518
transform 1 0 2332 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3669
timestamp 1713453518
transform 1 0 2436 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3670
timestamp 1713453518
transform 1 0 2356 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3671
timestamp 1713453518
transform 1 0 2420 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3672
timestamp 1713453518
transform 1 0 2380 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3673
timestamp 1713453518
transform 1 0 2324 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3674
timestamp 1713453518
transform 1 0 2524 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1713453518
transform 1 0 2324 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1713453518
transform 1 0 2596 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3677
timestamp 1713453518
transform 1 0 2420 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3678
timestamp 1713453518
transform 1 0 2316 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3679
timestamp 1713453518
transform 1 0 1532 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3680
timestamp 1713453518
transform 1 0 932 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3681
timestamp 1713453518
transform 1 0 1532 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3682
timestamp 1713453518
transform 1 0 1508 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1713453518
transform 1 0 1588 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3684
timestamp 1713453518
transform 1 0 1516 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3685
timestamp 1713453518
transform 1 0 3172 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1713453518
transform 1 0 2964 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_3687
timestamp 1713453518
transform 1 0 1828 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1713453518
transform 1 0 1708 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_3689
timestamp 1713453518
transform 1 0 1684 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3690
timestamp 1713453518
transform 1 0 1068 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3691
timestamp 1713453518
transform 1 0 1788 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1713453518
transform 1 0 1516 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1713453518
transform 1 0 1628 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3694
timestamp 1713453518
transform 1 0 1508 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3695
timestamp 1713453518
transform 1 0 2068 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3696
timestamp 1713453518
transform 1 0 2004 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1713453518
transform 1 0 1932 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1713453518
transform 1 0 1932 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3699
timestamp 1713453518
transform 1 0 1844 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3700
timestamp 1713453518
transform 1 0 1820 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3701
timestamp 1713453518
transform 1 0 1820 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3702
timestamp 1713453518
transform 1 0 1620 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_3703
timestamp 1713453518
transform 1 0 1636 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_3704
timestamp 1713453518
transform 1 0 1364 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_3705
timestamp 1713453518
transform 1 0 1308 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3706
timestamp 1713453518
transform 1 0 1244 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1713453518
transform 1 0 1204 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3708
timestamp 1713453518
transform 1 0 1972 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1713453518
transform 1 0 1772 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1713453518
transform 1 0 3196 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3711
timestamp 1713453518
transform 1 0 3148 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3712
timestamp 1713453518
transform 1 0 2916 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_3713
timestamp 1713453518
transform 1 0 2916 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1713453518
transform 1 0 1828 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1713453518
transform 1 0 1828 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3716
timestamp 1713453518
transform 1 0 1788 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3717
timestamp 1713453518
transform 1 0 1268 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3718
timestamp 1713453518
transform 1 0 1228 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3719
timestamp 1713453518
transform 1 0 1268 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3720
timestamp 1713453518
transform 1 0 1220 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3721
timestamp 1713453518
transform 1 0 1172 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3722
timestamp 1713453518
transform 1 0 1500 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3723
timestamp 1713453518
transform 1 0 892 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1713453518
transform 1 0 1572 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1713453518
transform 1 0 1484 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_3726
timestamp 1713453518
transform 1 0 1428 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1713453518
transform 1 0 1204 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3728
timestamp 1713453518
transform 1 0 3228 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_3729
timestamp 1713453518
transform 1 0 3204 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1713453518
transform 1 0 3204 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_3731
timestamp 1713453518
transform 1 0 2996 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1713453518
transform 1 0 2916 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1713453518
transform 1 0 2028 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1713453518
transform 1 0 2028 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3735
timestamp 1713453518
transform 1 0 1580 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3736
timestamp 1713453518
transform 1 0 1596 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3737
timestamp 1713453518
transform 1 0 1180 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1713453518
transform 1 0 1132 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3739
timestamp 1713453518
transform 1 0 1132 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3740
timestamp 1713453518
transform 1 0 1116 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1713453518
transform 1 0 1116 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3742
timestamp 1713453518
transform 1 0 1108 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3743
timestamp 1713453518
transform 1 0 1076 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1713453518
transform 1 0 1076 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3745
timestamp 1713453518
transform 1 0 1052 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3746
timestamp 1713453518
transform 1 0 1844 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1713453518
transform 1 0 1556 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_3748
timestamp 1713453518
transform 1 0 1628 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_3749
timestamp 1713453518
transform 1 0 1556 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_3750
timestamp 1713453518
transform 1 0 1636 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_3751
timestamp 1713453518
transform 1 0 1372 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_3752
timestamp 1713453518
transform 1 0 1356 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3753
timestamp 1713453518
transform 1 0 1316 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1713453518
transform 1 0 1292 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3755
timestamp 1713453518
transform 1 0 1204 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_3756
timestamp 1713453518
transform 1 0 1148 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1713453518
transform 1 0 1476 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_3758
timestamp 1713453518
transform 1 0 908 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_3759
timestamp 1713453518
transform 1 0 1956 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_3760
timestamp 1713453518
transform 1 0 1452 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_3761
timestamp 1713453518
transform 1 0 1380 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_3762
timestamp 1713453518
transform 1 0 1308 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_3763
timestamp 1713453518
transform 1 0 1732 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3764
timestamp 1713453518
transform 1 0 1500 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3765
timestamp 1713453518
transform 1 0 3116 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3766
timestamp 1713453518
transform 1 0 3092 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3767
timestamp 1713453518
transform 1 0 3084 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3768
timestamp 1713453518
transform 1 0 2996 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3769
timestamp 1713453518
transform 1 0 2996 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3770
timestamp 1713453518
transform 1 0 2796 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3771
timestamp 1713453518
transform 1 0 2796 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3772
timestamp 1713453518
transform 1 0 2708 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3773
timestamp 1713453518
transform 1 0 2700 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3774
timestamp 1713453518
transform 1 0 2428 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3775
timestamp 1713453518
transform 1 0 1820 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3776
timestamp 1713453518
transform 1 0 1860 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3777
timestamp 1713453518
transform 1 0 1244 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3778
timestamp 1713453518
transform 1 0 1372 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3779
timestamp 1713453518
transform 1 0 1372 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1713453518
transform 1 0 1340 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3781
timestamp 1713453518
transform 1 0 1276 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3782
timestamp 1713453518
transform 1 0 1236 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3783
timestamp 1713453518
transform 1 0 1228 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1713453518
transform 1 0 1180 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3785
timestamp 1713453518
transform 1 0 1148 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3786
timestamp 1713453518
transform 1 0 1108 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3787
timestamp 1713453518
transform 1 0 1092 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3788
timestamp 1713453518
transform 1 0 1068 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3789
timestamp 1713453518
transform 1 0 1028 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3790
timestamp 1713453518
transform 1 0 2012 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_3791
timestamp 1713453518
transform 1 0 1932 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_3792
timestamp 1713453518
transform 1 0 2092 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_3793
timestamp 1713453518
transform 1 0 1940 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1713453518
transform 1 0 2108 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_3795
timestamp 1713453518
transform 1 0 1444 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_3796
timestamp 1713453518
transform 1 0 2388 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1713453518
transform 1 0 2364 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1713453518
transform 1 0 2060 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3799
timestamp 1713453518
transform 1 0 2060 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1713453518
transform 1 0 2012 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1713453518
transform 1 0 1956 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3802
timestamp 1713453518
transform 1 0 1388 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_3803
timestamp 1713453518
transform 1 0 1356 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3804
timestamp 1713453518
transform 1 0 1300 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3805
timestamp 1713453518
transform 1 0 1244 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_3806
timestamp 1713453518
transform 1 0 1860 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3807
timestamp 1713453518
transform 1 0 1108 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3808
timestamp 1713453518
transform 1 0 2812 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3809
timestamp 1713453518
transform 1 0 1820 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3810
timestamp 1713453518
transform 1 0 1852 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3811
timestamp 1713453518
transform 1 0 1828 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3812
timestamp 1713453518
transform 1 0 2252 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1713453518
transform 1 0 1996 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1713453518
transform 1 0 2012 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1713453518
transform 1 0 1572 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3816
timestamp 1713453518
transform 1 0 1500 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_3817
timestamp 1713453518
transform 1 0 1492 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3818
timestamp 1713453518
transform 1 0 1460 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3819
timestamp 1713453518
transform 1 0 1300 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_3820
timestamp 1713453518
transform 1 0 1284 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3821
timestamp 1713453518
transform 1 0 1220 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1713453518
transform 1 0 1220 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1713453518
transform 1 0 1148 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_3824
timestamp 1713453518
transform 1 0 1404 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1713453518
transform 1 0 1276 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1713453518
transform 1 0 2972 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1713453518
transform 1 0 1468 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1713453518
transform 1 0 1316 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1713453518
transform 1 0 1300 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1713453518
transform 1 0 1268 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3831
timestamp 1713453518
transform 1 0 1252 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1713453518
transform 1 0 1196 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3833
timestamp 1713453518
transform 1 0 1196 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1713453518
transform 1 0 1172 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3835
timestamp 1713453518
transform 1 0 1148 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3836
timestamp 1713453518
transform 1 0 1084 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1713453518
transform 1 0 1076 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1713453518
transform 1 0 1044 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1713453518
transform 1 0 1044 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1713453518
transform 1 0 1036 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3841
timestamp 1713453518
transform 1 0 1036 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3842
timestamp 1713453518
transform 1 0 996 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1713453518
transform 1 0 996 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3844
timestamp 1713453518
transform 1 0 996 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3845
timestamp 1713453518
transform 1 0 2868 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3846
timestamp 1713453518
transform 1 0 2852 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1713453518
transform 1 0 2548 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1713453518
transform 1 0 1116 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_3849
timestamp 1713453518
transform 1 0 3140 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1713453518
transform 1 0 2516 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1713453518
transform 1 0 2428 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3852
timestamp 1713453518
transform 1 0 2100 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3853
timestamp 1713453518
transform 1 0 2628 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3854
timestamp 1713453518
transform 1 0 2524 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3855
timestamp 1713453518
transform 1 0 2972 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1713453518
transform 1 0 2540 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3857
timestamp 1713453518
transform 1 0 2284 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3858
timestamp 1713453518
transform 1 0 1716 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3859
timestamp 1713453518
transform 1 0 1436 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3860
timestamp 1713453518
transform 1 0 1124 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3861
timestamp 1713453518
transform 1 0 1084 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3862
timestamp 1713453518
transform 1 0 1084 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3863
timestamp 1713453518
transform 1 0 1068 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3864
timestamp 1713453518
transform 1 0 1060 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3865
timestamp 1713453518
transform 1 0 1060 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3866
timestamp 1713453518
transform 1 0 1060 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3867
timestamp 1713453518
transform 1 0 1028 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3868
timestamp 1713453518
transform 1 0 1028 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3869
timestamp 1713453518
transform 1 0 1020 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3870
timestamp 1713453518
transform 1 0 3244 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3871
timestamp 1713453518
transform 1 0 3132 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3872
timestamp 1713453518
transform 1 0 2204 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3873
timestamp 1713453518
transform 1 0 2140 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3874
timestamp 1713453518
transform 1 0 2076 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3875
timestamp 1713453518
transform 1 0 2076 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3876
timestamp 1713453518
transform 1 0 1404 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3877
timestamp 1713453518
transform 1 0 3172 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3878
timestamp 1713453518
transform 1 0 1348 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3879
timestamp 1713453518
transform 1 0 1420 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3880
timestamp 1713453518
transform 1 0 1420 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3881
timestamp 1713453518
transform 1 0 1316 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3882
timestamp 1713453518
transform 1 0 1316 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_3883
timestamp 1713453518
transform 1 0 1284 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_3884
timestamp 1713453518
transform 1 0 1276 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1713453518
transform 1 0 1532 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3886
timestamp 1713453518
transform 1 0 1508 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3887
timestamp 1713453518
transform 1 0 1492 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1713453518
transform 1 0 1428 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1713453518
transform 1 0 1428 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1713453518
transform 1 0 1332 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3891
timestamp 1713453518
transform 1 0 1300 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3892
timestamp 1713453518
transform 1 0 1300 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3893
timestamp 1713453518
transform 1 0 1268 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3894
timestamp 1713453518
transform 1 0 1244 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3895
timestamp 1713453518
transform 1 0 1236 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3896
timestamp 1713453518
transform 1 0 1212 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3897
timestamp 1713453518
transform 1 0 1204 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3898
timestamp 1713453518
transform 1 0 1196 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1713453518
transform 1 0 1188 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3900
timestamp 1713453518
transform 1 0 1188 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3901
timestamp 1713453518
transform 1 0 1164 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1713453518
transform 1 0 996 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3903
timestamp 1713453518
transform 1 0 996 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3904
timestamp 1713453518
transform 1 0 948 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3905
timestamp 1713453518
transform 1 0 948 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3906
timestamp 1713453518
transform 1 0 940 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3907
timestamp 1713453518
transform 1 0 940 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3908
timestamp 1713453518
transform 1 0 924 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1713453518
transform 1 0 924 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3910
timestamp 1713453518
transform 1 0 876 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3911
timestamp 1713453518
transform 1 0 860 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3912
timestamp 1713453518
transform 1 0 2556 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_3913
timestamp 1713453518
transform 1 0 1140 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_3914
timestamp 1713453518
transform 1 0 3332 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_3915
timestamp 1713453518
transform 1 0 2540 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_3916
timestamp 1713453518
transform 1 0 2572 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3917
timestamp 1713453518
transform 1 0 2388 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1713453518
transform 1 0 2748 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1713453518
transform 1 0 2660 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_3920
timestamp 1713453518
transform 1 0 3196 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_3921
timestamp 1713453518
transform 1 0 3124 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_3922
timestamp 1713453518
transform 1 0 2940 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_3923
timestamp 1713453518
transform 1 0 2916 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1713453518
transform 1 0 2796 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_3925
timestamp 1713453518
transform 1 0 2636 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_3926
timestamp 1713453518
transform 1 0 2596 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1713453518
transform 1 0 2532 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1713453518
transform 1 0 2524 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1713453518
transform 1 0 2476 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3930
timestamp 1713453518
transform 1 0 2420 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3931
timestamp 1713453518
transform 1 0 1860 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1713453518
transform 1 0 1860 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1713453518
transform 1 0 1756 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3934
timestamp 1713453518
transform 1 0 1756 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3935
timestamp 1713453518
transform 1 0 1188 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3936
timestamp 1713453518
transform 1 0 2948 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_3937
timestamp 1713453518
transform 1 0 2820 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1713453518
transform 1 0 2820 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1713453518
transform 1 0 2676 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1713453518
transform 1 0 3364 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_3941
timestamp 1713453518
transform 1 0 3196 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1713453518
transform 1 0 2940 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1713453518
transform 1 0 2940 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1713453518
transform 1 0 2764 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1713453518
transform 1 0 3372 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1713453518
transform 1 0 3012 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1713453518
transform 1 0 2420 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_3948
timestamp 1713453518
transform 1 0 1148 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3949
timestamp 1713453518
transform 1 0 1044 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1713453518
transform 1 0 1124 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1713453518
transform 1 0 1020 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1713453518
transform 1 0 1020 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3953
timestamp 1713453518
transform 1 0 988 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1713453518
transform 1 0 972 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3955
timestamp 1713453518
transform 1 0 3220 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_3956
timestamp 1713453518
transform 1 0 3068 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_3957
timestamp 1713453518
transform 1 0 2644 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1713453518
transform 1 0 2556 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_3959
timestamp 1713453518
transform 1 0 2556 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3960
timestamp 1713453518
transform 1 0 2476 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1713453518
transform 1 0 2388 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3962
timestamp 1713453518
transform 1 0 2364 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1713453518
transform 1 0 1396 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1713453518
transform 1 0 2748 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3965
timestamp 1713453518
transform 1 0 2732 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3966
timestamp 1713453518
transform 1 0 2692 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3967
timestamp 1713453518
transform 1 0 2588 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3968
timestamp 1713453518
transform 1 0 2580 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3969
timestamp 1713453518
transform 1 0 1276 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3970
timestamp 1713453518
transform 1 0 3220 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3971
timestamp 1713453518
transform 1 0 3212 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_3972
timestamp 1713453518
transform 1 0 3196 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3973
timestamp 1713453518
transform 1 0 3196 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_3974
timestamp 1713453518
transform 1 0 3124 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3975
timestamp 1713453518
transform 1 0 3084 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3976
timestamp 1713453518
transform 1 0 3076 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3977
timestamp 1713453518
transform 1 0 2508 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3978
timestamp 1713453518
transform 1 0 1452 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3979
timestamp 1713453518
transform 1 0 1452 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3980
timestamp 1713453518
transform 1 0 1124 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3981
timestamp 1713453518
transform 1 0 3116 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_3982
timestamp 1713453518
transform 1 0 2492 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_3983
timestamp 1713453518
transform 1 0 2524 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3984
timestamp 1713453518
transform 1 0 2316 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3985
timestamp 1713453518
transform 1 0 2724 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_3986
timestamp 1713453518
transform 1 0 2628 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_3987
timestamp 1713453518
transform 1 0 2876 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3988
timestamp 1713453518
transform 1 0 2844 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_3989
timestamp 1713453518
transform 1 0 3388 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3990
timestamp 1713453518
transform 1 0 3364 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3991
timestamp 1713453518
transform 1 0 3052 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1713453518
transform 1 0 2924 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_3993
timestamp 1713453518
transform 1 0 3356 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1713453518
transform 1 0 3308 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_3995
timestamp 1713453518
transform 1 0 2540 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_3996
timestamp 1713453518
transform 1 0 2436 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_3997
timestamp 1713453518
transform 1 0 2260 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_3998
timestamp 1713453518
transform 1 0 1276 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3999
timestamp 1713453518
transform 1 0 1140 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_4000
timestamp 1713453518
transform 1 0 1140 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4001
timestamp 1713453518
transform 1 0 1108 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4002
timestamp 1713453518
transform 1 0 1092 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4003
timestamp 1713453518
transform 1 0 1092 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4004
timestamp 1713453518
transform 1 0 1076 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4005
timestamp 1713453518
transform 1 0 1076 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4006
timestamp 1713453518
transform 1 0 1068 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4007
timestamp 1713453518
transform 1 0 1068 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4008
timestamp 1713453518
transform 1 0 1020 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4009
timestamp 1713453518
transform 1 0 1020 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4010
timestamp 1713453518
transform 1 0 1020 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4011
timestamp 1713453518
transform 1 0 1020 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4012
timestamp 1713453518
transform 1 0 988 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4013
timestamp 1713453518
transform 1 0 988 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4014
timestamp 1713453518
transform 1 0 956 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1713453518
transform 1 0 956 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4016
timestamp 1713453518
transform 1 0 948 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4017
timestamp 1713453518
transform 1 0 3388 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_4018
timestamp 1713453518
transform 1 0 3124 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1713453518
transform 1 0 2780 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4020
timestamp 1713453518
transform 1 0 2748 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4021
timestamp 1713453518
transform 1 0 2708 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4022
timestamp 1713453518
transform 1 0 2492 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4023
timestamp 1713453518
transform 1 0 2492 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4024
timestamp 1713453518
transform 1 0 2460 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1713453518
transform 1 0 2452 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4026
timestamp 1713453518
transform 1 0 2444 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4027
timestamp 1713453518
transform 1 0 1308 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4028
timestamp 1713453518
transform 1 0 2804 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4029
timestamp 1713453518
transform 1 0 2804 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4030
timestamp 1713453518
transform 1 0 2788 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4031
timestamp 1713453518
transform 1 0 2764 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4032
timestamp 1713453518
transform 1 0 2756 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4033
timestamp 1713453518
transform 1 0 2708 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4034
timestamp 1713453518
transform 1 0 2708 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4035
timestamp 1713453518
transform 1 0 2516 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4036
timestamp 1713453518
transform 1 0 2516 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4037
timestamp 1713453518
transform 1 0 2460 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4038
timestamp 1713453518
transform 1 0 2452 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1713453518
transform 1 0 1260 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4040
timestamp 1713453518
transform 1 0 2564 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1713453518
transform 1 0 1076 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_4042
timestamp 1713453518
transform 1 0 3236 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_4043
timestamp 1713453518
transform 1 0 2540 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_4044
timestamp 1713453518
transform 1 0 2452 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_4045
timestamp 1713453518
transform 1 0 2140 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_4046
timestamp 1713453518
transform 1 0 2620 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_4047
timestamp 1713453518
transform 1 0 2532 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_4048
timestamp 1713453518
transform 1 0 3100 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4049
timestamp 1713453518
transform 1 0 3092 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_4050
timestamp 1713453518
transform 1 0 3020 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_4051
timestamp 1713453518
transform 1 0 2924 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_4052
timestamp 1713453518
transform 1 0 2796 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4053
timestamp 1713453518
transform 1 0 2796 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4054
timestamp 1713453518
transform 1 0 2660 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_4055
timestamp 1713453518
transform 1 0 2596 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_4056
timestamp 1713453518
transform 1 0 2596 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4057
timestamp 1713453518
transform 1 0 2348 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_4058
timestamp 1713453518
transform 1 0 3340 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_4059
timestamp 1713453518
transform 1 0 3300 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_4060
timestamp 1713453518
transform 1 0 3052 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_4061
timestamp 1713453518
transform 1 0 2668 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_4062
timestamp 1713453518
transform 1 0 1524 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_4063
timestamp 1713453518
transform 1 0 2276 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_4064
timestamp 1713453518
transform 1 0 1516 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_4065
timestamp 1713453518
transform 1 0 3300 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_4066
timestamp 1713453518
transform 1 0 3244 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_4067
timestamp 1713453518
transform 1 0 2356 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_4068
timestamp 1713453518
transform 1 0 3324 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_4069
timestamp 1713453518
transform 1 0 3204 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_4070
timestamp 1713453518
transform 1 0 3236 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_4071
timestamp 1713453518
transform 1 0 3212 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_4072
timestamp 1713453518
transform 1 0 1548 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_4073
timestamp 1713453518
transform 1 0 1436 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_4074
timestamp 1713453518
transform 1 0 1476 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1713453518
transform 1 0 1308 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4076
timestamp 1713453518
transform 1 0 1324 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4077
timestamp 1713453518
transform 1 0 1292 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4078
timestamp 1713453518
transform 1 0 1908 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_4079
timestamp 1713453518
transform 1 0 1092 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_4080
timestamp 1713453518
transform 1 0 3268 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_4081
timestamp 1713453518
transform 1 0 2516 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_4082
timestamp 1713453518
transform 1 0 2484 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_4083
timestamp 1713453518
transform 1 0 2300 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_4084
timestamp 1713453518
transform 1 0 2292 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4085
timestamp 1713453518
transform 1 0 1876 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4086
timestamp 1713453518
transform 1 0 2028 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_4087
timestamp 1713453518
transform 1 0 1884 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1713453518
transform 1 0 2076 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_4089
timestamp 1713453518
transform 1 0 1996 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_4090
timestamp 1713453518
transform 1 0 2460 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_4091
timestamp 1713453518
transform 1 0 2124 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_4092
timestamp 1713453518
transform 1 0 3332 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_4093
timestamp 1713453518
transform 1 0 3308 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_4094
timestamp 1713453518
transform 1 0 3124 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1713453518
transform 1 0 2444 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_4096
timestamp 1713453518
transform 1 0 1628 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_4097
timestamp 1713453518
transform 1 0 1540 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4098
timestamp 1713453518
transform 1 0 1492 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1713453518
transform 1 0 1556 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4100
timestamp 1713453518
transform 1 0 1124 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1713453518
transform 1 0 1516 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4102
timestamp 1713453518
transform 1 0 1444 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4103
timestamp 1713453518
transform 1 0 1372 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1713453518
transform 1 0 3364 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_4105
timestamp 1713453518
transform 1 0 3236 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_4106
timestamp 1713453518
transform 1 0 3212 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_4107
timestamp 1713453518
transform 1 0 3092 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_4108
timestamp 1713453518
transform 1 0 1644 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_4109
timestamp 1713453518
transform 1 0 1364 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_4110
timestamp 1713453518
transform 1 0 1604 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4111
timestamp 1713453518
transform 1 0 1388 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1713453518
transform 1 0 1564 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4113
timestamp 1713453518
transform 1 0 1348 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4114
timestamp 1713453518
transform 1 0 1324 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1713453518
transform 1 0 1188 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4116
timestamp 1713453518
transform 1 0 1852 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_4117
timestamp 1713453518
transform 1 0 1052 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_4118
timestamp 1713453518
transform 1 0 3268 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_4119
timestamp 1713453518
transform 1 0 1812 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1713453518
transform 1 0 1924 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4121
timestamp 1713453518
transform 1 0 1836 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4122
timestamp 1713453518
transform 1 0 2460 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4123
timestamp 1713453518
transform 1 0 1892 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4124
timestamp 1713453518
transform 1 0 3268 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4125
timestamp 1713453518
transform 1 0 3132 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_4126
timestamp 1713453518
transform 1 0 3132 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4127
timestamp 1713453518
transform 1 0 3132 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4128
timestamp 1713453518
transform 1 0 2884 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4129
timestamp 1713453518
transform 1 0 2796 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_4130
timestamp 1713453518
transform 1 0 2796 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4131
timestamp 1713453518
transform 1 0 2556 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4132
timestamp 1713453518
transform 1 0 2508 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4133
timestamp 1713453518
transform 1 0 1692 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_4134
timestamp 1713453518
transform 1 0 2628 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4135
timestamp 1713453518
transform 1 0 2532 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4136
timestamp 1713453518
transform 1 0 1540 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_4137
timestamp 1713453518
transform 1 0 3412 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4138
timestamp 1713453518
transform 1 0 3348 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4139
timestamp 1713453518
transform 1 0 3156 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_4140
timestamp 1713453518
transform 1 0 3156 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4141
timestamp 1713453518
transform 1 0 2540 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_4142
timestamp 1713453518
transform 1 0 1468 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1713453518
transform 1 0 1636 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1713453518
transform 1 0 1116 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4145
timestamp 1713453518
transform 1 0 1508 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1713453518
transform 1 0 1228 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4147
timestamp 1713453518
transform 1 0 1228 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4148
timestamp 1713453518
transform 1 0 1180 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4149
timestamp 1713453518
transform 1 0 3412 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_4150
timestamp 1713453518
transform 1 0 3260 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_4151
timestamp 1713453518
transform 1 0 3236 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_4152
timestamp 1713453518
transform 1 0 3148 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1713453518
transform 1 0 3084 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_4154
timestamp 1713453518
transform 1 0 2796 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_4155
timestamp 1713453518
transform 1 0 1548 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4156
timestamp 1713453518
transform 1 0 1420 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_4157
timestamp 1713453518
transform 1 0 1428 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1713453518
transform 1 0 1340 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4159
timestamp 1713453518
transform 1 0 1588 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4160
timestamp 1713453518
transform 1 0 1548 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4161
timestamp 1713453518
transform 1 0 1484 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4162
timestamp 1713453518
transform 1 0 1196 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4163
timestamp 1713453518
transform 1 0 1276 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4164
timestamp 1713453518
transform 1 0 1188 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4165
timestamp 1713453518
transform 1 0 2020 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4166
timestamp 1713453518
transform 1 0 1044 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1713453518
transform 1 0 2892 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_4168
timestamp 1713453518
transform 1 0 1988 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_4169
timestamp 1713453518
transform 1 0 2356 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4170
timestamp 1713453518
transform 1 0 2292 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4171
timestamp 1713453518
transform 1 0 2292 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4172
timestamp 1713453518
transform 1 0 2100 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_4173
timestamp 1713453518
transform 1 0 3036 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4174
timestamp 1713453518
transform 1 0 2892 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4175
timestamp 1713453518
transform 1 0 2692 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4176
timestamp 1713453518
transform 1 0 2444 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4177
timestamp 1713453518
transform 1 0 1748 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4178
timestamp 1713453518
transform 1 0 1788 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4179
timestamp 1713453518
transform 1 0 1548 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4180
timestamp 1713453518
transform 1 0 1724 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4181
timestamp 1713453518
transform 1 0 1156 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4182
timestamp 1713453518
transform 1 0 1508 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4183
timestamp 1713453518
transform 1 0 1492 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1713453518
transform 1 0 1492 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4185
timestamp 1713453518
transform 1 0 1348 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4186
timestamp 1713453518
transform 1 0 1244 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4187
timestamp 1713453518
transform 1 0 2988 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4188
timestamp 1713453518
transform 1 0 2860 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1713453518
transform 1 0 2852 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4190
timestamp 1713453518
transform 1 0 2788 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4191
timestamp 1713453518
transform 1 0 2756 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4192
timestamp 1713453518
transform 1 0 2644 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_4193
timestamp 1713453518
transform 1 0 1828 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4194
timestamp 1713453518
transform 1 0 1636 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4195
timestamp 1713453518
transform 1 0 1724 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1713453518
transform 1 0 1628 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4197
timestamp 1713453518
transform 1 0 1540 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4198
timestamp 1713453518
transform 1 0 1492 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4199
timestamp 1713453518
transform 1 0 1460 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4200
timestamp 1713453518
transform 1 0 1292 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1713453518
transform 1 0 1524 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1713453518
transform 1 0 1460 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4203
timestamp 1713453518
transform 1 0 2196 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4204
timestamp 1713453518
transform 1 0 1116 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4205
timestamp 1713453518
transform 1 0 1116 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4206
timestamp 1713453518
transform 1 0 1092 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4207
timestamp 1713453518
transform 1 0 2828 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4208
timestamp 1713453518
transform 1 0 2172 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4209
timestamp 1713453518
transform 1 0 2316 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1713453518
transform 1 0 2100 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1713453518
transform 1 0 2932 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4212
timestamp 1713453518
transform 1 0 2892 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4213
timestamp 1713453518
transform 1 0 2828 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1713453518
transform 1 0 2348 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1713453518
transform 1 0 1740 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4216
timestamp 1713453518
transform 1 0 1868 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4217
timestamp 1713453518
transform 1 0 1772 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4218
timestamp 1713453518
transform 1 0 1644 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4219
timestamp 1713453518
transform 1 0 1604 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4220
timestamp 1713453518
transform 1 0 1652 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4221
timestamp 1713453518
transform 1 0 1140 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4222
timestamp 1713453518
transform 1 0 1572 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4223
timestamp 1713453518
transform 1 0 1396 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4224
timestamp 1713453518
transform 1 0 1372 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1713453518
transform 1 0 3012 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4226
timestamp 1713453518
transform 1 0 2796 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4227
timestamp 1713453518
transform 1 0 2788 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4228
timestamp 1713453518
transform 1 0 2756 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4229
timestamp 1713453518
transform 1 0 1756 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4230
timestamp 1713453518
transform 1 0 1628 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4231
timestamp 1713453518
transform 1 0 1716 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1713453518
transform 1 0 1340 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4233
timestamp 1713453518
transform 1 0 1356 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4234
timestamp 1713453518
transform 1 0 1268 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4235
timestamp 1713453518
transform 1 0 1236 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4236
timestamp 1713453518
transform 1 0 1756 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4237
timestamp 1713453518
transform 1 0 1716 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1713453518
transform 1 0 1596 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4239
timestamp 1713453518
transform 1 0 1508 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1713453518
transform 1 0 1212 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4241
timestamp 1713453518
transform 1 0 1172 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4242
timestamp 1713453518
transform 1 0 2100 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4243
timestamp 1713453518
transform 1 0 1068 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4244
timestamp 1713453518
transform 1 0 3028 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4245
timestamp 1713453518
transform 1 0 2060 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4246
timestamp 1713453518
transform 1 0 2316 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4247
timestamp 1713453518
transform 1 0 2156 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4248
timestamp 1713453518
transform 1 0 2540 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4249
timestamp 1713453518
transform 1 0 2460 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4250
timestamp 1713453518
transform 1 0 2276 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4251
timestamp 1713453518
transform 1 0 3316 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4252
timestamp 1713453518
transform 1 0 3076 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4253
timestamp 1713453518
transform 1 0 3076 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1713453518
transform 1 0 2908 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4255
timestamp 1713453518
transform 1 0 2908 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4256
timestamp 1713453518
transform 1 0 2564 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4257
timestamp 1713453518
transform 1 0 1476 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4258
timestamp 1713453518
transform 1 0 2012 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4259
timestamp 1713453518
transform 1 0 1716 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1713453518
transform 1 0 1652 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4261
timestamp 1713453518
transform 1 0 1116 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4262
timestamp 1713453518
transform 1 0 3148 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4263
timestamp 1713453518
transform 1 0 3004 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4264
timestamp 1713453518
transform 1 0 1428 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4265
timestamp 1713453518
transform 1 0 1396 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4266
timestamp 1713453518
transform 1 0 1804 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4267
timestamp 1713453518
transform 1 0 1012 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4268
timestamp 1713453518
transform 1 0 3300 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4269
timestamp 1713453518
transform 1 0 1788 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4270
timestamp 1713453518
transform 1 0 1940 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4271
timestamp 1713453518
transform 1 0 1868 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4272
timestamp 1713453518
transform 1 0 2460 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4273
timestamp 1713453518
transform 1 0 1868 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4274
timestamp 1713453518
transform 1 0 3340 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4275
timestamp 1713453518
transform 1 0 3316 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1713453518
transform 1 0 3092 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4277
timestamp 1713453518
transform 1 0 2796 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4278
timestamp 1713453518
transform 1 0 2772 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1713453518
transform 1 0 2036 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4280
timestamp 1713453518
transform 1 0 1772 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4281
timestamp 1713453518
transform 1 0 1668 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4282
timestamp 1713453518
transform 1 0 1564 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4283
timestamp 1713453518
transform 1 0 1724 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4284
timestamp 1713453518
transform 1 0 1076 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4285
timestamp 1713453518
transform 1 0 3412 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4286
timestamp 1713453518
transform 1 0 3292 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4287
timestamp 1713453518
transform 1 0 3316 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4288
timestamp 1713453518
transform 1 0 3260 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4289
timestamp 1713453518
transform 1 0 3228 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4290
timestamp 1713453518
transform 1 0 3116 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4291
timestamp 1713453518
transform 1 0 3332 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4292
timestamp 1713453518
transform 1 0 3300 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4293
timestamp 1713453518
transform 1 0 3268 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4294
timestamp 1713453518
transform 1 0 3252 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4295
timestamp 1713453518
transform 1 0 3140 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4296
timestamp 1713453518
transform 1 0 3108 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4297
timestamp 1713453518
transform 1 0 3108 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1713453518
transform 1 0 3100 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4299
timestamp 1713453518
transform 1 0 2508 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4300
timestamp 1713453518
transform 1 0 1028 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1713453518
transform 1 0 3284 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4302
timestamp 1713453518
transform 1 0 2468 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4303
timestamp 1713453518
transform 1 0 2404 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4304
timestamp 1713453518
transform 1 0 2372 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4305
timestamp 1713453518
transform 1 0 2572 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1713453518
transform 1 0 2468 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4307
timestamp 1713453518
transform 1 0 3116 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4308
timestamp 1713453518
transform 1 0 3108 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4309
timestamp 1713453518
transform 1 0 2996 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4310
timestamp 1713453518
transform 1 0 2940 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4311
timestamp 1713453518
transform 1 0 2876 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4312
timestamp 1713453518
transform 1 0 2716 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4313
timestamp 1713453518
transform 1 0 2708 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4314
timestamp 1713453518
transform 1 0 2676 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4315
timestamp 1713453518
transform 1 0 2444 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4316
timestamp 1713453518
transform 1 0 1836 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4317
timestamp 1713453518
transform 1 0 2908 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4318
timestamp 1713453518
transform 1 0 2764 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4319
timestamp 1713453518
transform 1 0 3348 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4320
timestamp 1713453518
transform 1 0 3324 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4321
timestamp 1713453518
transform 1 0 3132 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4322
timestamp 1713453518
transform 1 0 2892 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1713453518
transform 1 0 2356 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4324
timestamp 1713453518
transform 1 0 1836 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4325
timestamp 1713453518
transform 1 0 1724 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4326
timestamp 1713453518
transform 1 0 1604 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4327
timestamp 1713453518
transform 1 0 1732 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4328
timestamp 1713453518
transform 1 0 1124 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4329
timestamp 1713453518
transform 1 0 3412 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1713453518
transform 1 0 3244 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4331
timestamp 1713453518
transform 1 0 3260 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4332
timestamp 1713453518
transform 1 0 3244 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1713453518
transform 1 0 3228 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4334
timestamp 1713453518
transform 1 0 3180 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4335
timestamp 1713453518
transform 1 0 1772 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4336
timestamp 1713453518
transform 1 0 1700 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4337
timestamp 1713453518
transform 1 0 1612 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4338
timestamp 1713453518
transform 1 0 1612 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4339
timestamp 1713453518
transform 1 0 1532 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4340
timestamp 1713453518
transform 1 0 1188 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4341
timestamp 1713453518
transform 1 0 2404 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1713453518
transform 1 0 1068 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4343
timestamp 1713453518
transform 1 0 3228 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1713453518
transform 1 0 2348 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4345
timestamp 1713453518
transform 1 0 2428 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4346
timestamp 1713453518
transform 1 0 2148 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4347
timestamp 1713453518
transform 1 0 2876 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4348
timestamp 1713453518
transform 1 0 2604 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4349
timestamp 1713453518
transform 1 0 1900 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4350
timestamp 1713453518
transform 1 0 3316 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4351
timestamp 1713453518
transform 1 0 3284 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4352
timestamp 1713453518
transform 1 0 2908 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4353
timestamp 1713453518
transform 1 0 2908 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4354
timestamp 1713453518
transform 1 0 2764 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4355
timestamp 1713453518
transform 1 0 2764 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4356
timestamp 1713453518
transform 1 0 2644 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4357
timestamp 1713453518
transform 1 0 1412 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4358
timestamp 1713453518
transform 1 0 2388 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4359
timestamp 1713453518
transform 1 0 1820 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4360
timestamp 1713453518
transform 1 0 3412 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4361
timestamp 1713453518
transform 1 0 3196 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4362
timestamp 1713453518
transform 1 0 3228 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4363
timestamp 1713453518
transform 1 0 3204 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4364
timestamp 1713453518
transform 1 0 1852 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4365
timestamp 1713453518
transform 1 0 1684 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4366
timestamp 1713453518
transform 1 0 1324 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4367
timestamp 1713453518
transform 1 0 1268 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4368
timestamp 1713453518
transform 1 0 2356 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4369
timestamp 1713453518
transform 1 0 1092 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4370
timestamp 1713453518
transform 1 0 2980 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4371
timestamp 1713453518
transform 1 0 2316 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1713453518
transform 1 0 2244 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4373
timestamp 1713453518
transform 1 0 2052 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4374
timestamp 1713453518
transform 1 0 2516 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4375
timestamp 1713453518
transform 1 0 2316 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4376
timestamp 1713453518
transform 1 0 3340 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4377
timestamp 1713453518
transform 1 0 3300 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4378
timestamp 1713453518
transform 1 0 2796 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4379
timestamp 1713453518
transform 1 0 2548 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4380
timestamp 1713453518
transform 1 0 1700 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4381
timestamp 1713453518
transform 1 0 1796 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4382
timestamp 1713453518
transform 1 0 1764 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4383
timestamp 1713453518
transform 1 0 1852 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4384
timestamp 1713453518
transform 1 0 1164 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4385
timestamp 1713453518
transform 1 0 1788 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4386
timestamp 1713453518
transform 1 0 1652 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4387
timestamp 1713453518
transform 1 0 1588 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4388
timestamp 1713453518
transform 1 0 1484 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1713453518
transform 1 0 1468 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4390
timestamp 1713453518
transform 1 0 1444 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4391
timestamp 1713453518
transform 1 0 3340 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4392
timestamp 1713453518
transform 1 0 3012 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4393
timestamp 1713453518
transform 1 0 3092 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4394
timestamp 1713453518
transform 1 0 3060 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4395
timestamp 1713453518
transform 1 0 3092 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4396
timestamp 1713453518
transform 1 0 2940 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4397
timestamp 1713453518
transform 1 0 1772 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4398
timestamp 1713453518
transform 1 0 1612 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4399
timestamp 1713453518
transform 1 0 1644 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4400
timestamp 1713453518
transform 1 0 1580 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1713453518
transform 1 0 1708 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4402
timestamp 1713453518
transform 1 0 1612 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4403
timestamp 1713453518
transform 1 0 1476 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4404
timestamp 1713453518
transform 1 0 1476 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4405
timestamp 1713453518
transform 1 0 1460 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4406
timestamp 1713453518
transform 1 0 1444 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4407
timestamp 1713453518
transform 1 0 1444 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4408
timestamp 1713453518
transform 1 0 1548 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1713453518
transform 1 0 1476 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4410
timestamp 1713453518
transform 1 0 2340 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4411
timestamp 1713453518
transform 1 0 1092 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4412
timestamp 1713453518
transform 1 0 3284 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4413
timestamp 1713453518
transform 1 0 2348 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4414
timestamp 1713453518
transform 1 0 2260 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4415
timestamp 1713453518
transform 1 0 2156 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4416
timestamp 1713453518
transform 1 0 2500 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1713453518
transform 1 0 2324 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4418
timestamp 1713453518
transform 1 0 2716 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1713453518
transform 1 0 2604 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4420
timestamp 1713453518
transform 1 0 1764 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4421
timestamp 1713453518
transform 1 0 3316 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1713453518
transform 1 0 3316 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4423
timestamp 1713453518
transform 1 0 3284 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4424
timestamp 1713453518
transform 1 0 3132 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4425
timestamp 1713453518
transform 1 0 2588 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4426
timestamp 1713453518
transform 1 0 1804 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1713453518
transform 1 0 1836 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4428
timestamp 1713453518
transform 1 0 1196 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4429
timestamp 1713453518
transform 1 0 3356 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4430
timestamp 1713453518
transform 1 0 3300 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1713453518
transform 1 0 3316 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4432
timestamp 1713453518
transform 1 0 3244 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4433
timestamp 1713453518
transform 1 0 1724 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4434
timestamp 1713453518
transform 1 0 1580 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4435
timestamp 1713453518
transform 1 0 1764 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4436
timestamp 1713453518
transform 1 0 1700 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4437
timestamp 1713453518
transform 1 0 1676 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4438
timestamp 1713453518
transform 1 0 1588 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4439
timestamp 1713453518
transform 1 0 1412 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4440
timestamp 1713453518
transform 1 0 1556 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4441
timestamp 1713453518
transform 1 0 1508 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4442
timestamp 1713453518
transform 1 0 2340 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4443
timestamp 1713453518
transform 1 0 1092 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_4444
timestamp 1713453518
transform 1 0 1076 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4445
timestamp 1713453518
transform 1 0 1060 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1713453518
transform 1 0 3068 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1713453518
transform 1 0 2316 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4448
timestamp 1713453518
transform 1 0 2252 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4449
timestamp 1713453518
transform 1 0 2124 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4450
timestamp 1713453518
transform 1 0 2428 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4451
timestamp 1713453518
transform 1 0 2308 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4452
timestamp 1713453518
transform 1 0 2596 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4453
timestamp 1713453518
transform 1 0 2412 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4454
timestamp 1713453518
transform 1 0 2324 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4455
timestamp 1713453518
transform 1 0 2324 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4456
timestamp 1713453518
transform 1 0 1740 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4457
timestamp 1713453518
transform 1 0 3268 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4458
timestamp 1713453518
transform 1 0 3204 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4459
timestamp 1713453518
transform 1 0 3204 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1713453518
transform 1 0 2988 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4461
timestamp 1713453518
transform 1 0 2468 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4462
timestamp 1713453518
transform 1 0 1780 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_4463
timestamp 1713453518
transform 1 0 2196 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4464
timestamp 1713453518
transform 1 0 1868 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1713453518
transform 1 0 1756 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1713453518
transform 1 0 1692 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4467
timestamp 1713453518
transform 1 0 1820 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4468
timestamp 1713453518
transform 1 0 1124 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4469
timestamp 1713453518
transform 1 0 1628 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4470
timestamp 1713453518
transform 1 0 1532 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4471
timestamp 1713453518
transform 1 0 1332 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4472
timestamp 1713453518
transform 1 0 1252 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1713453518
transform 1 0 1180 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4474
timestamp 1713453518
transform 1 0 3260 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4475
timestamp 1713453518
transform 1 0 3044 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4476
timestamp 1713453518
transform 1 0 3020 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4477
timestamp 1713453518
transform 1 0 2900 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4478
timestamp 1713453518
transform 1 0 1700 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4479
timestamp 1713453518
transform 1 0 1596 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4480
timestamp 1713453518
transform 1 0 1764 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4481
timestamp 1713453518
transform 1 0 1572 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1713453518
transform 1 0 1612 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4483
timestamp 1713453518
transform 1 0 1508 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4484
timestamp 1713453518
transform 1 0 1316 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4485
timestamp 1713453518
transform 1 0 1492 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1713453518
transform 1 0 1420 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4487
timestamp 1713453518
transform 1 0 1908 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4488
timestamp 1713453518
transform 1 0 1044 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4489
timestamp 1713453518
transform 1 0 2636 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4490
timestamp 1713453518
transform 1 0 1892 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4491
timestamp 1713453518
transform 1 0 2012 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4492
timestamp 1713453518
transform 1 0 1932 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4493
timestamp 1713453518
transform 1 0 2380 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4494
timestamp 1713453518
transform 1 0 1972 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4495
timestamp 1713453518
transform 1 0 2596 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4496
timestamp 1713453518
transform 1 0 2324 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4497
timestamp 1713453518
transform 1 0 1764 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4498
timestamp 1713453518
transform 1 0 2980 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1713453518
transform 1 0 2852 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4500
timestamp 1713453518
transform 1 0 2756 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1713453518
transform 1 0 2452 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4502
timestamp 1713453518
transform 1 0 2404 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4503
timestamp 1713453518
transform 1 0 1660 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4504
timestamp 1713453518
transform 1 0 2028 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4505
timestamp 1713453518
transform 1 0 1868 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4506
timestamp 1713453518
transform 1 0 1772 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4507
timestamp 1713453518
transform 1 0 1684 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4508
timestamp 1713453518
transform 1 0 1796 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1713453518
transform 1 0 1100 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4510
timestamp 1713453518
transform 1 0 1668 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4511
timestamp 1713453518
transform 1 0 1316 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4512
timestamp 1713453518
transform 1 0 2964 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4513
timestamp 1713453518
transform 1 0 2676 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4514
timestamp 1713453518
transform 1 0 2756 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4515
timestamp 1713453518
transform 1 0 2708 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4516
timestamp 1713453518
transform 1 0 1700 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4517
timestamp 1713453518
transform 1 0 1564 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4518
timestamp 1713453518
transform 1 0 1604 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4519
timestamp 1713453518
transform 1 0 1292 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4520
timestamp 1713453518
transform 1 0 1132 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4521
timestamp 1713453518
transform 1 0 1092 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4522
timestamp 1713453518
transform 1 0 1276 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4523
timestamp 1713453518
transform 1 0 1252 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4524
timestamp 1713453518
transform 1 0 1244 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4525
timestamp 1713453518
transform 1 0 1188 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4526
timestamp 1713453518
transform 1 0 1244 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4527
timestamp 1713453518
transform 1 0 1172 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4528
timestamp 1713453518
transform 1 0 1652 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4529
timestamp 1713453518
transform 1 0 1644 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4530
timestamp 1713453518
transform 1 0 1556 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4531
timestamp 1713453518
transform 1 0 1532 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4532
timestamp 1713453518
transform 1 0 1532 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4533
timestamp 1713453518
transform 1 0 1244 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1713453518
transform 1 0 1852 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4535
timestamp 1713453518
transform 1 0 1012 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4536
timestamp 1713453518
transform 1 0 2812 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4537
timestamp 1713453518
transform 1 0 1804 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_4538
timestamp 1713453518
transform 1 0 1964 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4539
timestamp 1713453518
transform 1 0 1844 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4540
timestamp 1713453518
transform 1 0 1948 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4541
timestamp 1713453518
transform 1 0 1916 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4542
timestamp 1713453518
transform 1 0 2316 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4543
timestamp 1713453518
transform 1 0 2036 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4544
timestamp 1713453518
transform 1 0 3412 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4545
timestamp 1713453518
transform 1 0 3412 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4546
timestamp 1713453518
transform 1 0 3340 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4547
timestamp 1713453518
transform 1 0 2788 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4548
timestamp 1713453518
transform 1 0 2668 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4549
timestamp 1713453518
transform 1 0 2668 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4550
timestamp 1713453518
transform 1 0 2620 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4551
timestamp 1713453518
transform 1 0 2620 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4552
timestamp 1713453518
transform 1 0 2564 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4553
timestamp 1713453518
transform 1 0 2524 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4554
timestamp 1713453518
transform 1 0 2468 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4555
timestamp 1713453518
transform 1 0 2444 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4556
timestamp 1713453518
transform 1 0 2444 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4557
timestamp 1713453518
transform 1 0 2236 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4558
timestamp 1713453518
transform 1 0 1796 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4559
timestamp 1713453518
transform 1 0 2884 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4560
timestamp 1713453518
transform 1 0 2836 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4561
timestamp 1713453518
transform 1 0 2636 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4562
timestamp 1713453518
transform 1 0 2444 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4563
timestamp 1713453518
transform 1 0 1460 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4564
timestamp 1713453518
transform 1 0 1764 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4565
timestamp 1713453518
transform 1 0 1076 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4566
timestamp 1713453518
transform 1 0 2932 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4567
timestamp 1713453518
transform 1 0 2804 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4568
timestamp 1713453518
transform 1 0 2820 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4569
timestamp 1713453518
transform 1 0 2788 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_4570
timestamp 1713453518
transform 1 0 2756 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1713453518
transform 1 0 2732 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1713453518
transform 1 0 1412 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4573
timestamp 1713453518
transform 1 0 1308 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4574
timestamp 1713453518
transform 1 0 1236 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4575
timestamp 1713453518
transform 1 0 1100 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4576
timestamp 1713453518
transform 1 0 1252 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4577
timestamp 1713453518
transform 1 0 1196 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4578
timestamp 1713453518
transform 1 0 2052 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4579
timestamp 1713453518
transform 1 0 1900 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4580
timestamp 1713453518
transform 1 0 1900 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4581
timestamp 1713453518
transform 1 0 1084 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4582
timestamp 1713453518
transform 1 0 3284 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4583
timestamp 1713453518
transform 1 0 2012 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4584
timestamp 1713453518
transform 1 0 2324 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4585
timestamp 1713453518
transform 1 0 2100 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4586
timestamp 1713453518
transform 1 0 2604 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4587
timestamp 1713453518
transform 1 0 2532 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4588
timestamp 1713453518
transform 1 0 2500 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4589
timestamp 1713453518
transform 1 0 3292 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4590
timestamp 1713453518
transform 1 0 3236 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4591
timestamp 1713453518
transform 1 0 3108 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4592
timestamp 1713453518
transform 1 0 2588 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4593
timestamp 1713453518
transform 1 0 2076 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4594
timestamp 1713453518
transform 1 0 1812 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4595
timestamp 1713453518
transform 1 0 1764 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4596
timestamp 1713453518
transform 1 0 1084 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4597
timestamp 1713453518
transform 1 0 3420 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4598
timestamp 1713453518
transform 1 0 3300 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4599
timestamp 1713453518
transform 1 0 1212 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4600
timestamp 1713453518
transform 1 0 1180 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1713453518
transform 1 0 1284 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1713453518
transform 1 0 1204 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1713453518
transform 1 0 1204 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4604
timestamp 1713453518
transform 1 0 1132 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1713453518
transform 1 0 1140 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1713453518
transform 1 0 1092 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4607
timestamp 1713453518
transform 1 0 1092 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4608
timestamp 1713453518
transform 1 0 1068 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1713453518
transform 1 0 1052 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4610
timestamp 1713453518
transform 1 0 1052 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4611
timestamp 1713453518
transform 1 0 1212 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4612
timestamp 1713453518
transform 1 0 1180 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4613
timestamp 1713453518
transform 1 0 3372 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1713453518
transform 1 0 3364 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4615
timestamp 1713453518
transform 1 0 3228 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4616
timestamp 1713453518
transform 1 0 3228 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1713453518
transform 1 0 3148 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4618
timestamp 1713453518
transform 1 0 3148 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4619
timestamp 1713453518
transform 1 0 3132 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1713453518
transform 1 0 2276 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1713453518
transform 1 0 988 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1713453518
transform 1 0 3092 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1713453518
transform 1 0 2236 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4624
timestamp 1713453518
transform 1 0 2268 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4625
timestamp 1713453518
transform 1 0 2132 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1713453518
transform 1 0 2132 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4627
timestamp 1713453518
transform 1 0 2108 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1713453518
transform 1 0 2636 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4629
timestamp 1713453518
transform 1 0 2548 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4630
timestamp 1713453518
transform 1 0 2420 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4631
timestamp 1713453518
transform 1 0 3204 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1713453518
transform 1 0 3052 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1713453518
transform 1 0 2940 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4634
timestamp 1713453518
transform 1 0 2940 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1713453518
transform 1 0 2476 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4636
timestamp 1713453518
transform 1 0 2444 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4637
timestamp 1713453518
transform 1 0 2140 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4638
timestamp 1713453518
transform 1 0 1812 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4639
timestamp 1713453518
transform 1 0 1700 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4640
timestamp 1713453518
transform 1 0 1068 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4641
timestamp 1713453518
transform 1 0 3124 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4642
timestamp 1713453518
transform 1 0 3068 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4643
timestamp 1713453518
transform 1 0 3292 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4644
timestamp 1713453518
transform 1 0 3180 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4645
timestamp 1713453518
transform 1 0 3332 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4646
timestamp 1713453518
transform 1 0 3300 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4647
timestamp 1713453518
transform 1 0 3324 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4648
timestamp 1713453518
transform 1 0 3300 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4649
timestamp 1713453518
transform 1 0 1220 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4650
timestamp 1713453518
transform 1 0 1196 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4651
timestamp 1713453518
transform 1 0 1260 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4652
timestamp 1713453518
transform 1 0 1180 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4653
timestamp 1713453518
transform 1 0 1188 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4654
timestamp 1713453518
transform 1 0 1180 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4655
timestamp 1713453518
transform 1 0 1164 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4656
timestamp 1713453518
transform 1 0 1156 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4657
timestamp 1713453518
transform 1 0 1804 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4658
timestamp 1713453518
transform 1 0 1132 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4659
timestamp 1713453518
transform 1 0 3012 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4660
timestamp 1713453518
transform 1 0 1764 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4661
timestamp 1713453518
transform 1 0 2332 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4662
timestamp 1713453518
transform 1 0 1884 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4663
timestamp 1713453518
transform 1 0 2612 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4664
timestamp 1713453518
transform 1 0 2276 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4665
timestamp 1713453518
transform 1 0 1780 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4666
timestamp 1713453518
transform 1 0 2884 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4667
timestamp 1713453518
transform 1 0 2852 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4668
timestamp 1713453518
transform 1 0 2460 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4669
timestamp 1713453518
transform 1 0 2460 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4670
timestamp 1713453518
transform 1 0 2412 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4671
timestamp 1713453518
transform 1 0 1628 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4672
timestamp 1713453518
transform 1 0 1628 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4673
timestamp 1713453518
transform 1 0 1476 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4674
timestamp 1713453518
transform 1 0 2204 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4675
timestamp 1713453518
transform 1 0 1668 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4676
timestamp 1713453518
transform 1 0 3092 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1713453518
transform 1 0 3052 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4678
timestamp 1713453518
transform 1 0 3212 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4679
timestamp 1713453518
transform 1 0 3124 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4680
timestamp 1713453518
transform 1 0 1380 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4681
timestamp 1713453518
transform 1 0 1300 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4682
timestamp 1713453518
transform 1 0 2212 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4683
timestamp 1713453518
transform 1 0 1020 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4684
timestamp 1713453518
transform 1 0 2740 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4685
timestamp 1713453518
transform 1 0 2180 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4686
timestamp 1713453518
transform 1 0 2164 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4687
timestamp 1713453518
transform 1 0 2092 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1713453518
transform 1 0 2300 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4689
timestamp 1713453518
transform 1 0 2196 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4690
timestamp 1713453518
transform 1 0 3164 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4691
timestamp 1713453518
transform 1 0 2700 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4692
timestamp 1713453518
transform 1 0 2604 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4693
timestamp 1713453518
transform 1 0 2604 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4694
timestamp 1713453518
transform 1 0 2596 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4695
timestamp 1713453518
transform 1 0 2500 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4696
timestamp 1713453518
transform 1 0 2420 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4697
timestamp 1713453518
transform 1 0 2356 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1713453518
transform 1 0 2324 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4699
timestamp 1713453518
transform 1 0 2260 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4700
timestamp 1713453518
transform 1 0 2260 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4701
timestamp 1713453518
transform 1 0 2012 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4702
timestamp 1713453518
transform 1 0 2460 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4703
timestamp 1713453518
transform 1 0 2276 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4704
timestamp 1713453518
transform 1 0 1756 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4705
timestamp 1713453518
transform 1 0 2788 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4706
timestamp 1713453518
transform 1 0 2660 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4707
timestamp 1713453518
transform 1 0 2340 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1713453518
transform 1 0 1788 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4709
timestamp 1713453518
transform 1 0 2116 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4710
timestamp 1713453518
transform 1 0 2012 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4711
timestamp 1713453518
transform 1 0 1956 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4712
timestamp 1713453518
transform 1 0 1716 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4713
timestamp 1713453518
transform 1 0 1972 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4714
timestamp 1713453518
transform 1 0 1084 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4715
timestamp 1713453518
transform 1 0 1252 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4716
timestamp 1713453518
transform 1 0 1148 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4717
timestamp 1713453518
transform 1 0 1140 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4718
timestamp 1713453518
transform 1 0 1132 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_4719
timestamp 1713453518
transform 1 0 1132 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4720
timestamp 1713453518
transform 1 0 1084 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4721
timestamp 1713453518
transform 1 0 1196 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4722
timestamp 1713453518
transform 1 0 1148 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_4723
timestamp 1713453518
transform 1 0 1132 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4724
timestamp 1713453518
transform 1 0 1116 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4725
timestamp 1713453518
transform 1 0 1660 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4726
timestamp 1713453518
transform 1 0 1596 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1713453518
transform 1 0 1580 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1713453518
transform 1 0 1380 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4729
timestamp 1713453518
transform 1 0 2820 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1713453518
transform 1 0 2716 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1713453518
transform 1 0 2748 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4732
timestamp 1713453518
transform 1 0 2700 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4733
timestamp 1713453518
transform 1 0 1740 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4734
timestamp 1713453518
transform 1 0 1516 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4735
timestamp 1713453518
transform 1 0 1772 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4736
timestamp 1713453518
transform 1 0 1604 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4737
timestamp 1713453518
transform 1 0 1660 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1713453518
transform 1 0 1572 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1713453518
transform 1 0 1436 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4740
timestamp 1713453518
transform 1 0 1516 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4741
timestamp 1713453518
transform 1 0 1452 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4742
timestamp 1713453518
transform 1 0 2196 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4743
timestamp 1713453518
transform 1 0 1052 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4744
timestamp 1713453518
transform 1 0 2692 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4745
timestamp 1713453518
transform 1 0 2180 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4746
timestamp 1713453518
transform 1 0 2340 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4747
timestamp 1713453518
transform 1 0 2212 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4748
timestamp 1713453518
transform 1 0 3188 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4749
timestamp 1713453518
transform 1 0 2740 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4750
timestamp 1713453518
transform 1 0 2740 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4751
timestamp 1713453518
transform 1 0 2716 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4752
timestamp 1713453518
transform 1 0 2708 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4753
timestamp 1713453518
transform 1 0 2660 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4754
timestamp 1713453518
transform 1 0 2460 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4755
timestamp 1713453518
transform 1 0 2436 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4756
timestamp 1713453518
transform 1 0 2404 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4757
timestamp 1713453518
transform 1 0 2388 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4758
timestamp 1713453518
transform 1 0 2388 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4759
timestamp 1713453518
transform 1 0 2324 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4760
timestamp 1713453518
transform 1 0 1852 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4761
timestamp 1713453518
transform 1 0 2580 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4762
timestamp 1713453518
transform 1 0 2372 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4763
timestamp 1713453518
transform 1 0 1748 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4764
timestamp 1713453518
transform 1 0 2756 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4765
timestamp 1713453518
transform 1 0 2684 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4766
timestamp 1713453518
transform 1 0 2476 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4767
timestamp 1713453518
transform 1 0 1804 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4768
timestamp 1713453518
transform 1 0 2092 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4769
timestamp 1713453518
transform 1 0 1820 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_4770
timestamp 1713453518
transform 1 0 1772 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4771
timestamp 1713453518
transform 1 0 1668 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4772
timestamp 1713453518
transform 1 0 1796 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4773
timestamp 1713453518
transform 1 0 1156 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4774
timestamp 1713453518
transform 1 0 1628 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4775
timestamp 1713453518
transform 1 0 1620 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4776
timestamp 1713453518
transform 1 0 1580 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1713453518
transform 1 0 1580 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4778
timestamp 1713453518
transform 1 0 1436 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4779
timestamp 1713453518
transform 1 0 1428 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4780
timestamp 1713453518
transform 1 0 2820 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1713453518
transform 1 0 2676 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4782
timestamp 1713453518
transform 1 0 1740 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4783
timestamp 1713453518
transform 1 0 1516 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4784
timestamp 1713453518
transform 1 0 1764 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4785
timestamp 1713453518
transform 1 0 1692 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1713453518
transform 1 0 1636 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1713453518
transform 1 0 1596 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4788
timestamp 1713453518
transform 1 0 1660 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4789
timestamp 1713453518
transform 1 0 1636 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1713453518
transform 1 0 1700 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4791
timestamp 1713453518
transform 1 0 1668 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4792
timestamp 1713453518
transform 1 0 1660 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4793
timestamp 1713453518
transform 1 0 1588 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4794
timestamp 1713453518
transform 1 0 1452 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4795
timestamp 1713453518
transform 1 0 1356 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1713453518
transform 1 0 1564 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4797
timestamp 1713453518
transform 1 0 1460 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4798
timestamp 1713453518
transform 1 0 2308 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_4799
timestamp 1713453518
transform 1 0 1028 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_4800
timestamp 1713453518
transform 1 0 2788 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4801
timestamp 1713453518
transform 1 0 2276 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4802
timestamp 1713453518
transform 1 0 2244 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4803
timestamp 1713453518
transform 1 0 2124 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4804
timestamp 1713453518
transform 1 0 3084 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4805
timestamp 1713453518
transform 1 0 2532 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4806
timestamp 1713453518
transform 1 0 2492 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4807
timestamp 1713453518
transform 1 0 2404 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4808
timestamp 1713453518
transform 1 0 2404 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4809
timestamp 1713453518
transform 1 0 2340 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4810
timestamp 1713453518
transform 1 0 2308 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4811
timestamp 1713453518
transform 1 0 2220 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4812
timestamp 1713453518
transform 1 0 2204 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4813
timestamp 1713453518
transform 1 0 1852 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4814
timestamp 1713453518
transform 1 0 2516 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1713453518
transform 1 0 2332 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4816
timestamp 1713453518
transform 1 0 2188 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1713453518
transform 1 0 2188 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4818
timestamp 1713453518
transform 1 0 2028 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4819
timestamp 1713453518
transform 1 0 2028 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4820
timestamp 1713453518
transform 1 0 1660 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4821
timestamp 1713453518
transform 1 0 2948 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4822
timestamp 1713453518
transform 1 0 2884 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1713453518
transform 1 0 2884 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4824
timestamp 1713453518
transform 1 0 2572 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1713453518
transform 1 0 2572 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4826
timestamp 1713453518
transform 1 0 2540 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4827
timestamp 1713453518
transform 1 0 2428 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4828
timestamp 1713453518
transform 1 0 1780 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4829
timestamp 1713453518
transform 1 0 2068 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1713453518
transform 1 0 1860 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1713453518
transform 1 0 1812 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4832
timestamp 1713453518
transform 1 0 1652 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4833
timestamp 1713453518
transform 1 0 1820 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4834
timestamp 1713453518
transform 1 0 1068 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4835
timestamp 1713453518
transform 1 0 1628 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4836
timestamp 1713453518
transform 1 0 1604 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1713453518
transform 1 0 1604 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4838
timestamp 1713453518
transform 1 0 1540 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4839
timestamp 1713453518
transform 1 0 1540 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4840
timestamp 1713453518
transform 1 0 1452 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4841
timestamp 1713453518
transform 1 0 1452 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4842
timestamp 1713453518
transform 1 0 1380 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4843
timestamp 1713453518
transform 1 0 1340 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4844
timestamp 1713453518
transform 1 0 2932 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4845
timestamp 1713453518
transform 1 0 2756 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4846
timestamp 1713453518
transform 1 0 2732 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4847
timestamp 1713453518
transform 1 0 2668 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4848
timestamp 1713453518
transform 1 0 1700 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4849
timestamp 1713453518
transform 1 0 1636 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4850
timestamp 1713453518
transform 1 0 1764 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4851
timestamp 1713453518
transform 1 0 1676 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4852
timestamp 1713453518
transform 1 0 1620 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4853
timestamp 1713453518
transform 1 0 1596 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4854
timestamp 1713453518
transform 1 0 1724 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4855
timestamp 1713453518
transform 1 0 1724 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1713453518
transform 1 0 1700 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4857
timestamp 1713453518
transform 1 0 1620 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4858
timestamp 1713453518
transform 1 0 1580 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4859
timestamp 1713453518
transform 1 0 1564 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4860
timestamp 1713453518
transform 1 0 1564 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4861
timestamp 1713453518
transform 1 0 1564 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4862
timestamp 1713453518
transform 1 0 1292 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4863
timestamp 1713453518
transform 1 0 1276 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1713453518
transform 1 0 1556 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4865
timestamp 1713453518
transform 1 0 1508 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4866
timestamp 1713453518
transform 1 0 1820 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4867
timestamp 1713453518
transform 1 0 988 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4868
timestamp 1713453518
transform 1 0 2932 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4869
timestamp 1713453518
transform 1 0 1804 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4870
timestamp 1713453518
transform 1 0 2004 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4871
timestamp 1713453518
transform 1 0 1780 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4872
timestamp 1713453518
transform 1 0 1804 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4873
timestamp 1713453518
transform 1 0 1796 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4874
timestamp 1713453518
transform 1 0 1772 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4875
timestamp 1713453518
transform 1 0 1772 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4876
timestamp 1713453518
transform 1 0 1732 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4877
timestamp 1713453518
transform 1 0 1508 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4878
timestamp 1713453518
transform 1 0 1572 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4879
timestamp 1713453518
transform 1 0 1484 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4880
timestamp 1713453518
transform 1 0 2020 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4881
timestamp 1713453518
transform 1 0 2020 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4882
timestamp 1713453518
transform 1 0 1980 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4883
timestamp 1713453518
transform 1 0 1964 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4884
timestamp 1713453518
transform 1 0 1892 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4885
timestamp 1713453518
transform 1 0 1652 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4886
timestamp 1713453518
transform 1 0 2180 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4887
timestamp 1713453518
transform 1 0 2004 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_4888
timestamp 1713453518
transform 1 0 2060 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_4889
timestamp 1713453518
transform 1 0 1756 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_4890
timestamp 1713453518
transform 1 0 1732 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4891
timestamp 1713453518
transform 1 0 1316 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4892
timestamp 1713453518
transform 1 0 3124 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4893
timestamp 1713453518
transform 1 0 2852 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4894
timestamp 1713453518
transform 1 0 2844 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4895
timestamp 1713453518
transform 1 0 2772 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4896
timestamp 1713453518
transform 1 0 2508 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4897
timestamp 1713453518
transform 1 0 2228 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4898
timestamp 1713453518
transform 1 0 1836 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4899
timestamp 1713453518
transform 1 0 1836 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4900
timestamp 1713453518
transform 1 0 1780 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4901
timestamp 1713453518
transform 1 0 1660 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4902
timestamp 1713453518
transform 1 0 1356 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4903
timestamp 1713453518
transform 1 0 3012 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4904
timestamp 1713453518
transform 1 0 2980 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4905
timestamp 1713453518
transform 1 0 2596 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4906
timestamp 1713453518
transform 1 0 2500 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4907
timestamp 1713453518
transform 1 0 2380 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4908
timestamp 1713453518
transform 1 0 2300 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4909
timestamp 1713453518
transform 1 0 3044 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4910
timestamp 1713453518
transform 1 0 3012 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4911
timestamp 1713453518
transform 1 0 2820 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1713453518
transform 1 0 1524 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_4913
timestamp 1713453518
transform 1 0 2644 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4914
timestamp 1713453518
transform 1 0 2468 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4915
timestamp 1713453518
transform 1 0 2372 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4916
timestamp 1713453518
transform 1 0 2316 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4917
timestamp 1713453518
transform 1 0 2260 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4918
timestamp 1713453518
transform 1 0 2452 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4919
timestamp 1713453518
transform 1 0 2420 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4920
timestamp 1713453518
transform 1 0 2356 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4921
timestamp 1713453518
transform 1 0 1508 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1713453518
transform 1 0 1300 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4923
timestamp 1713453518
transform 1 0 1244 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4924
timestamp 1713453518
transform 1 0 1220 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4925
timestamp 1713453518
transform 1 0 1228 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4926
timestamp 1713453518
transform 1 0 1196 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4927
timestamp 1713453518
transform 1 0 1188 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_4928
timestamp 1713453518
transform 1 0 1132 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4929
timestamp 1713453518
transform 1 0 1116 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4930
timestamp 1713453518
transform 1 0 1436 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4931
timestamp 1713453518
transform 1 0 1404 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_4932
timestamp 1713453518
transform 1 0 1716 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4933
timestamp 1713453518
transform 1 0 1716 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4934
timestamp 1713453518
transform 1 0 1636 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4935
timestamp 1713453518
transform 1 0 1492 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4936
timestamp 1713453518
transform 1 0 1460 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4937
timestamp 1713453518
transform 1 0 1372 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1713453518
transform 1 0 1372 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4939
timestamp 1713453518
transform 1 0 1220 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4940
timestamp 1713453518
transform 1 0 2684 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4941
timestamp 1713453518
transform 1 0 2476 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4942
timestamp 1713453518
transform 1 0 2476 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4943
timestamp 1713453518
transform 1 0 2444 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1713453518
transform 1 0 2444 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4945
timestamp 1713453518
transform 1 0 2324 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1713453518
transform 1 0 1860 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4947
timestamp 1713453518
transform 1 0 1052 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4948
timestamp 1713453518
transform 1 0 2004 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4949
timestamp 1713453518
transform 1 0 1852 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4950
timestamp 1713453518
transform 1 0 2068 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4951
timestamp 1713453518
transform 1 0 1972 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4952
timestamp 1713453518
transform 1 0 2180 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4953
timestamp 1713453518
transform 1 0 1988 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4954
timestamp 1713453518
transform 1 0 1996 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4955
timestamp 1713453518
transform 1 0 1940 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4956
timestamp 1713453518
transform 1 0 1836 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4957
timestamp 1713453518
transform 1 0 1716 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4958
timestamp 1713453518
transform 1 0 1836 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1713453518
transform 1 0 1076 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4960
timestamp 1713453518
transform 1 0 3220 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4961
timestamp 1713453518
transform 1 0 2572 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4962
timestamp 1713453518
transform 1 0 2532 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4963
timestamp 1713453518
transform 1 0 2516 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4964
timestamp 1713453518
transform 1 0 2436 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4965
timestamp 1713453518
transform 1 0 1980 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4966
timestamp 1713453518
transform 1 0 1812 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4967
timestamp 1713453518
transform 1 0 2276 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4968
timestamp 1713453518
transform 1 0 2052 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_4969
timestamp 1713453518
transform 1 0 2036 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4970
timestamp 1713453518
transform 1 0 1956 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4971
timestamp 1713453518
transform 1 0 1924 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4972
timestamp 1713453518
transform 1 0 1732 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4973
timestamp 1713453518
transform 1 0 1524 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4974
timestamp 1713453518
transform 1 0 1940 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1713453518
transform 1 0 1412 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4976
timestamp 1713453518
transform 1 0 2484 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4977
timestamp 1713453518
transform 1 0 1956 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4978
timestamp 1713453518
transform 1 0 1956 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4979
timestamp 1713453518
transform 1 0 1892 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4980
timestamp 1713453518
transform 1 0 1852 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4981
timestamp 1713453518
transform 1 0 1420 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1713453518
transform 1 0 1268 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1713453518
transform 1 0 1172 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4984
timestamp 1713453518
transform 1 0 1148 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4985
timestamp 1713453518
transform 1 0 1204 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4986
timestamp 1713453518
transform 1 0 1156 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4987
timestamp 1713453518
transform 1 0 1156 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_4988
timestamp 1713453518
transform 1 0 1124 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4989
timestamp 1713453518
transform 1 0 1396 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4990
timestamp 1713453518
transform 1 0 1348 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4991
timestamp 1713453518
transform 1 0 1428 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4992
timestamp 1713453518
transform 1 0 1364 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4993
timestamp 1713453518
transform 1 0 1252 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_4994
timestamp 1713453518
transform 1 0 1828 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4995
timestamp 1713453518
transform 1 0 1812 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_4996
timestamp 1713453518
transform 1 0 1788 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4997
timestamp 1713453518
transform 1 0 1756 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4998
timestamp 1713453518
transform 1 0 1676 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_4999
timestamp 1713453518
transform 1 0 1452 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_5000
timestamp 1713453518
transform 1 0 1924 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5001
timestamp 1713453518
transform 1 0 1092 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5002
timestamp 1713453518
transform 1 0 2124 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5003
timestamp 1713453518
transform 1 0 1916 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5004
timestamp 1713453518
transform 1 0 2172 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_5005
timestamp 1713453518
transform 1 0 2116 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_5006
timestamp 1713453518
transform 1 0 2220 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5007
timestamp 1713453518
transform 1 0 2124 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5008
timestamp 1713453518
transform 1 0 2148 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5009
timestamp 1713453518
transform 1 0 2100 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5010
timestamp 1713453518
transform 1 0 2092 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5011
timestamp 1713453518
transform 1 0 1756 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5012
timestamp 1713453518
transform 1 0 1716 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5013
timestamp 1713453518
transform 1 0 1052 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5014
timestamp 1713453518
transform 1 0 3084 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5015
timestamp 1713453518
transform 1 0 2916 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5016
timestamp 1713453518
transform 1 0 2484 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_5017
timestamp 1713453518
transform 1 0 2460 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5018
timestamp 1713453518
transform 1 0 2404 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5019
timestamp 1713453518
transform 1 0 2404 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5020
timestamp 1713453518
transform 1 0 2292 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5021
timestamp 1713453518
transform 1 0 2268 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_5022
timestamp 1713453518
transform 1 0 2044 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_5023
timestamp 1713453518
transform 1 0 2044 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_5024
timestamp 1713453518
transform 1 0 1956 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_5025
timestamp 1713453518
transform 1 0 2340 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5026
timestamp 1713453518
transform 1 0 2148 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5027
timestamp 1713453518
transform 1 0 3220 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5028
timestamp 1713453518
transform 1 0 3180 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5029
timestamp 1713453518
transform 1 0 3148 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5030
timestamp 1713453518
transform 1 0 3124 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5031
timestamp 1713453518
transform 1 0 3092 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5032
timestamp 1713453518
transform 1 0 3092 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5033
timestamp 1713453518
transform 1 0 3212 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5034
timestamp 1713453518
transform 1 0 3164 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5035
timestamp 1713453518
transform 1 0 2084 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5036
timestamp 1713453518
transform 1 0 1956 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5037
timestamp 1713453518
transform 1 0 1948 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_5038
timestamp 1713453518
transform 1 0 1828 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1713453518
transform 1 0 1284 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_5040
timestamp 1713453518
transform 1 0 1908 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5041
timestamp 1713453518
transform 1 0 1436 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5042
timestamp 1713453518
transform 1 0 1444 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_5043
timestamp 1713453518
transform 1 0 1284 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_5044
timestamp 1713453518
transform 1 0 1428 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5045
timestamp 1713453518
transform 1 0 1372 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5046
timestamp 1713453518
transform 1 0 1436 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5047
timestamp 1713453518
transform 1 0 1396 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5048
timestamp 1713453518
transform 1 0 1260 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5049
timestamp 1713453518
transform 1 0 1260 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5050
timestamp 1713453518
transform 1 0 1100 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5051
timestamp 1713453518
transform 1 0 1332 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5052
timestamp 1713453518
transform 1 0 1236 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5053
timestamp 1713453518
transform 1 0 1196 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5054
timestamp 1713453518
transform 1 0 1940 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5055
timestamp 1713453518
transform 1 0 1924 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5056
timestamp 1713453518
transform 1 0 1828 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_5057
timestamp 1713453518
transform 1 0 1716 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_5058
timestamp 1713453518
transform 1 0 3324 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5059
timestamp 1713453518
transform 1 0 3284 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5060
timestamp 1713453518
transform 1 0 1620 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5061
timestamp 1713453518
transform 1 0 1460 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5062
timestamp 1713453518
transform 1 0 1860 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_5063
timestamp 1713453518
transform 1 0 1036 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_5064
timestamp 1713453518
transform 1 0 1860 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5065
timestamp 1713453518
transform 1 0 1836 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5066
timestamp 1713453518
transform 1 0 1996 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5067
timestamp 1713453518
transform 1 0 1836 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5068
timestamp 1713453518
transform 1 0 2156 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_5069
timestamp 1713453518
transform 1 0 1948 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_5070
timestamp 1713453518
transform 1 0 1924 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5071
timestamp 1713453518
transform 1 0 1820 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5072
timestamp 1713453518
transform 1 0 1764 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5073
timestamp 1713453518
transform 1 0 1716 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5074
timestamp 1713453518
transform 1 0 1812 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5075
timestamp 1713453518
transform 1 0 1020 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5076
timestamp 1713453518
transform 1 0 2092 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_5077
timestamp 1713453518
transform 1 0 2052 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_5078
timestamp 1713453518
transform 1 0 2388 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5079
timestamp 1713453518
transform 1 0 2132 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5080
timestamp 1713453518
transform 1 0 2044 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5081
timestamp 1713453518
transform 1 0 1884 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5082
timestamp 1713453518
transform 1 0 1868 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_5083
timestamp 1713453518
transform 1 0 1812 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_5084
timestamp 1713453518
transform 1 0 1812 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_5085
timestamp 1713453518
transform 1 0 1060 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_5086
timestamp 1713453518
transform 1 0 1860 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_5087
timestamp 1713453518
transform 1 0 1316 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_5088
timestamp 1713453518
transform 1 0 1332 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5089
timestamp 1713453518
transform 1 0 1268 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5090
timestamp 1713453518
transform 1 0 1284 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5091
timestamp 1713453518
transform 1 0 1172 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5092
timestamp 1713453518
transform 1 0 1172 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_5093
timestamp 1713453518
transform 1 0 1156 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5094
timestamp 1713453518
transform 1 0 1332 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5095
timestamp 1713453518
transform 1 0 1316 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5096
timestamp 1713453518
transform 1 0 1444 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5097
timestamp 1713453518
transform 1 0 1356 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5098
timestamp 1713453518
transform 1 0 1252 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1713453518
transform 1 0 1868 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_5100
timestamp 1713453518
transform 1 0 1836 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_5101
timestamp 1713453518
transform 1 0 1748 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5102
timestamp 1713453518
transform 1 0 1684 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_5103
timestamp 1713453518
transform 1 0 2084 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5104
timestamp 1713453518
transform 1 0 876 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5105
timestamp 1713453518
transform 1 0 2228 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5106
timestamp 1713453518
transform 1 0 2068 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5107
timestamp 1713453518
transform 1 0 2212 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5108
timestamp 1713453518
transform 1 0 1820 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5109
timestamp 1713453518
transform 1 0 2332 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_5110
timestamp 1713453518
transform 1 0 2228 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_5111
timestamp 1713453518
transform 1 0 1836 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_5112
timestamp 1713453518
transform 1 0 1628 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_5113
timestamp 1713453518
transform 1 0 1940 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_5114
timestamp 1713453518
transform 1 0 1828 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_5115
timestamp 1713453518
transform 1 0 1596 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_5116
timestamp 1713453518
transform 1 0 1548 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_5117
timestamp 1713453518
transform 1 0 1532 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_5118
timestamp 1713453518
transform 1 0 1956 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_5119
timestamp 1713453518
transform 1 0 1748 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_5120
timestamp 1713453518
transform 1 0 3300 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5121
timestamp 1713453518
transform 1 0 3236 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5122
timestamp 1713453518
transform 1 0 1364 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5123
timestamp 1713453518
transform 1 0 1316 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5124
timestamp 1713453518
transform 1 0 932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5125
timestamp 1713453518
transform 1 0 2924 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5126
timestamp 1713453518
transform 1 0 2852 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5127
timestamp 1713453518
transform 1 0 884 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5128
timestamp 1713453518
transform 1 0 868 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5129
timestamp 1713453518
transform 1 0 3172 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5130
timestamp 1713453518
transform 1 0 3156 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5131
timestamp 1713453518
transform 1 0 3252 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5132
timestamp 1713453518
transform 1 0 3180 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5133
timestamp 1713453518
transform 1 0 3188 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5134
timestamp 1713453518
transform 1 0 2564 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5135
timestamp 1713453518
transform 1 0 2620 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5136
timestamp 1713453518
transform 1 0 2516 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5137
timestamp 1713453518
transform 1 0 2508 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_5138
timestamp 1713453518
transform 1 0 2372 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_5139
timestamp 1713453518
transform 1 0 3308 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_5140
timestamp 1713453518
transform 1 0 3228 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_5141
timestamp 1713453518
transform 1 0 2380 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_5142
timestamp 1713453518
transform 1 0 2164 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_5143
timestamp 1713453518
transform 1 0 2228 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_5144
timestamp 1713453518
transform 1 0 2188 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_5145
timestamp 1713453518
transform 1 0 2068 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_5146
timestamp 1713453518
transform 1 0 1988 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_5147
timestamp 1713453518
transform 1 0 1964 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_5148
timestamp 1713453518
transform 1 0 1876 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_5149
timestamp 1713453518
transform 1 0 2116 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5150
timestamp 1713453518
transform 1 0 2052 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5151
timestamp 1713453518
transform 1 0 1980 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5152
timestamp 1713453518
transform 1 0 2084 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_5153
timestamp 1713453518
transform 1 0 1948 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_5154
timestamp 1713453518
transform 1 0 3140 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5155
timestamp 1713453518
transform 1 0 3028 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5156
timestamp 1713453518
transform 1 0 3044 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5157
timestamp 1713453518
transform 1 0 3012 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1713453518
transform 1 0 2860 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5159
timestamp 1713453518
transform 1 0 2860 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_5160
timestamp 1713453518
transform 1 0 2716 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5161
timestamp 1713453518
transform 1 0 2588 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5162
timestamp 1713453518
transform 1 0 1956 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5163
timestamp 1713453518
transform 1 0 3092 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5164
timestamp 1713453518
transform 1 0 3036 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5165
timestamp 1713453518
transform 1 0 2908 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5166
timestamp 1713453518
transform 1 0 2724 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5167
timestamp 1713453518
transform 1 0 2724 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5168
timestamp 1713453518
transform 1 0 2620 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5169
timestamp 1713453518
transform 1 0 2172 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_5170
timestamp 1713453518
transform 1 0 2996 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5171
timestamp 1713453518
transform 1 0 2900 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5172
timestamp 1713453518
transform 1 0 2684 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5173
timestamp 1713453518
transform 1 0 2612 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5174
timestamp 1713453518
transform 1 0 2140 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_5175
timestamp 1713453518
transform 1 0 2004 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_5176
timestamp 1713453518
transform 1 0 2164 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5177
timestamp 1713453518
transform 1 0 2044 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1713453518
transform 1 0 2036 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5179
timestamp 1713453518
transform 1 0 1908 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_5180
timestamp 1713453518
transform 1 0 1964 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5181
timestamp 1713453518
transform 1 0 1892 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5182
timestamp 1713453518
transform 1 0 2444 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_5183
timestamp 1713453518
transform 1 0 2116 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_5184
timestamp 1713453518
transform 1 0 636 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5185
timestamp 1713453518
transform 1 0 556 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5186
timestamp 1713453518
transform 1 0 660 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_5187
timestamp 1713453518
transform 1 0 612 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_5188
timestamp 1713453518
transform 1 0 436 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5189
timestamp 1713453518
transform 1 0 308 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5190
timestamp 1713453518
transform 1 0 820 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1713453518
transform 1 0 692 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5192
timestamp 1713453518
transform 1 0 636 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5193
timestamp 1713453518
transform 1 0 476 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5194
timestamp 1713453518
transform 1 0 356 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5195
timestamp 1713453518
transform 1 0 308 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5196
timestamp 1713453518
transform 1 0 324 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5197
timestamp 1713453518
transform 1 0 276 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5198
timestamp 1713453518
transform 1 0 292 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5199
timestamp 1713453518
transform 1 0 252 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5200
timestamp 1713453518
transform 1 0 812 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5201
timestamp 1713453518
transform 1 0 508 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5202
timestamp 1713453518
transform 1 0 756 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5203
timestamp 1713453518
transform 1 0 316 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5204
timestamp 1713453518
transform 1 0 812 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5205
timestamp 1713453518
transform 1 0 196 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5206
timestamp 1713453518
transform 1 0 340 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5207
timestamp 1713453518
transform 1 0 284 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5208
timestamp 1713453518
transform 1 0 356 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5209
timestamp 1713453518
transform 1 0 316 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5210
timestamp 1713453518
transform 1 0 348 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5211
timestamp 1713453518
transform 1 0 276 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5212
timestamp 1713453518
transform 1 0 348 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5213
timestamp 1713453518
transform 1 0 300 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5214
timestamp 1713453518
transform 1 0 516 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5215
timestamp 1713453518
transform 1 0 460 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5216
timestamp 1713453518
transform 1 0 284 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5217
timestamp 1713453518
transform 1 0 244 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5218
timestamp 1713453518
transform 1 0 356 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5219
timestamp 1713453518
transform 1 0 300 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5220
timestamp 1713453518
transform 1 0 412 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5221
timestamp 1713453518
transform 1 0 364 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5222
timestamp 1713453518
transform 1 0 348 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5223
timestamp 1713453518
transform 1 0 308 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5224
timestamp 1713453518
transform 1 0 476 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5225
timestamp 1713453518
transform 1 0 428 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5226
timestamp 1713453518
transform 1 0 332 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5227
timestamp 1713453518
transform 1 0 284 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5228
timestamp 1713453518
transform 1 0 316 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5229
timestamp 1713453518
transform 1 0 276 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5230
timestamp 1713453518
transform 1 0 252 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5231
timestamp 1713453518
transform 1 0 212 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5232
timestamp 1713453518
transform 1 0 372 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5233
timestamp 1713453518
transform 1 0 300 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5234
timestamp 1713453518
transform 1 0 596 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5235
timestamp 1713453518
transform 1 0 556 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_5236
timestamp 1713453518
transform 1 0 444 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5237
timestamp 1713453518
transform 1 0 444 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_5238
timestamp 1713453518
transform 1 0 252 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5239
timestamp 1713453518
transform 1 0 244 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_5240
timestamp 1713453518
transform 1 0 244 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_5241
timestamp 1713453518
transform 1 0 220 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5242
timestamp 1713453518
transform 1 0 196 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5243
timestamp 1713453518
transform 1 0 188 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_5244
timestamp 1713453518
transform 1 0 180 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5245
timestamp 1713453518
transform 1 0 580 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5246
timestamp 1713453518
transform 1 0 508 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5247
timestamp 1713453518
transform 1 0 468 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5248
timestamp 1713453518
transform 1 0 388 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5249
timestamp 1713453518
transform 1 0 532 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5250
timestamp 1713453518
transform 1 0 340 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5251
timestamp 1713453518
transform 1 0 332 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5252
timestamp 1713453518
transform 1 0 164 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5253
timestamp 1713453518
transform 1 0 372 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5254
timestamp 1713453518
transform 1 0 308 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5255
timestamp 1713453518
transform 1 0 492 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5256
timestamp 1713453518
transform 1 0 404 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5257
timestamp 1713453518
transform 1 0 364 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5258
timestamp 1713453518
transform 1 0 324 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5259
timestamp 1713453518
transform 1 0 148 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5260
timestamp 1713453518
transform 1 0 108 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_5261
timestamp 1713453518
transform 1 0 364 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1713453518
transform 1 0 124 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5263
timestamp 1713453518
transform 1 0 588 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5264
timestamp 1713453518
transform 1 0 356 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5265
timestamp 1713453518
transform 1 0 548 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5266
timestamp 1713453518
transform 1 0 492 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5267
timestamp 1713453518
transform 1 0 484 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_5268
timestamp 1713453518
transform 1 0 476 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5269
timestamp 1713453518
transform 1 0 412 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_5270
timestamp 1713453518
transform 1 0 412 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5271
timestamp 1713453518
transform 1 0 660 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1713453518
transform 1 0 660 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5273
timestamp 1713453518
transform 1 0 588 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5274
timestamp 1713453518
transform 1 0 556 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5275
timestamp 1713453518
transform 1 0 548 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5276
timestamp 1713453518
transform 1 0 468 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1713453518
transform 1 0 444 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_5278
timestamp 1713453518
transform 1 0 236 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_5279
timestamp 1713453518
transform 1 0 556 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1713453518
transform 1 0 452 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1713453518
transform 1 0 364 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5282
timestamp 1713453518
transform 1 0 308 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5283
timestamp 1713453518
transform 1 0 380 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5284
timestamp 1713453518
transform 1 0 340 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1713453518
transform 1 0 500 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1713453518
transform 1 0 500 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1713453518
transform 1 0 460 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_5288
timestamp 1713453518
transform 1 0 444 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5289
timestamp 1713453518
transform 1 0 572 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5290
timestamp 1713453518
transform 1 0 540 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5291
timestamp 1713453518
transform 1 0 652 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5292
timestamp 1713453518
transform 1 0 612 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5293
timestamp 1713453518
transform 1 0 428 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5294
timestamp 1713453518
transform 1 0 236 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1713453518
transform 1 0 676 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5296
timestamp 1713453518
transform 1 0 420 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5297
timestamp 1713453518
transform 1 0 644 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1713453518
transform 1 0 620 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1713453518
transform 1 0 588 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1713453518
transform 1 0 676 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1713453518
transform 1 0 604 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5302
timestamp 1713453518
transform 1 0 620 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1713453518
transform 1 0 604 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5304
timestamp 1713453518
transform 1 0 596 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5305
timestamp 1713453518
transform 1 0 548 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5306
timestamp 1713453518
transform 1 0 540 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5307
timestamp 1713453518
transform 1 0 460 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5308
timestamp 1713453518
transform 1 0 260 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5309
timestamp 1713453518
transform 1 0 620 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5310
timestamp 1713453518
transform 1 0 572 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5311
timestamp 1713453518
transform 1 0 572 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5312
timestamp 1713453518
transform 1 0 452 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5313
timestamp 1713453518
transform 1 0 628 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_5314
timestamp 1713453518
transform 1 0 556 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_5315
timestamp 1713453518
transform 1 0 420 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5316
timestamp 1713453518
transform 1 0 228 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5317
timestamp 1713453518
transform 1 0 580 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5318
timestamp 1713453518
transform 1 0 412 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5319
timestamp 1713453518
transform 1 0 580 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5320
timestamp 1713453518
transform 1 0 548 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5321
timestamp 1713453518
transform 1 0 396 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5322
timestamp 1713453518
transform 1 0 180 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5323
timestamp 1713453518
transform 1 0 676 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5324
timestamp 1713453518
transform 1 0 396 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5325
timestamp 1713453518
transform 1 0 684 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1713453518
transform 1 0 644 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5327
timestamp 1713453518
transform 1 0 652 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5328
timestamp 1713453518
transform 1 0 588 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1713453518
transform 1 0 588 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5330
timestamp 1713453518
transform 1 0 564 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5331
timestamp 1713453518
transform 1 0 612 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5332
timestamp 1713453518
transform 1 0 516 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5333
timestamp 1713453518
transform 1 0 516 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5334
timestamp 1713453518
transform 1 0 452 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5335
timestamp 1713453518
transform 1 0 716 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5336
timestamp 1713453518
transform 1 0 628 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5337
timestamp 1713453518
transform 1 0 620 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5338
timestamp 1713453518
transform 1 0 572 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5339
timestamp 1713453518
transform 1 0 572 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5340
timestamp 1713453518
transform 1 0 604 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5341
timestamp 1713453518
transform 1 0 428 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5342
timestamp 1713453518
transform 1 0 428 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5343
timestamp 1713453518
transform 1 0 412 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5344
timestamp 1713453518
transform 1 0 700 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5345
timestamp 1713453518
transform 1 0 692 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5346
timestamp 1713453518
transform 1 0 652 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5347
timestamp 1713453518
transform 1 0 644 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5348
timestamp 1713453518
transform 1 0 644 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5349
timestamp 1713453518
transform 1 0 620 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5350
timestamp 1713453518
transform 1 0 612 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5351
timestamp 1713453518
transform 1 0 740 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5352
timestamp 1713453518
transform 1 0 380 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5353
timestamp 1713453518
transform 1 0 740 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5354
timestamp 1713453518
transform 1 0 700 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5355
timestamp 1713453518
transform 1 0 348 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5356
timestamp 1713453518
transform 1 0 252 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5357
timestamp 1713453518
transform 1 0 644 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5358
timestamp 1713453518
transform 1 0 340 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5359
timestamp 1713453518
transform 1 0 676 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5360
timestamp 1713453518
transform 1 0 644 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5361
timestamp 1713453518
transform 1 0 428 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5362
timestamp 1713453518
transform 1 0 252 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5363
timestamp 1713453518
transform 1 0 692 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5364
timestamp 1713453518
transform 1 0 436 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5365
timestamp 1713453518
transform 1 0 708 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5366
timestamp 1713453518
transform 1 0 692 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5367
timestamp 1713453518
transform 1 0 724 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5368
timestamp 1713453518
transform 1 0 556 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5369
timestamp 1713453518
transform 1 0 540 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5370
timestamp 1713453518
transform 1 0 492 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5371
timestamp 1713453518
transform 1 0 780 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5372
timestamp 1713453518
transform 1 0 740 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5373
timestamp 1713453518
transform 1 0 676 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5374
timestamp 1713453518
transform 1 0 588 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5375
timestamp 1713453518
transform 1 0 748 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5376
timestamp 1713453518
transform 1 0 684 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5377
timestamp 1713453518
transform 1 0 652 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5378
timestamp 1713453518
transform 1 0 636 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5379
timestamp 1713453518
transform 1 0 628 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5380
timestamp 1713453518
transform 1 0 572 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5381
timestamp 1713453518
transform 1 0 572 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5382
timestamp 1713453518
transform 1 0 460 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5383
timestamp 1713453518
transform 1 0 260 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5384
timestamp 1713453518
transform 1 0 596 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1713453518
transform 1 0 460 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5386
timestamp 1713453518
transform 1 0 724 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5387
timestamp 1713453518
transform 1 0 644 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5388
timestamp 1713453518
transform 1 0 596 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5389
timestamp 1713453518
transform 1 0 572 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5390
timestamp 1713453518
transform 1 0 572 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5391
timestamp 1713453518
transform 1 0 460 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5392
timestamp 1713453518
transform 1 0 260 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5393
timestamp 1713453518
transform 1 0 700 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5394
timestamp 1713453518
transform 1 0 452 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5395
timestamp 1713453518
transform 1 0 460 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5396
timestamp 1713453518
transform 1 0 252 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5397
timestamp 1713453518
transform 1 0 748 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5398
timestamp 1713453518
transform 1 0 452 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5399
timestamp 1713453518
transform 1 0 500 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_5400
timestamp 1713453518
transform 1 0 420 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_5401
timestamp 1713453518
transform 1 0 708 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5402
timestamp 1713453518
transform 1 0 492 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5403
timestamp 1713453518
transform 1 0 756 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_5404
timestamp 1713453518
transform 1 0 724 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_5405
timestamp 1713453518
transform 1 0 596 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5406
timestamp 1713453518
transform 1 0 572 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5407
timestamp 1713453518
transform 1 0 788 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5408
timestamp 1713453518
transform 1 0 604 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5409
timestamp 1713453518
transform 1 0 524 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5410
timestamp 1713453518
transform 1 0 500 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5411
timestamp 1713453518
transform 1 0 476 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5412
timestamp 1713453518
transform 1 0 468 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5413
timestamp 1713453518
transform 1 0 460 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5414
timestamp 1713453518
transform 1 0 788 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5415
timestamp 1713453518
transform 1 0 692 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5416
timestamp 1713453518
transform 1 0 596 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5417
timestamp 1713453518
transform 1 0 252 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5418
timestamp 1713453518
transform 1 0 628 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5419
timestamp 1713453518
transform 1 0 604 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5420
timestamp 1713453518
transform 1 0 780 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5421
timestamp 1713453518
transform 1 0 780 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5422
timestamp 1713453518
transform 1 0 748 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5423
timestamp 1713453518
transform 1 0 676 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5424
timestamp 1713453518
transform 1 0 676 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5425
timestamp 1713453518
transform 1 0 612 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5426
timestamp 1713453518
transform 1 0 412 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5427
timestamp 1713453518
transform 1 0 244 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5428
timestamp 1713453518
transform 1 0 660 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5429
timestamp 1713453518
transform 1 0 396 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_5430
timestamp 1713453518
transform 1 0 684 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5431
timestamp 1713453518
transform 1 0 660 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5432
timestamp 1713453518
transform 1 0 444 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1713453518
transform 1 0 300 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5434
timestamp 1713453518
transform 1 0 772 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_5435
timestamp 1713453518
transform 1 0 436 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_5436
timestamp 1713453518
transform 1 0 788 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5437
timestamp 1713453518
transform 1 0 764 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5438
timestamp 1713453518
transform 1 0 500 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_5439
timestamp 1713453518
transform 1 0 300 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_5440
timestamp 1713453518
transform 1 0 740 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_5441
timestamp 1713453518
transform 1 0 492 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_5442
timestamp 1713453518
transform 1 0 780 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5443
timestamp 1713453518
transform 1 0 740 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5444
timestamp 1713453518
transform 1 0 604 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5445
timestamp 1713453518
transform 1 0 580 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5446
timestamp 1713453518
transform 1 0 716 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5447
timestamp 1713453518
transform 1 0 644 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5448
timestamp 1713453518
transform 1 0 540 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5449
timestamp 1713453518
transform 1 0 540 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5450
timestamp 1713453518
transform 1 0 508 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5451
timestamp 1713453518
transform 1 0 676 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5452
timestamp 1713453518
transform 1 0 636 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5453
timestamp 1713453518
transform 1 0 780 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5454
timestamp 1713453518
transform 1 0 772 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5455
timestamp 1713453518
transform 1 0 692 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5456
timestamp 1713453518
transform 1 0 692 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5457
timestamp 1713453518
transform 1 0 588 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5458
timestamp 1713453518
transform 1 0 564 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5459
timestamp 1713453518
transform 1 0 460 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5460
timestamp 1713453518
transform 1 0 252 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5461
timestamp 1713453518
transform 1 0 708 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5462
timestamp 1713453518
transform 1 0 460 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5463
timestamp 1713453518
transform 1 0 732 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5464
timestamp 1713453518
transform 1 0 660 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5465
timestamp 1713453518
transform 1 0 660 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5466
timestamp 1713453518
transform 1 0 628 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5467
timestamp 1713453518
transform 1 0 820 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1713453518
transform 1 0 652 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_5469
timestamp 1713453518
transform 1 0 836 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5470
timestamp 1713453518
transform 1 0 620 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5471
timestamp 1713453518
transform 1 0 836 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5472
timestamp 1713453518
transform 1 0 756 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5473
timestamp 1713453518
transform 1 0 860 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5474
timestamp 1713453518
transform 1 0 508 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5475
timestamp 1713453518
transform 1 0 868 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5476
timestamp 1713453518
transform 1 0 692 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5477
timestamp 1713453518
transform 1 0 708 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5478
timestamp 1713453518
transform 1 0 660 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5479
timestamp 1713453518
transform 1 0 596 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_5480
timestamp 1713453518
transform 1 0 588 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1713453518
transform 1 0 532 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5482
timestamp 1713453518
transform 1 0 532 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1713453518
transform 1 0 740 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5484
timestamp 1713453518
transform 1 0 556 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1713453518
transform 1 0 516 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1713453518
transform 1 0 668 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5487
timestamp 1713453518
transform 1 0 604 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5488
timestamp 1713453518
transform 1 0 556 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1713453518
transform 1 0 540 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1713453518
transform 1 0 532 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5491
timestamp 1713453518
transform 1 0 500 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5492
timestamp 1713453518
transform 1 0 420 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5493
timestamp 1713453518
transform 1 0 268 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5494
timestamp 1713453518
transform 1 0 548 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1713453518
transform 1 0 420 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5496
timestamp 1713453518
transform 1 0 596 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5497
timestamp 1713453518
transform 1 0 556 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5498
timestamp 1713453518
transform 1 0 532 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1713453518
transform 1 0 532 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5500
timestamp 1713453518
transform 1 0 220 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1713453518
transform 1 0 636 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5502
timestamp 1713453518
transform 1 0 548 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5503
timestamp 1713453518
transform 1 0 468 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1713453518
transform 1 0 220 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5505
timestamp 1713453518
transform 1 0 604 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5506
timestamp 1713453518
transform 1 0 460 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5507
timestamp 1713453518
transform 1 0 476 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5508
timestamp 1713453518
transform 1 0 236 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5509
timestamp 1713453518
transform 1 0 588 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1713453518
transform 1 0 468 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5511
timestamp 1713453518
transform 1 0 692 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5512
timestamp 1713453518
transform 1 0 588 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5513
timestamp 1713453518
transform 1 0 580 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5514
timestamp 1713453518
transform 1 0 540 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5515
timestamp 1713453518
transform 1 0 524 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5516
timestamp 1713453518
transform 1 0 524 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_5517
timestamp 1713453518
transform 1 0 772 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5518
timestamp 1713453518
transform 1 0 588 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_5519
timestamp 1713453518
transform 1 0 524 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5520
timestamp 1713453518
transform 1 0 500 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5521
timestamp 1713453518
transform 1 0 484 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5522
timestamp 1713453518
transform 1 0 484 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5523
timestamp 1713453518
transform 1 0 460 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5524
timestamp 1713453518
transform 1 0 428 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5525
timestamp 1713453518
transform 1 0 540 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5526
timestamp 1713453518
transform 1 0 500 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5527
timestamp 1713453518
transform 1 0 412 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5528
timestamp 1713453518
transform 1 0 604 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_5529
timestamp 1713453518
transform 1 0 540 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_5530
timestamp 1713453518
transform 1 0 604 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5531
timestamp 1713453518
transform 1 0 580 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5532
timestamp 1713453518
transform 1 0 676 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5533
timestamp 1713453518
transform 1 0 596 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5534
timestamp 1713453518
transform 1 0 612 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5535
timestamp 1713453518
transform 1 0 524 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5536
timestamp 1713453518
transform 1 0 524 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5537
timestamp 1713453518
transform 1 0 484 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5538
timestamp 1713453518
transform 1 0 492 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5539
timestamp 1713453518
transform 1 0 396 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_5540
timestamp 1713453518
transform 1 0 476 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5541
timestamp 1713453518
transform 1 0 380 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5542
timestamp 1713453518
transform 1 0 420 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_5543
timestamp 1713453518
transform 1 0 380 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1713453518
transform 1 0 508 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_5545
timestamp 1713453518
transform 1 0 460 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5546
timestamp 1713453518
transform 1 0 364 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_5547
timestamp 1713453518
transform 1 0 364 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5548
timestamp 1713453518
transform 1 0 468 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5549
timestamp 1713453518
transform 1 0 428 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5550
timestamp 1713453518
transform 1 0 532 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5551
timestamp 1713453518
transform 1 0 460 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5552
timestamp 1713453518
transform 1 0 508 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5553
timestamp 1713453518
transform 1 0 436 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5554
timestamp 1713453518
transform 1 0 660 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5555
timestamp 1713453518
transform 1 0 540 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5556
timestamp 1713453518
transform 1 0 516 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5557
timestamp 1713453518
transform 1 0 484 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5558
timestamp 1713453518
transform 1 0 676 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_5559
timestamp 1713453518
transform 1 0 652 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5560
timestamp 1713453518
transform 1 0 580 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5561
timestamp 1713453518
transform 1 0 492 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5562
timestamp 1713453518
transform 1 0 484 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_5563
timestamp 1713453518
transform 1 0 452 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5564
timestamp 1713453518
transform 1 0 316 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5565
timestamp 1713453518
transform 1 0 316 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5566
timestamp 1713453518
transform 1 0 284 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5567
timestamp 1713453518
transform 1 0 276 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5568
timestamp 1713453518
transform 1 0 268 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_5569
timestamp 1713453518
transform 1 0 268 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5570
timestamp 1713453518
transform 1 0 260 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5571
timestamp 1713453518
transform 1 0 260 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5572
timestamp 1713453518
transform 1 0 244 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5573
timestamp 1713453518
transform 1 0 244 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5574
timestamp 1713453518
transform 1 0 236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_5575
timestamp 1713453518
transform 1 0 164 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5576
timestamp 1713453518
transform 1 0 156 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5577
timestamp 1713453518
transform 1 0 564 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5578
timestamp 1713453518
transform 1 0 532 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5579
timestamp 1713453518
transform 1 0 500 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5580
timestamp 1713453518
transform 1 0 804 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5581
timestamp 1713453518
transform 1 0 772 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5582
timestamp 1713453518
transform 1 0 644 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5583
timestamp 1713453518
transform 1 0 604 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5584
timestamp 1713453518
transform 1 0 324 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5585
timestamp 1713453518
transform 1 0 212 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5586
timestamp 1713453518
transform 1 0 452 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5587
timestamp 1713453518
transform 1 0 356 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_5588
timestamp 1713453518
transform 1 0 220 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5589
timestamp 1713453518
transform 1 0 156 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5590
timestamp 1713453518
transform 1 0 236 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5591
timestamp 1713453518
transform 1 0 116 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_5592
timestamp 1713453518
transform 1 0 260 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5593
timestamp 1713453518
transform 1 0 148 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5594
timestamp 1713453518
transform 1 0 236 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5595
timestamp 1713453518
transform 1 0 116 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5596
timestamp 1713453518
transform 1 0 164 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5597
timestamp 1713453518
transform 1 0 116 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5598
timestamp 1713453518
transform 1 0 372 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5599
timestamp 1713453518
transform 1 0 260 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5600
timestamp 1713453518
transform 1 0 356 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5601
timestamp 1713453518
transform 1 0 252 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5602
timestamp 1713453518
transform 1 0 252 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5603
timestamp 1713453518
transform 1 0 148 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5604
timestamp 1713453518
transform 1 0 252 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5605
timestamp 1713453518
transform 1 0 140 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5606
timestamp 1713453518
transform 1 0 252 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5607
timestamp 1713453518
transform 1 0 148 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5608
timestamp 1713453518
transform 1 0 260 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5609
timestamp 1713453518
transform 1 0 148 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5610
timestamp 1713453518
transform 1 0 252 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5611
timestamp 1713453518
transform 1 0 116 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5612
timestamp 1713453518
transform 1 0 420 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5613
timestamp 1713453518
transform 1 0 316 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5614
timestamp 1713453518
transform 1 0 244 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5615
timestamp 1713453518
transform 1 0 140 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5616
timestamp 1713453518
transform 1 0 244 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5617
timestamp 1713453518
transform 1 0 140 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5618
timestamp 1713453518
transform 1 0 300 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5619
timestamp 1713453518
transform 1 0 148 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5620
timestamp 1713453518
transform 1 0 284 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5621
timestamp 1713453518
transform 1 0 164 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5622
timestamp 1713453518
transform 1 0 244 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5623
timestamp 1713453518
transform 1 0 132 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5624
timestamp 1713453518
transform 1 0 620 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5625
timestamp 1713453518
transform 1 0 572 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5626
timestamp 1713453518
transform 1 0 668 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5627
timestamp 1713453518
transform 1 0 564 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_5628
timestamp 1713453518
transform 1 0 468 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5629
timestamp 1713453518
transform 1 0 356 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5630
timestamp 1713453518
transform 1 0 268 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5631
timestamp 1713453518
transform 1 0 228 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5632
timestamp 1713453518
transform 1 0 220 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_5633
timestamp 1713453518
transform 1 0 132 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_5634
timestamp 1713453518
transform 1 0 212 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5635
timestamp 1713453518
transform 1 0 132 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5636
timestamp 1713453518
transform 1 0 236 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5637
timestamp 1713453518
transform 1 0 132 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5638
timestamp 1713453518
transform 1 0 572 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_5639
timestamp 1713453518
transform 1 0 516 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_5640
timestamp 1713453518
transform 1 0 1244 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5641
timestamp 1713453518
transform 1 0 1004 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5642
timestamp 1713453518
transform 1 0 1260 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5643
timestamp 1713453518
transform 1 0 1220 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5644
timestamp 1713453518
transform 1 0 1292 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_5645
timestamp 1713453518
transform 1 0 1260 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_5646
timestamp 1713453518
transform 1 0 724 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5647
timestamp 1713453518
transform 1 0 572 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5648
timestamp 1713453518
transform 1 0 420 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5649
timestamp 1713453518
transform 1 0 220 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5650
timestamp 1713453518
transform 1 0 460 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_5651
timestamp 1713453518
transform 1 0 204 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1713453518
transform 1 0 404 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_5653
timestamp 1713453518
transform 1 0 372 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_5654
timestamp 1713453518
transform 1 0 764 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5655
timestamp 1713453518
transform 1 0 700 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5656
timestamp 1713453518
transform 1 0 684 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_5657
timestamp 1713453518
transform 1 0 524 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_5658
timestamp 1713453518
transform 1 0 804 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_5659
timestamp 1713453518
transform 1 0 724 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1713453518
transform 1 0 1604 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_5661
timestamp 1713453518
transform 1 0 1580 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_5662
timestamp 1713453518
transform 1 0 1420 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_5663
timestamp 1713453518
transform 1 0 620 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5664
timestamp 1713453518
transform 1 0 412 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_5665
timestamp 1713453518
transform 1 0 404 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5666
timestamp 1713453518
transform 1 0 268 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_5667
timestamp 1713453518
transform 1 0 252 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5668
timestamp 1713453518
transform 1 0 1612 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5669
timestamp 1713453518
transform 1 0 1540 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5670
timestamp 1713453518
transform 1 0 1892 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5671
timestamp 1713453518
transform 1 0 1836 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5672
timestamp 1713453518
transform 1 0 1516 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5673
timestamp 1713453518
transform 1 0 1420 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_5674
timestamp 1713453518
transform 1 0 1548 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5675
timestamp 1713453518
transform 1 0 1516 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5676
timestamp 1713453518
transform 1 0 1556 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5677
timestamp 1713453518
transform 1 0 1468 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5678
timestamp 1713453518
transform 1 0 1428 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5679
timestamp 1713453518
transform 1 0 1380 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5680
timestamp 1713453518
transform 1 0 1444 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5681
timestamp 1713453518
transform 1 0 1388 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5682
timestamp 1713453518
transform 1 0 1420 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_5683
timestamp 1713453518
transform 1 0 1388 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_5684
timestamp 1713453518
transform 1 0 1436 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_5685
timestamp 1713453518
transform 1 0 1396 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_5686
timestamp 1713453518
transform 1 0 1492 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_5687
timestamp 1713453518
transform 1 0 1380 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_5688
timestamp 1713453518
transform 1 0 1412 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1713453518
transform 1 0 1364 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_5690
timestamp 1713453518
transform 1 0 3036 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5691
timestamp 1713453518
transform 1 0 2964 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1713453518
transform 1 0 2596 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1713453518
transform 1 0 2396 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1713453518
transform 1 0 2236 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5695
timestamp 1713453518
transform 1 0 2228 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_5696
timestamp 1713453518
transform 1 0 1636 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_5697
timestamp 1713453518
transform 1 0 1284 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_5698
timestamp 1713453518
transform 1 0 972 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_5699
timestamp 1713453518
transform 1 0 1316 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_5700
timestamp 1713453518
transform 1 0 1044 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_5701
timestamp 1713453518
transform 1 0 1708 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_5702
timestamp 1713453518
transform 1 0 1572 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1713453518
transform 1 0 1580 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5704
timestamp 1713453518
transform 1 0 948 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_5705
timestamp 1713453518
transform 1 0 948 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_5706
timestamp 1713453518
transform 1 0 772 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5707
timestamp 1713453518
transform 1 0 764 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1713453518
transform 1 0 724 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_5709
timestamp 1713453518
transform 1 0 724 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5710
timestamp 1713453518
transform 1 0 652 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1713453518
transform 1 0 620 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_5712
timestamp 1713453518
transform 1 0 868 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5713
timestamp 1713453518
transform 1 0 860 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1713453518
transform 1 0 836 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5715
timestamp 1713453518
transform 1 0 836 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1713453518
transform 1 0 812 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5717
timestamp 1713453518
transform 1 0 812 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5718
timestamp 1713453518
transform 1 0 780 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5719
timestamp 1713453518
transform 1 0 756 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5720
timestamp 1713453518
transform 1 0 756 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5721
timestamp 1713453518
transform 1 0 1412 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5722
timestamp 1713453518
transform 1 0 1076 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5723
timestamp 1713453518
transform 1 0 756 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5724
timestamp 1713453518
transform 1 0 756 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1713453518
transform 1 0 692 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5726
timestamp 1713453518
transform 1 0 652 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5727
timestamp 1713453518
transform 1 0 628 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5728
timestamp 1713453518
transform 1 0 1372 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5729
timestamp 1713453518
transform 1 0 1044 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5730
timestamp 1713453518
transform 1 0 1044 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5731
timestamp 1713453518
transform 1 0 996 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5732
timestamp 1713453518
transform 1 0 820 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1713453518
transform 1 0 812 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5734
timestamp 1713453518
transform 1 0 804 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5735
timestamp 1713453518
transform 1 0 788 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5736
timestamp 1713453518
transform 1 0 780 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5737
timestamp 1713453518
transform 1 0 780 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5738
timestamp 1713453518
transform 1 0 780 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5739
timestamp 1713453518
transform 1 0 676 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5740
timestamp 1713453518
transform 1 0 652 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_5741
timestamp 1713453518
transform 1 0 1300 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5742
timestamp 1713453518
transform 1 0 988 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5743
timestamp 1713453518
transform 1 0 748 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5744
timestamp 1713453518
transform 1 0 732 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1713453518
transform 1 0 652 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5746
timestamp 1713453518
transform 1 0 636 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5747
timestamp 1713453518
transform 1 0 636 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5748
timestamp 1713453518
transform 1 0 1276 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5749
timestamp 1713453518
transform 1 0 996 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1713453518
transform 1 0 932 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5751
timestamp 1713453518
transform 1 0 932 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1713453518
transform 1 0 892 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5753
timestamp 1713453518
transform 1 0 884 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5754
timestamp 1713453518
transform 1 0 740 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5755
timestamp 1713453518
transform 1 0 724 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5756
timestamp 1713453518
transform 1 0 940 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_5757
timestamp 1713453518
transform 1 0 772 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_5758
timestamp 1713453518
transform 1 0 692 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5759
timestamp 1713453518
transform 1 0 692 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_5760
timestamp 1713453518
transform 1 0 580 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5761
timestamp 1713453518
transform 1 0 524 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5762
timestamp 1713453518
transform 1 0 524 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_5763
timestamp 1713453518
transform 1 0 1468 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_5764
timestamp 1713453518
transform 1 0 1004 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_5765
timestamp 1713453518
transform 1 0 996 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_5766
timestamp 1713453518
transform 1 0 788 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_5767
timestamp 1713453518
transform 1 0 692 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_5768
timestamp 1713453518
transform 1 0 684 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_5769
timestamp 1713453518
transform 1 0 460 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_5770
timestamp 1713453518
transform 1 0 900 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5771
timestamp 1713453518
transform 1 0 748 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5772
timestamp 1713453518
transform 1 0 724 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5773
timestamp 1713453518
transform 1 0 572 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5774
timestamp 1713453518
transform 1 0 836 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5775
timestamp 1713453518
transform 1 0 772 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5776
timestamp 1713453518
transform 1 0 684 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5777
timestamp 1713453518
transform 1 0 588 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5778
timestamp 1713453518
transform 1 0 1236 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5779
timestamp 1713453518
transform 1 0 1084 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5780
timestamp 1713453518
transform 1 0 1060 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5781
timestamp 1713453518
transform 1 0 852 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_5782
timestamp 1713453518
transform 1 0 852 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5783
timestamp 1713453518
transform 1 0 748 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_5784
timestamp 1713453518
transform 1 0 676 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_5785
timestamp 1713453518
transform 1 0 676 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5786
timestamp 1713453518
transform 1 0 484 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_5787
timestamp 1713453518
transform 1 0 892 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5788
timestamp 1713453518
transform 1 0 844 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_5789
timestamp 1713453518
transform 1 0 844 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5790
timestamp 1713453518
transform 1 0 700 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5791
timestamp 1713453518
transform 1 0 628 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5792
timestamp 1713453518
transform 1 0 1412 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5793
timestamp 1713453518
transform 1 0 1324 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5794
timestamp 1713453518
transform 1 0 1052 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5795
timestamp 1713453518
transform 1 0 1044 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5796
timestamp 1713453518
transform 1 0 820 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5797
timestamp 1713453518
transform 1 0 684 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5798
timestamp 1713453518
transform 1 0 500 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5799
timestamp 1713453518
transform 1 0 492 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5800
timestamp 1713453518
transform 1 0 444 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5801
timestamp 1713453518
transform 1 0 1236 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5802
timestamp 1713453518
transform 1 0 1052 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5803
timestamp 1713453518
transform 1 0 940 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_5804
timestamp 1713453518
transform 1 0 1108 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5805
timestamp 1713453518
transform 1 0 1004 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_5806
timestamp 1713453518
transform 1 0 1212 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5807
timestamp 1713453518
transform 1 0 1132 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5808
timestamp 1713453518
transform 1 0 1084 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5809
timestamp 1713453518
transform 1 0 916 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5810
timestamp 1713453518
transform 1 0 1476 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5811
timestamp 1713453518
transform 1 0 1044 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5812
timestamp 1713453518
transform 1 0 924 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5813
timestamp 1713453518
transform 1 0 1268 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5814
timestamp 1713453518
transform 1 0 1052 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5815
timestamp 1713453518
transform 1 0 892 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5816
timestamp 1713453518
transform 1 0 1132 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5817
timestamp 1713453518
transform 1 0 1004 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5818
timestamp 1713453518
transform 1 0 868 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5819
timestamp 1713453518
transform 1 0 844 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5820
timestamp 1713453518
transform 1 0 812 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5821
timestamp 1713453518
transform 1 0 1092 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5822
timestamp 1713453518
transform 1 0 988 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5823
timestamp 1713453518
transform 1 0 988 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5824
timestamp 1713453518
transform 1 0 836 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5825
timestamp 1713453518
transform 1 0 812 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5826
timestamp 1713453518
transform 1 0 1540 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5827
timestamp 1713453518
transform 1 0 1052 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1713453518
transform 1 0 1052 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5829
timestamp 1713453518
transform 1 0 860 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5830
timestamp 1713453518
transform 1 0 844 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_5831
timestamp 1713453518
transform 1 0 844 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5832
timestamp 1713453518
transform 1 0 764 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_5833
timestamp 1713453518
transform 1 0 1052 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5834
timestamp 1713453518
transform 1 0 1004 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5835
timestamp 1713453518
transform 1 0 908 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5836
timestamp 1713453518
transform 1 0 884 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5837
timestamp 1713453518
transform 1 0 580 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_5838
timestamp 1713453518
transform 1 0 1460 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5839
timestamp 1713453518
transform 1 0 1052 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5840
timestamp 1713453518
transform 1 0 1028 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5841
timestamp 1713453518
transform 1 0 860 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_5842
timestamp 1713453518
transform 1 0 844 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5843
timestamp 1713453518
transform 1 0 732 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5844
timestamp 1713453518
transform 1 0 692 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5845
timestamp 1713453518
transform 1 0 1628 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5846
timestamp 1713453518
transform 1 0 956 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5847
timestamp 1713453518
transform 1 0 820 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5848
timestamp 1713453518
transform 1 0 788 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5849
timestamp 1713453518
transform 1 0 756 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5850
timestamp 1713453518
transform 1 0 732 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5851
timestamp 1713453518
transform 1 0 1020 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5852
timestamp 1713453518
transform 1 0 820 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5853
timestamp 1713453518
transform 1 0 812 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5854
timestamp 1713453518
transform 1 0 788 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5855
timestamp 1713453518
transform 1 0 788 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5856
timestamp 1713453518
transform 1 0 740 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5857
timestamp 1713453518
transform 1 0 740 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5858
timestamp 1713453518
transform 1 0 660 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5859
timestamp 1713453518
transform 1 0 644 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5860
timestamp 1713453518
transform 1 0 1292 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1713453518
transform 1 0 1004 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1713453518
transform 1 0 1004 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1713453518
transform 1 0 804 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5864
timestamp 1713453518
transform 1 0 804 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5865
timestamp 1713453518
transform 1 0 716 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5866
timestamp 1713453518
transform 1 0 564 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5867
timestamp 1713453518
transform 1 0 1212 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5868
timestamp 1713453518
transform 1 0 1076 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5869
timestamp 1713453518
transform 1 0 1044 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5870
timestamp 1713453518
transform 1 0 868 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5871
timestamp 1713453518
transform 1 0 1444 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5872
timestamp 1713453518
transform 1 0 1052 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5873
timestamp 1713453518
transform 1 0 908 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5874
timestamp 1713453518
transform 1 0 1412 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5875
timestamp 1713453518
transform 1 0 1052 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5876
timestamp 1713453518
transform 1 0 1052 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5877
timestamp 1713453518
transform 1 0 1004 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5878
timestamp 1713453518
transform 1 0 884 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5879
timestamp 1713453518
transform 1 0 1444 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5880
timestamp 1713453518
transform 1 0 996 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5881
timestamp 1713453518
transform 1 0 1476 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5882
timestamp 1713453518
transform 1 0 964 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5883
timestamp 1713453518
transform 1 0 964 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5884
timestamp 1713453518
transform 1 0 780 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5885
timestamp 1713453518
transform 1 0 732 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5886
timestamp 1713453518
transform 1 0 660 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5887
timestamp 1713453518
transform 1 0 1524 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5888
timestamp 1713453518
transform 1 0 1044 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5889
timestamp 1713453518
transform 1 0 868 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_5890
timestamp 1713453518
transform 1 0 708 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5891
timestamp 1713453518
transform 1 0 708 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_5892
timestamp 1713453518
transform 1 0 692 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5893
timestamp 1713453518
transform 1 0 564 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_5894
timestamp 1713453518
transform 1 0 836 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5895
timestamp 1713453518
transform 1 0 788 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5896
timestamp 1713453518
transform 1 0 692 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5897
timestamp 1713453518
transform 1 0 380 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5898
timestamp 1713453518
transform 1 0 380 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_5899
timestamp 1713453518
transform 1 0 356 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_5900
timestamp 1713453518
transform 1 0 700 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5901
timestamp 1713453518
transform 1 0 460 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_5902
timestamp 1713453518
transform 1 0 420 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_5903
timestamp 1713453518
transform 1 0 348 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_5904
timestamp 1713453518
transform 1 0 764 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5905
timestamp 1713453518
transform 1 0 732 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_5906
timestamp 1713453518
transform 1 0 732 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5907
timestamp 1713453518
transform 1 0 684 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_5908
timestamp 1713453518
transform 1 0 1548 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5909
timestamp 1713453518
transform 1 0 708 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_5910
timestamp 1713453518
transform 1 0 708 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_5911
timestamp 1713453518
transform 1 0 636 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5912
timestamp 1713453518
transform 1 0 596 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_5913
timestamp 1713453518
transform 1 0 1020 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5914
timestamp 1713453518
transform 1 0 940 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5915
timestamp 1713453518
transform 1 0 916 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5916
timestamp 1713453518
transform 1 0 700 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5917
timestamp 1713453518
transform 1 0 612 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5918
timestamp 1713453518
transform 1 0 548 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5919
timestamp 1713453518
transform 1 0 508 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5920
timestamp 1713453518
transform 1 0 404 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5921
timestamp 1713453518
transform 1 0 1044 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5922
timestamp 1713453518
transform 1 0 756 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5923
timestamp 1713453518
transform 1 0 524 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5924
timestamp 1713453518
transform 1 0 428 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_5925
timestamp 1713453518
transform 1 0 1068 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5926
timestamp 1713453518
transform 1 0 708 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5927
timestamp 1713453518
transform 1 0 628 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_5928
timestamp 1713453518
transform 1 0 1292 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_5929
timestamp 1713453518
transform 1 0 804 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5930
timestamp 1713453518
transform 1 0 620 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5931
timestamp 1713453518
transform 1 0 612 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_5932
timestamp 1713453518
transform 1 0 572 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_5933
timestamp 1713453518
transform 1 0 572 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5934
timestamp 1713453518
transform 1 0 340 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5935
timestamp 1713453518
transform 1 0 1044 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5936
timestamp 1713453518
transform 1 0 948 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5937
timestamp 1713453518
transform 1 0 684 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_5938
timestamp 1713453518
transform 1 0 684 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5939
timestamp 1713453518
transform 1 0 644 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_5940
timestamp 1713453518
transform 1 0 444 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_5941
timestamp 1713453518
transform 1 0 316 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_5942
timestamp 1713453518
transform 1 0 1116 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5943
timestamp 1713453518
transform 1 0 748 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5944
timestamp 1713453518
transform 1 0 564 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_5945
timestamp 1713453518
transform 1 0 436 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5946
timestamp 1713453518
transform 1 0 420 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5947
timestamp 1713453518
transform 1 0 1084 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5948
timestamp 1713453518
transform 1 0 804 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5949
timestamp 1713453518
transform 1 0 660 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5950
timestamp 1713453518
transform 1 0 388 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5951
timestamp 1713453518
transform 1 0 652 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5952
timestamp 1713453518
transform 1 0 652 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5953
timestamp 1713453518
transform 1 0 580 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5954
timestamp 1713453518
transform 1 0 428 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5955
timestamp 1713453518
transform 1 0 1052 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5956
timestamp 1713453518
transform 1 0 724 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5957
timestamp 1713453518
transform 1 0 708 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5958
timestamp 1713453518
transform 1 0 692 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5959
timestamp 1713453518
transform 1 0 652 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5960
timestamp 1713453518
transform 1 0 508 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5961
timestamp 1713453518
transform 1 0 1044 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5962
timestamp 1713453518
transform 1 0 748 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5963
timestamp 1713453518
transform 1 0 700 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5964
timestamp 1713453518
transform 1 0 700 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5965
timestamp 1713453518
transform 1 0 700 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5966
timestamp 1713453518
transform 1 0 516 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5967
timestamp 1713453518
transform 1 0 516 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5968
timestamp 1713453518
transform 1 0 428 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5969
timestamp 1713453518
transform 1 0 404 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5970
timestamp 1713453518
transform 1 0 1108 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5971
timestamp 1713453518
transform 1 0 764 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5972
timestamp 1713453518
transform 1 0 740 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5973
timestamp 1713453518
transform 1 0 668 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5974
timestamp 1713453518
transform 1 0 420 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5975
timestamp 1713453518
transform 1 0 420 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5976
timestamp 1713453518
transform 1 0 1092 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5977
timestamp 1713453518
transform 1 0 988 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5978
timestamp 1713453518
transform 1 0 708 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5979
timestamp 1713453518
transform 1 0 652 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5980
timestamp 1713453518
transform 1 0 644 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5981
timestamp 1713453518
transform 1 0 636 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5982
timestamp 1713453518
transform 1 0 628 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5983
timestamp 1713453518
transform 1 0 620 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5984
timestamp 1713453518
transform 1 0 612 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5985
timestamp 1713453518
transform 1 0 428 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5986
timestamp 1713453518
transform 1 0 428 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5987
timestamp 1713453518
transform 1 0 1108 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5988
timestamp 1713453518
transform 1 0 1068 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5989
timestamp 1713453518
transform 1 0 668 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5990
timestamp 1713453518
transform 1 0 404 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5991
timestamp 1713453518
transform 1 0 396 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5992
timestamp 1713453518
transform 1 0 1204 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5993
timestamp 1713453518
transform 1 0 1108 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5994
timestamp 1713453518
transform 1 0 804 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_5995
timestamp 1713453518
transform 1 0 764 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_5996
timestamp 1713453518
transform 1 0 764 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5997
timestamp 1713453518
transform 1 0 748 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5998
timestamp 1713453518
transform 1 0 660 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5999
timestamp 1713453518
transform 1 0 652 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_6000
timestamp 1713453518
transform 1 0 380 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_6001
timestamp 1713453518
transform 1 0 1116 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_6002
timestamp 1713453518
transform 1 0 1020 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_6003
timestamp 1713453518
transform 1 0 788 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_6004
timestamp 1713453518
transform 1 0 788 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_6005
timestamp 1713453518
transform 1 0 780 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6006
timestamp 1713453518
transform 1 0 756 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6007
timestamp 1713453518
transform 1 0 700 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_6008
timestamp 1713453518
transform 1 0 444 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_6009
timestamp 1713453518
transform 1 0 444 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_6010
timestamp 1713453518
transform 1 0 652 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6011
timestamp 1713453518
transform 1 0 524 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6012
timestamp 1713453518
transform 1 0 524 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_6013
timestamp 1713453518
transform 1 0 524 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_6014
timestamp 1713453518
transform 1 0 476 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_6015
timestamp 1713453518
transform 1 0 1108 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_6016
timestamp 1713453518
transform 1 0 836 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_6017
timestamp 1713453518
transform 1 0 836 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_6018
timestamp 1713453518
transform 1 0 836 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_6019
timestamp 1713453518
transform 1 0 820 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_6020
timestamp 1713453518
transform 1 0 820 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_6021
timestamp 1713453518
transform 1 0 796 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6022
timestamp 1713453518
transform 1 0 796 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_6023
timestamp 1713453518
transform 1 0 780 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6024
timestamp 1713453518
transform 1 0 468 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_6025
timestamp 1713453518
transform 1 0 1044 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6026
timestamp 1713453518
transform 1 0 820 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6027
timestamp 1713453518
transform 1 0 740 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6028
timestamp 1713453518
transform 1 0 652 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6029
timestamp 1713453518
transform 1 0 468 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6030
timestamp 1713453518
transform 1 0 76 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_6031
timestamp 1713453518
transform 1 0 76 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_6032
timestamp 1713453518
transform 1 0 1116 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_6033
timestamp 1713453518
transform 1 0 884 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_6034
timestamp 1713453518
transform 1 0 876 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_6035
timestamp 1713453518
transform 1 0 708 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_6036
timestamp 1713453518
transform 1 0 652 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_6037
timestamp 1713453518
transform 1 0 508 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_6038
timestamp 1713453518
transform 1 0 508 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_6039
timestamp 1713453518
transform 1 0 1108 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_6040
timestamp 1713453518
transform 1 0 876 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_6041
timestamp 1713453518
transform 1 0 604 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_6042
timestamp 1713453518
transform 1 0 604 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6043
timestamp 1713453518
transform 1 0 548 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6044
timestamp 1713453518
transform 1 0 348 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6045
timestamp 1713453518
transform 1 0 348 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6046
timestamp 1713453518
transform 1 0 1124 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_6047
timestamp 1713453518
transform 1 0 844 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_6048
timestamp 1713453518
transform 1 0 700 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_6049
timestamp 1713453518
transform 1 0 652 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_6050
timestamp 1713453518
transform 1 0 628 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_6051
timestamp 1713453518
transform 1 0 628 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_6052
timestamp 1713453518
transform 1 0 612 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_6053
timestamp 1713453518
transform 1 0 420 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_6054
timestamp 1713453518
transform 1 0 1068 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6055
timestamp 1713453518
transform 1 0 876 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6056
timestamp 1713453518
transform 1 0 772 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6057
timestamp 1713453518
transform 1 0 716 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6058
timestamp 1713453518
transform 1 0 660 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_6059
timestamp 1713453518
transform 1 0 620 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_6060
timestamp 1713453518
transform 1 0 620 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6061
timestamp 1713453518
transform 1 0 452 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6062
timestamp 1713453518
transform 1 0 1092 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_6063
timestamp 1713453518
transform 1 0 900 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_6064
timestamp 1713453518
transform 1 0 756 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_6065
timestamp 1713453518
transform 1 0 756 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_6066
timestamp 1713453518
transform 1 0 692 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_6067
timestamp 1713453518
transform 1 0 580 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6068
timestamp 1713453518
transform 1 0 508 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_6069
timestamp 1713453518
transform 1 0 508 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_6070
timestamp 1713453518
transform 1 0 460 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6071
timestamp 1713453518
transform 1 0 460 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_6072
timestamp 1713453518
transform 1 0 884 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6073
timestamp 1713453518
transform 1 0 780 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6074
timestamp 1713453518
transform 1 0 652 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6075
timestamp 1713453518
transform 1 0 468 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6076
timestamp 1713453518
transform 1 0 1140 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6077
timestamp 1713453518
transform 1 0 860 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6078
timestamp 1713453518
transform 1 0 788 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6079
timestamp 1713453518
transform 1 0 740 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6080
timestamp 1713453518
transform 1 0 724 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6081
timestamp 1713453518
transform 1 0 724 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6082
timestamp 1713453518
transform 1 0 684 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6083
timestamp 1713453518
transform 1 0 668 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6084
timestamp 1713453518
transform 1 0 1036 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6085
timestamp 1713453518
transform 1 0 780 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6086
timestamp 1713453518
transform 1 0 756 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6087
timestamp 1713453518
transform 1 0 756 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_6088
timestamp 1713453518
transform 1 0 724 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_6089
timestamp 1713453518
transform 1 0 668 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_6090
timestamp 1713453518
transform 1 0 636 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_6091
timestamp 1713453518
transform 1 0 1100 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_6092
timestamp 1713453518
transform 1 0 980 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_6093
timestamp 1713453518
transform 1 0 980 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_6094
timestamp 1713453518
transform 1 0 772 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_6095
timestamp 1713453518
transform 1 0 764 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_6096
timestamp 1713453518
transform 1 0 748 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_6097
timestamp 1713453518
transform 1 0 748 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6098
timestamp 1713453518
transform 1 0 676 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6099
timestamp 1713453518
transform 1 0 564 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6100
timestamp 1713453518
transform 1 0 428 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6101
timestamp 1713453518
transform 1 0 1220 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_6102
timestamp 1713453518
transform 1 0 1204 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_6103
timestamp 1713453518
transform 1 0 1092 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_6104
timestamp 1713453518
transform 1 0 1092 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_6105
timestamp 1713453518
transform 1 0 964 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_6106
timestamp 1713453518
transform 1 0 860 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_6107
timestamp 1713453518
transform 1 0 588 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_6108
timestamp 1713453518
transform 1 0 1172 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6109
timestamp 1713453518
transform 1 0 1156 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6110
timestamp 1713453518
transform 1 0 852 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_6111
timestamp 1713453518
transform 1 0 732 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_6112
timestamp 1713453518
transform 1 0 732 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6113
timestamp 1713453518
transform 1 0 732 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6114
timestamp 1713453518
transform 1 0 676 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6115
timestamp 1713453518
transform 1 0 500 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6116
timestamp 1713453518
transform 1 0 1180 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6117
timestamp 1713453518
transform 1 0 1052 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6118
timestamp 1713453518
transform 1 0 1052 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_6119
timestamp 1713453518
transform 1 0 836 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_6120
timestamp 1713453518
transform 1 0 788 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_6121
timestamp 1713453518
transform 1 0 788 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_6122
timestamp 1713453518
transform 1 0 668 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6123
timestamp 1713453518
transform 1 0 524 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6124
timestamp 1713453518
transform 1 0 2780 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_6125
timestamp 1713453518
transform 1 0 1372 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_6126
timestamp 1713453518
transform 1 0 1276 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_6127
timestamp 1713453518
transform 1 0 1268 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_6128
timestamp 1713453518
transform 1 0 1108 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_6129
timestamp 1713453518
transform 1 0 892 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_6130
timestamp 1713453518
transform 1 0 892 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_6131
timestamp 1713453518
transform 1 0 604 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_6132
timestamp 1713453518
transform 1 0 508 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_6133
timestamp 1713453518
transform 1 0 452 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_6134
timestamp 1713453518
transform 1 0 668 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6135
timestamp 1713453518
transform 1 0 76 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6136
timestamp 1713453518
transform 1 0 76 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_6137
timestamp 1713453518
transform 1 0 1268 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_6138
timestamp 1713453518
transform 1 0 1036 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_6139
timestamp 1713453518
transform 1 0 1036 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_6140
timestamp 1713453518
transform 1 0 684 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_6141
timestamp 1713453518
transform 1 0 380 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_6142
timestamp 1713453518
transform 1 0 372 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_6143
timestamp 1713453518
transform 1 0 348 0 1 915
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1713453518
transform 1 0 2744 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1713453518
transform 1 0 2592 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1713453518
transform 1 0 2760 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1713453518
transform 1 0 2296 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1713453518
transform 1 0 2240 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1713453518
transform 1 0 2240 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1713453518
transform 1 0 1872 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1713453518
transform 1 0 2400 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1713453518
transform 1 0 2120 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1713453518
transform 1 0 3416 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1713453518
transform 1 0 2536 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1713453518
transform 1 0 2640 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1713453518
transform 1 0 1656 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1713453518
transform 1 0 1200 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1713453518
transform 1 0 1576 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1713453518
transform 1 0 1184 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1713453518
transform 1 0 1840 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1713453518
transform 1 0 1248 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1713453518
transform 1 0 1920 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1713453518
transform 1 0 1992 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1713453518
transform 1 0 2816 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1713453518
transform 1 0 2744 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1713453518
transform 1 0 2456 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1713453518
transform 1 0 2528 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1713453518
transform 1 0 1104 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1713453518
transform 1 0 3128 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1713453518
transform 1 0 3152 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1713453518
transform 1 0 2584 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1713453518
transform 1 0 2800 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1713453518
transform 1 0 2416 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1713453518
transform 1 0 1200 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1713453518
transform 1 0 1152 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1713453518
transform 1 0 3320 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1713453518
transform 1 0 3344 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1713453518
transform 1 0 3176 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1713453518
transform 1 0 2576 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1713453518
transform 1 0 2824 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1713453518
transform 1 0 2256 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1713453518
transform 1 0 1240 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1713453518
transform 1 0 1096 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1713453518
transform 1 0 3120 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1713453518
transform 1 0 3344 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1713453518
transform 1 0 3368 0 -1 3370
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1713453518
transform 1 0 3208 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1713453518
transform 1 0 2472 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1713453518
transform 1 0 2640 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1713453518
transform 1 0 3216 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1713453518
transform 1 0 1528 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1713453518
transform 1 0 3280 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1713453518
transform 1 0 3304 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1713453518
transform 1 0 3216 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1713453518
transform 1 0 2072 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1713453518
transform 1 0 2568 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1713453518
transform 1 0 1480 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1713453518
transform 1 0 3232 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1713453518
transform 1 0 1624 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1713453518
transform 1 0 3312 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1713453518
transform 1 0 3288 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1713453518
transform 1 0 1584 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1713453518
transform 1 0 1296 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1713453518
transform 1 0 3104 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1713453518
transform 1 0 1832 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1713453518
transform 1 0 2512 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1713453518
transform 1 0 1504 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1713453518
transform 1 0 3256 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1713453518
transform 1 0 1520 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1713453518
transform 1 0 3392 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1713453518
transform 1 0 3328 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1713453518
transform 1 0 1408 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1713453518
transform 1 0 1128 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1713453518
transform 1 0 1728 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1713453518
transform 1 0 2056 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1713453518
transform 1 0 1488 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1713453518
transform 1 0 2856 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1713453518
transform 1 0 2864 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1713453518
transform 1 0 3000 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1713453518
transform 1 0 1704 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1713453518
transform 1 0 1360 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1713453518
transform 1 0 1720 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1713453518
transform 1 0 3192 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1713453518
transform 1 0 2080 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1713453518
transform 1 0 1552 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1713453518
transform 1 0 2792 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1713453518
transform 1 0 2912 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1713453518
transform 1 0 2872 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1713453518
transform 1 0 1696 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1713453518
transform 1 0 1200 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1713453518
transform 1 0 1880 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_88
timestamp 1713453518
transform 1 0 3120 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_89
timestamp 1713453518
transform 1 0 2136 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1713453518
transform 1 0 2440 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_91
timestamp 1713453518
transform 1 0 1568 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_92
timestamp 1713453518
transform 1 0 3000 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1713453518
transform 1 0 3296 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_94
timestamp 1713453518
transform 1 0 3056 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_95
timestamp 1713453518
transform 1 0 1384 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1713453518
transform 1 0 1248 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_97
timestamp 1713453518
transform 1 0 2904 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_98
timestamp 1713453518
transform 1 0 1856 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1713453518
transform 1 0 2688 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_100
timestamp 1713453518
transform 1 0 1544 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_101
timestamp 1713453518
transform 1 0 1352 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1713453518
transform 1 0 3288 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_103
timestamp 1713453518
transform 1 0 3320 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1713453518
transform 1 0 3296 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1713453518
transform 1 0 3016 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_106
timestamp 1713453518
transform 1 0 3096 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_107
timestamp 1713453518
transform 1 0 2448 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_108
timestamp 1713453518
transform 1 0 2696 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_109
timestamp 1713453518
transform 1 0 1568 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_110
timestamp 1713453518
transform 1 0 1168 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_111
timestamp 1713453518
transform 1 0 3240 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_112
timestamp 1713453518
transform 1 0 3304 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1713453518
transform 1 0 3328 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_114
timestamp 1713453518
transform 1 0 1168 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_115
timestamp 1713453518
transform 1 0 3280 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_116
timestamp 1713453518
transform 1 0 2424 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_117
timestamp 1713453518
transform 1 0 2584 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1713453518
transform 1 0 3200 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_119
timestamp 1713453518
transform 1 0 1824 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_120
timestamp 1713453518
transform 1 0 3296 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1713453518
transform 1 0 3248 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_122
timestamp 1713453518
transform 1 0 3264 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1713453518
transform 1 0 3272 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1713453518
transform 1 0 2248 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1713453518
transform 1 0 1696 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_126
timestamp 1713453518
transform 1 0 3008 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_127
timestamp 1713453518
transform 1 0 3280 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_128
timestamp 1713453518
transform 1 0 3320 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_129
timestamp 1713453518
transform 1 0 1624 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_130
timestamp 1713453518
transform 1 0 1264 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_131
timestamp 1713453518
transform 1 0 2992 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_132
timestamp 1713453518
transform 1 0 2280 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_133
timestamp 1713453518
transform 1 0 2560 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_134
timestamp 1713453518
transform 1 0 1768 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_135
timestamp 1713453518
transform 1 0 3296 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_136
timestamp 1713453518
transform 1 0 1704 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_137
timestamp 1713453518
transform 1 0 3256 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_138
timestamp 1713453518
transform 1 0 3296 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_139
timestamp 1713453518
transform 1 0 1728 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_140
timestamp 1713453518
transform 1 0 1160 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_141
timestamp 1713453518
transform 1 0 3200 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_142
timestamp 1713453518
transform 1 0 3248 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_143
timestamp 1713453518
transform 1 0 2288 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_144
timestamp 1713453518
transform 1 0 2392 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_145
timestamp 1713453518
transform 1 0 1680 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_146
timestamp 1713453518
transform 1 0 3040 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_147
timestamp 1713453518
transform 1 0 1680 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_148
timestamp 1713453518
transform 1 0 3176 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_149
timestamp 1713453518
transform 1 0 3248 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_150
timestamp 1713453518
transform 1 0 1744 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_151
timestamp 1713453518
transform 1 0 1368 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_152
timestamp 1713453518
transform 1 0 3200 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_153
timestamp 1713453518
transform 1 0 1936 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_154
timestamp 1713453518
transform 1 0 2304 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_155
timestamp 1713453518
transform 1 0 1656 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_156
timestamp 1713453518
transform 1 0 2672 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_157
timestamp 1713453518
transform 1 0 1680 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_158
timestamp 1713453518
transform 1 0 2832 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_159
timestamp 1713453518
transform 1 0 2960 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_160
timestamp 1713453518
transform 1 0 1584 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_161
timestamp 1713453518
transform 1 0 1192 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_162
timestamp 1713453518
transform 1 0 2688 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_163
timestamp 1713453518
transform 1 0 3104 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_164
timestamp 1713453518
transform 1 0 1968 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_165
timestamp 1713453518
transform 1 0 2240 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_166
timestamp 1713453518
transform 1 0 1648 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_167
timestamp 1713453518
transform 1 0 2800 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_168
timestamp 1713453518
transform 1 0 2864 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_169
timestamp 1713453518
transform 1 0 2816 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_170
timestamp 1713453518
transform 1 0 1304 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_171
timestamp 1713453518
transform 1 0 1232 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_172
timestamp 1713453518
transform 1 0 2688 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_173
timestamp 1713453518
transform 1 0 3128 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_174
timestamp 1713453518
transform 1 0 2048 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_175
timestamp 1713453518
transform 1 0 2456 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_176
timestamp 1713453518
transform 1 0 1680 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_177
timestamp 1713453518
transform 1 0 1416 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_178
timestamp 1713453518
transform 1 0 3272 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_179
timestamp 1713453518
transform 1 0 3208 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_180
timestamp 1713453518
transform 1 0 3080 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_181
timestamp 1713453518
transform 1 0 2752 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_182
timestamp 1713453518
transform 1 0 2264 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_183
timestamp 1713453518
transform 1 0 2384 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_184
timestamp 1713453518
transform 1 0 1656 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_185
timestamp 1713453518
transform 1 0 1368 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_186
timestamp 1713453518
transform 1 0 3136 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_187
timestamp 1713453518
transform 1 0 2912 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_188
timestamp 1713453518
transform 1 0 3040 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_189
timestamp 1713453518
transform 1 0 2872 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_190
timestamp 1713453518
transform 1 0 3384 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_191
timestamp 1713453518
transform 1 0 1824 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_192
timestamp 1713453518
transform 1 0 2256 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_193
timestamp 1713453518
transform 1 0 3024 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_194
timestamp 1713453518
transform 1 0 1696 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_195
timestamp 1713453518
transform 1 0 2800 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_196
timestamp 1713453518
transform 1 0 2856 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_197
timestamp 1713453518
transform 1 0 1200 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_198
timestamp 1713453518
transform 1 0 2568 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_199
timestamp 1713453518
transform 1 0 3400 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_200
timestamp 1713453518
transform 1 0 2160 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_201
timestamp 1713453518
transform 1 0 2256 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_202
timestamp 1713453518
transform 1 0 1096 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_203
timestamp 1713453518
transform 1 0 1672 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_204
timestamp 1713453518
transform 1 0 2704 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_205
timestamp 1713453518
transform 1 0 1720 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_206
timestamp 1713453518
transform 1 0 2776 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_207
timestamp 1713453518
transform 1 0 2768 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_208
timestamp 1713453518
transform 1 0 1752 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_209
timestamp 1713453518
transform 1 0 1304 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_210
timestamp 1713453518
transform 1 0 2744 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_211
timestamp 1713453518
transform 1 0 2192 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_212
timestamp 1713453518
transform 1 0 2360 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_213
timestamp 1713453518
transform 1 0 1648 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_214
timestamp 1713453518
transform 1 0 2680 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_215
timestamp 1713453518
transform 1 0 1720 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_216
timestamp 1713453518
transform 1 0 2760 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_217
timestamp 1713453518
transform 1 0 2736 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_218
timestamp 1713453518
transform 1 0 1744 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_219
timestamp 1713453518
transform 1 0 1208 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_220
timestamp 1713453518
transform 1 0 2768 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_221
timestamp 1713453518
transform 1 0 3368 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_222
timestamp 1713453518
transform 1 0 2280 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_223
timestamp 1713453518
transform 1 0 2304 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_224
timestamp 1713453518
transform 1 0 1632 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_225
timestamp 1713453518
transform 1 0 2752 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_226
timestamp 1713453518
transform 1 0 1680 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_227
timestamp 1713453518
transform 1 0 2928 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_228
timestamp 1713453518
transform 1 0 2864 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_229
timestamp 1713453518
transform 1 0 1744 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_230
timestamp 1713453518
transform 1 0 1344 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_231
timestamp 1713453518
transform 1 0 2560 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_232
timestamp 1713453518
transform 1 0 3352 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_233
timestamp 1713453518
transform 1 0 1552 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_234
timestamp 1713453518
transform 1 0 1640 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_235
timestamp 1713453518
transform 1 0 2912 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_236
timestamp 1713453518
transform 1 0 3016 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_237
timestamp 1713453518
transform 1 0 2784 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_238
timestamp 1713453518
transform 1 0 2992 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_239
timestamp 1713453518
transform 1 0 1304 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_240
timestamp 1713453518
transform 1 0 1384 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_241
timestamp 1713453518
transform 1 0 2808 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_242
timestamp 1713453518
transform 1 0 2512 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_243
timestamp 1713453518
transform 1 0 1664 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_244
timestamp 1713453518
transform 1 0 2400 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_245
timestamp 1713453518
transform 1 0 2184 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_246
timestamp 1713453518
transform 1 0 3192 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_247
timestamp 1713453518
transform 1 0 1288 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_248
timestamp 1713453518
transform 1 0 2456 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_249
timestamp 1713453518
transform 1 0 1656 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_250
timestamp 1713453518
transform 1 0 2424 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_251
timestamp 1713453518
transform 1 0 2216 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_252
timestamp 1713453518
transform 1 0 1344 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_253
timestamp 1713453518
transform 1 0 3216 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_254
timestamp 1713453518
transform 1 0 2488 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_255
timestamp 1713453518
transform 1 0 1696 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_256
timestamp 1713453518
transform 1 0 2472 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_257
timestamp 1713453518
transform 1 0 1928 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_258
timestamp 1713453518
transform 1 0 3160 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_259
timestamp 1713453518
transform 1 0 1368 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_260
timestamp 1713453518
transform 1 0 3088 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_261
timestamp 1713453518
transform 1 0 2112 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_262
timestamp 1713453518
transform 1 0 2344 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_263
timestamp 1713453518
transform 1 0 3208 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_264
timestamp 1713453518
transform 1 0 2232 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_265
timestamp 1713453518
transform 1 0 1344 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_266
timestamp 1713453518
transform 1 0 1528 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_267
timestamp 1713453518
transform 1 0 1336 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_268
timestamp 1713453518
transform 1 0 2488 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_269
timestamp 1713453518
transform 1 0 2256 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_270
timestamp 1713453518
transform 1 0 2312 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_271
timestamp 1713453518
transform 1 0 3088 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_272
timestamp 1713453518
transform 1 0 1272 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_273
timestamp 1713453518
transform 1 0 1208 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_274
timestamp 1713453518
transform 1 0 1584 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_275
timestamp 1713453518
transform 1 0 2208 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_276
timestamp 1713453518
transform 1 0 3112 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_277
timestamp 1713453518
transform 1 0 3120 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_278
timestamp 1713453518
transform 1 0 880 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_279
timestamp 1713453518
transform 1 0 3352 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_280
timestamp 1713453518
transform 1 0 3248 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_281
timestamp 1713453518
transform 1 0 3360 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_282
timestamp 1713453518
transform 1 0 3128 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_283
timestamp 1713453518
transform 1 0 3408 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_284
timestamp 1713453518
transform 1 0 1600 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_285
timestamp 1713453518
transform 1 0 1496 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_286
timestamp 1713453518
transform 1 0 1968 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_287
timestamp 1713453518
transform 1 0 2000 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_288
timestamp 1713453518
transform 1 0 2048 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_289
timestamp 1713453518
transform 1 0 2152 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_290
timestamp 1713453518
transform 1 0 344 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_291
timestamp 1713453518
transform 1 0 544 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_292
timestamp 1713453518
transform 1 0 216 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_293
timestamp 1713453518
transform 1 0 520 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_294
timestamp 1713453518
transform 1 0 648 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_295
timestamp 1713453518
transform 1 0 600 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_296
timestamp 1713453518
transform 1 0 504 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_297
timestamp 1713453518
transform 1 0 632 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_298
timestamp 1713453518
transform 1 0 672 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_299
timestamp 1713453518
transform 1 0 464 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_300
timestamp 1713453518
transform 1 0 464 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_301
timestamp 1713453518
transform 1 0 808 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_302
timestamp 1713453518
transform 1 0 872 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_303
timestamp 1713453518
transform 1 0 1352 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_304
timestamp 1713453518
transform 1 0 1352 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_305
timestamp 1713453518
transform 1 0 1328 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_306
timestamp 1713453518
transform 1 0 960 0 -1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1713453518
transform 1 0 3016 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1713453518
transform 1 0 2048 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1713453518
transform 1 0 2648 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1713453518
transform 1 0 2728 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1713453518
transform 1 0 2704 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1713453518
transform 1 0 2272 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1713453518
transform 1 0 2408 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1713453518
transform 1 0 2504 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1713453518
transform 1 0 1936 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1713453518
transform 1 0 1984 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1713453518
transform 1 0 2112 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1713453518
transform 1 0 1904 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1713453518
transform 1 0 2960 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1713453518
transform 1 0 3408 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1713453518
transform 1 0 3008 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1713453518
transform 1 0 2952 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1713453518
transform 1 0 2936 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1713453518
transform 1 0 2912 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1713453518
transform 1 0 3400 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1713453518
transform 1 0 3056 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1713453518
transform 1 0 2760 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1713453518
transform 1 0 2536 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1713453518
transform 1 0 1776 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1713453518
transform 1 0 3200 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1713453518
transform 1 0 2952 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1713453518
transform 1 0 3192 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1713453518
transform 1 0 3184 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1713453518
transform 1 0 2904 0 -1 3370
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1713453518
transform 1 0 3080 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1713453518
transform 1 0 2688 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1713453518
transform 1 0 2336 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1713453518
transform 1 0 1448 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1713453518
transform 1 0 3032 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1713453518
transform 1 0 2416 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1713453518
transform 1 0 3152 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1713453518
transform 1 0 1360 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1713453518
transform 1 0 2568 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1713453518
transform 1 0 3152 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1713453518
transform 1 0 1216 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1713453518
transform 1 0 2464 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1713453518
transform 1 0 2680 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1713453518
transform 1 0 1504 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1713453518
transform 1 0 2400 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1713453518
transform 1 0 2808 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1713453518
transform 1 0 2568 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1713453518
transform 1 0 2936 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1713453518
transform 1 0 1360 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1713453518
transform 1 0 2752 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_48
timestamp 1713453518
transform 1 0 3128 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_49
timestamp 1713453518
transform 1 0 2872 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_50
timestamp 1713453518
transform 1 0 3168 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_51
timestamp 1713453518
transform 1 0 2640 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_52
timestamp 1713453518
transform 1 0 2440 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_53
timestamp 1713453518
transform 1 0 1744 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_54
timestamp 1713453518
transform 1 0 2944 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1713453518
transform 1 0 2568 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_56
timestamp 1713453518
transform 1 0 2816 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_57
timestamp 1713453518
transform 1 0 1456 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_58
timestamp 1713453518
transform 1 0 2568 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_59
timestamp 1713453518
transform 1 0 3120 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_60
timestamp 1713453518
transform 1 0 1608 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_61
timestamp 1713453518
transform 1 0 2488 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_62
timestamp 1713453518
transform 1 0 3008 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_63
timestamp 1713453518
transform 1 0 1520 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_64
timestamp 1713453518
transform 1 0 2440 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_65
timestamp 1713453518
transform 1 0 2784 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_66
timestamp 1713453518
transform 1 0 2472 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_67
timestamp 1713453518
transform 1 0 2664 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_68
timestamp 1713453518
transform 1 0 1280 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_69
timestamp 1713453518
transform 1 0 1296 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_70
timestamp 1713453518
transform 1 0 2568 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_71
timestamp 1713453518
transform 1 0 3320 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_72
timestamp 1713453518
transform 1 0 2424 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_73
timestamp 1713453518
transform 1 0 3184 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_74
timestamp 1713453518
transform 1 0 2392 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_75
timestamp 1713453518
transform 1 0 2200 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_76
timestamp 1713453518
transform 1 0 1640 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_77
timestamp 1713453518
transform 1 0 2840 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_78
timestamp 1713453518
transform 1 0 2352 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_79
timestamp 1713453518
transform 1 0 2616 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_80
timestamp 1713453518
transform 1 0 1568 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_81
timestamp 1713453518
transform 1 0 2456 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_82
timestamp 1713453518
transform 1 0 2704 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_83
timestamp 1713453518
transform 1 0 1600 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_84
timestamp 1713453518
transform 1 0 2408 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_85
timestamp 1713453518
transform 1 0 2568 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_86
timestamp 1713453518
transform 1 0 1592 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_87
timestamp 1713453518
transform 1 0 2880 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_88
timestamp 1713453518
transform 1 0 2840 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_89
timestamp 1713453518
transform 1 0 1128 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_90
timestamp 1713453518
transform 1 0 1976 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_91
timestamp 1713453518
transform 1 0 1120 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_92
timestamp 1713453518
transform 1 0 2104 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_93
timestamp 1713453518
transform 1 0 3184 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_94
timestamp 1713453518
transform 1 0 1096 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_95
timestamp 1713453518
transform 1 0 1168 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_96
timestamp 1713453518
transform 1 0 3296 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_97
timestamp 1713453518
transform 1 0 1192 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_98
timestamp 1713453518
transform 1 0 1952 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_99
timestamp 1713453518
transform 1 0 3384 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_100
timestamp 1713453518
transform 1 0 1144 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_101
timestamp 1713453518
transform 1 0 1232 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_102
timestamp 1713453518
transform 1 0 3264 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_103
timestamp 1713453518
transform 1 0 1112 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_104
timestamp 1713453518
transform 1 0 2440 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_105
timestamp 1713453518
transform 1 0 3408 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_106
timestamp 1713453518
transform 1 0 1080 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_107
timestamp 1713453518
transform 1 0 3272 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_108
timestamp 1713453518
transform 1 0 1712 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_109
timestamp 1713453518
transform 1 0 1712 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_110
timestamp 1713453518
transform 1 0 1256 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_111
timestamp 1713453518
transform 1 0 1160 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_112
timestamp 1713453518
transform 1 0 1168 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_113
timestamp 1713453518
transform 1 0 3304 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_114
timestamp 1713453518
transform 1 0 3376 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_115
timestamp 1713453518
transform 1 0 2504 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_116
timestamp 1713453518
transform 1 0 3232 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_117
timestamp 1713453518
transform 1 0 2120 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_118
timestamp 1713453518
transform 1 0 2072 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_119
timestamp 1713453518
transform 1 0 2032 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_120
timestamp 1713453518
transform 1 0 1912 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_121
timestamp 1713453518
transform 1 0 1912 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_122
timestamp 1713453518
transform 1 0 2032 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_123
timestamp 1713453518
transform 1 0 1848 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_124
timestamp 1713453518
transform 1 0 576 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_125
timestamp 1713453518
transform 1 0 496 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_126
timestamp 1713453518
transform 1 0 496 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_127
timestamp 1713453518
transform 1 0 512 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_128
timestamp 1713453518
transform 1 0 528 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_129
timestamp 1713453518
transform 1 0 544 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_130
timestamp 1713453518
transform 1 0 480 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_131
timestamp 1713453518
transform 1 0 632 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_132
timestamp 1713453518
transform 1 0 440 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_133
timestamp 1713453518
transform 1 0 744 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_134
timestamp 1713453518
transform 1 0 664 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_135
timestamp 1713453518
transform 1 0 696 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_136
timestamp 1713453518
transform 1 0 696 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_137
timestamp 1713453518
transform 1 0 688 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_138
timestamp 1713453518
transform 1 0 760 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_139
timestamp 1713453518
transform 1 0 600 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_140
timestamp 1713453518
transform 1 0 544 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_141
timestamp 1713453518
transform 1 0 536 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_142
timestamp 1713453518
transform 1 0 568 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_143
timestamp 1713453518
transform 1 0 704 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_144
timestamp 1713453518
transform 1 0 808 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_145
timestamp 1713453518
transform 1 0 984 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_146
timestamp 1713453518
transform 1 0 728 0 1 370
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1713453518
transform 1 0 2944 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1713453518
transform 1 0 2488 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1713453518
transform 1 0 2704 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1713453518
transform 1 0 1920 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1713453518
transform 1 0 2640 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1713453518
transform 1 0 2760 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1713453518
transform 1 0 2392 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1713453518
transform 1 0 2104 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1713453518
transform 1 0 2224 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1713453518
transform 1 0 2288 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1713453518
transform 1 0 2016 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1713453518
transform 1 0 2064 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1713453518
transform 1 0 1920 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1713453518
transform 1 0 2016 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1713453518
transform 1 0 2056 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1713453518
transform 1 0 2072 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1713453518
transform 1 0 1896 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1713453518
transform 1 0 3400 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1713453518
transform 1 0 3400 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1713453518
transform 1 0 3424 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1713453518
transform 1 0 2944 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1713453518
transform 1 0 2528 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1713453518
transform 1 0 2920 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1713453518
transform 1 0 3416 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1713453518
transform 1 0 3328 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1713453518
transform 1 0 2704 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1713453518
transform 1 0 1992 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1713453518
transform 1 0 2576 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1713453518
transform 1 0 1680 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1713453518
transform 1 0 1872 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1713453518
transform 1 0 1720 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1713453518
transform 1 0 1872 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1713453518
transform 1 0 2216 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1713453518
transform 1 0 2200 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1713453518
transform 1 0 2960 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1713453518
transform 1 0 1344 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1713453518
transform 1 0 1232 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1713453518
transform 1 0 3000 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1713453518
transform 1 0 1248 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1713453518
transform 1 0 3024 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1713453518
transform 1 0 1144 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1713453518
transform 1 0 3056 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1713453518
transform 1 0 1208 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1713453518
transform 1 0 3032 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1713453518
transform 1 0 1400 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1713453518
transform 1 0 1480 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1713453518
transform 1 0 2464 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1713453518
transform 1 0 1256 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1713453518
transform 1 0 2392 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1713453518
transform 1 0 2768 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1713453518
transform 1 0 1120 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1713453518
transform 1 0 2248 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1713453518
transform 1 0 1872 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1713453518
transform 1 0 2608 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1713453518
transform 1 0 1112 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1713453518
transform 1 0 2288 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1713453518
transform 1 0 1824 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1713453518
transform 1 0 2648 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1713453518
transform 1 0 1560 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1713453518
transform 1 0 1992 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1713453518
transform 1 0 2816 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1713453518
transform 1 0 1464 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1713453518
transform 1 0 3072 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1713453518
transform 1 0 2024 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1713453518
transform 1 0 1656 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1713453518
transform 1 0 3064 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1713453518
transform 1 0 1688 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1713453518
transform 1 0 3040 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1713453518
transform 1 0 1344 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1713453518
transform 1 0 2408 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1713453518
transform 1 0 1920 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1713453518
transform 1 0 2784 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1713453518
transform 1 0 1248 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1713453518
transform 1 0 3160 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1713453518
transform 1 0 1456 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1713453518
transform 1 0 2824 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1713453518
transform 1 0 1440 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1713453518
transform 1 0 2664 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1713453518
transform 1 0 1472 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1713453518
transform 1 0 1472 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1713453518
transform 1 0 1128 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1713453518
transform 1 0 3096 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1713453518
transform 1 0 3328 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1713453518
transform 1 0 1552 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1713453518
transform 1 0 3320 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1713453518
transform 1 0 1576 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1713453518
transform 1 0 1600 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1713453518
transform 1 0 3144 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1713453518
transform 1 0 1440 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1713453518
transform 1 0 2096 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1713453518
transform 1 0 2696 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1713453518
transform 1 0 1368 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1713453518
transform 1 0 2072 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1713453518
transform 1 0 1144 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1713453518
transform 1 0 2624 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1713453518
transform 1 0 1320 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1713453518
transform 1 0 2048 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1713453518
transform 1 0 1096 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1713453518
transform 1 0 2592 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1713453518
transform 1 0 1272 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1713453518
transform 1 0 2008 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1713453518
transform 1 0 1072 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1713453518
transform 1 0 2712 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1713453518
transform 1 0 1112 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1713453518
transform 1 0 3160 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1713453518
transform 1 0 1248 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1713453518
transform 1 0 1120 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1713453518
transform 1 0 1472 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1713453518
transform 1 0 1096 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1713453518
transform 1 0 1272 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1713453518
transform 1 0 1232 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1713453518
transform 1 0 1200 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1713453518
transform 1 0 1128 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1713453518
transform 1 0 1224 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1713453518
transform 1 0 1232 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1713453518
transform 1 0 1048 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1713453518
transform 1 0 1064 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1713453518
transform 1 0 1208 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1713453518
transform 1 0 1216 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1713453518
transform 1 0 3184 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1713453518
transform 1 0 888 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1713453518
transform 1 0 3168 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1713453518
transform 1 0 3224 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1713453518
transform 1 0 2072 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1713453518
transform 1 0 360 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1713453518
transform 1 0 240 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_126
timestamp 1713453518
transform 1 0 416 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_127
timestamp 1713453518
transform 1 0 504 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_128
timestamp 1713453518
transform 1 0 528 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_129
timestamp 1713453518
transform 1 0 616 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_130
timestamp 1713453518
transform 1 0 616 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_131
timestamp 1713453518
transform 1 0 472 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_132
timestamp 1713453518
transform 1 0 496 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_133
timestamp 1713453518
transform 1 0 592 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_134
timestamp 1713453518
transform 1 0 680 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_135
timestamp 1713453518
transform 1 0 240 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_136
timestamp 1713453518
transform 1 0 224 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_137
timestamp 1713453518
transform 1 0 232 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_138
timestamp 1713453518
transform 1 0 296 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_139
timestamp 1713453518
transform 1 0 464 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_140
timestamp 1713453518
transform 1 0 656 0 -1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_141
timestamp 1713453518
transform 1 0 640 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_142
timestamp 1713453518
transform 1 0 256 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_143
timestamp 1713453518
transform 1 0 296 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_144
timestamp 1713453518
transform 1 0 304 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_145
timestamp 1713453518
transform 1 0 248 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_146
timestamp 1713453518
transform 1 0 184 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_147
timestamp 1713453518
transform 1 0 424 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_148
timestamp 1713453518
transform 1 0 256 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_149
timestamp 1713453518
transform 1 0 264 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_150
timestamp 1713453518
transform 1 0 264 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_151
timestamp 1713453518
transform 1 0 256 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_152
timestamp 1713453518
transform 1 0 144 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_153
timestamp 1713453518
transform 1 0 304 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_154
timestamp 1713453518
transform 1 0 472 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_155
timestamp 1713453518
transform 1 0 192 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_156
timestamp 1713453518
transform 1 0 240 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_157
timestamp 1713453518
transform 1 0 264 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_158
timestamp 1713453518
transform 1 0 240 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_159
timestamp 1713453518
transform 1 0 224 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_160
timestamp 1713453518
transform 1 0 88 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_161
timestamp 1713453518
transform 1 0 216 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_162
timestamp 1713453518
transform 1 0 112 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_163
timestamp 1713453518
transform 1 0 432 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_164
timestamp 1713453518
transform 1 0 376 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_165
timestamp 1713453518
transform 1 0 288 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_166
timestamp 1713453518
transform 1 0 576 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_167
timestamp 1713453518
transform 1 0 664 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_168
timestamp 1713453518
transform 1 0 680 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_169
timestamp 1713453518
transform 1 0 760 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_170
timestamp 1713453518
transform 1 0 520 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_171
timestamp 1713453518
transform 1 0 696 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_172
timestamp 1713453518
transform 1 0 720 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_173
timestamp 1713453518
transform 1 0 632 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_174
timestamp 1713453518
transform 1 0 1232 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_175
timestamp 1713453518
transform 1 0 848 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_176
timestamp 1713453518
transform 1 0 480 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_177
timestamp 1713453518
transform 1 0 640 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_178
timestamp 1713453518
transform 1 0 1712 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_179
timestamp 1713453518
transform 1 0 1808 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_180
timestamp 1713453518
transform 1 0 328 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_181
timestamp 1713453518
transform 1 0 1784 0 -1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_0
timestamp 1713453518
transform 1 0 2712 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1713453518
transform 1 0 1984 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1713453518
transform 1 0 2664 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1713453518
transform 1 0 2856 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1713453518
transform 1 0 1920 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1713453518
transform 1 0 2200 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1713453518
transform 1 0 2352 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1713453518
transform 1 0 1968 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1713453518
transform 1 0 2016 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1713453518
transform 1 0 1984 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1713453518
transform 1 0 2016 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1713453518
transform 1 0 1888 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1713453518
transform 1 0 1512 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1713453518
transform 1 0 2056 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1713453518
transform 1 0 1864 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1713453518
transform 1 0 3376 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1713453518
transform 1 0 3176 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1713453518
transform 1 0 3144 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1713453518
transform 1 0 3368 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1713453518
transform 1 0 3392 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1713453518
transform 1 0 2496 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1713453518
transform 1 0 2888 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1713453518
transform 1 0 2920 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1713453518
transform 1 0 3064 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1713453518
transform 1 0 3384 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1713453518
transform 1 0 3392 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1713453518
transform 1 0 2136 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1713453518
transform 1 0 3408 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1713453518
transform 1 0 3272 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1713453518
transform 1 0 2752 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1713453518
transform 1 0 2664 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1713453518
transform 1 0 1976 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1713453518
transform 1 0 2648 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1713453518
transform 1 0 2544 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1713453518
transform 1 0 888 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1713453518
transform 1 0 1504 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1713453518
transform 1 0 1568 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1713453518
transform 1 0 1024 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1713453518
transform 1 0 1296 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1713453518
transform 1 0 1768 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1713453518
transform 1 0 1312 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1713453518
transform 1 0 864 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1713453518
transform 1 0 1480 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1713453518
transform 1 0 1440 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1713453518
transform 1 0 1136 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1713453518
transform 1 0 1360 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1713453518
transform 1 0 1800 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1713453518
transform 1 0 1344 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1713453518
transform 1 0 880 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1713453518
transform 1 0 1448 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1713453518
transform 1 0 1432 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1713453518
transform 1 0 1176 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1713453518
transform 1 0 1984 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1713453518
transform 1 0 1376 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1713453518
transform 1 0 1040 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1713453518
transform 1 0 1816 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1713453518
transform 1 0 1512 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1713453518
transform 1 0 1424 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1713453518
transform 1 0 1248 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1713453518
transform 1 0 2752 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1713453518
transform 1 0 1312 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1713453518
transform 1 0 1184 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1713453518
transform 1 0 1240 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1713453518
transform 1 0 1072 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1713453518
transform 1 0 2512 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1713453518
transform 1 0 1072 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1713453518
transform 1 0 3080 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1713453518
transform 1 0 2192 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1713453518
transform 1 0 1280 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1713453518
transform 1 0 1256 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1713453518
transform 1 0 1120 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1713453518
transform 1 0 2536 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1713453518
transform 1 0 1160 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1713453518
transform 1 0 1008 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1713453518
transform 1 0 3224 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1713453518
transform 1 0 2608 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1713453518
transform 1 0 2680 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1713453518
transform 1 0 1096 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1713453518
transform 1 0 2488 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1713453518
transform 1 0 1264 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1713453518
transform 1 0 1112 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1713453518
transform 1 0 3096 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1713453518
transform 1 0 2768 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1713453518
transform 1 0 2832 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1713453518
transform 1 0 1040 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1713453518
transform 1 0 2536 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1713453518
transform 1 0 3112 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1713453518
transform 1 0 1464 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1713453518
transform 1 0 1064 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1713453518
transform 1 0 1888 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1713453518
transform 1 0 1584 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1713453518
transform 1 0 1056 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1713453518
transform 1 0 3064 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1713453518
transform 1 0 1352 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1713453518
transform 1 0 1024 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1713453518
transform 1 0 1808 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1713453518
transform 1 0 1632 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1713453518
transform 1 0 1048 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1713453518
transform 1 0 3096 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1713453518
transform 1 0 1280 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1713453518
transform 1 0 1016 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1713453518
transform 1 0 1992 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1713453518
transform 1 0 1784 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1713453518
transform 1 0 1096 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1713453518
transform 1 0 2768 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1713453518
transform 1 0 1568 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1713453518
transform 1 0 1064 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1713453518
transform 1 0 2168 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1713453518
transform 1 0 1696 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1713453518
transform 1 0 1072 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1713453518
transform 1 0 2672 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1713453518
transform 1 0 1304 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1713453518
transform 1 0 1176 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1713453518
transform 1 0 1040 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1713453518
transform 1 0 2064 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1713453518
transform 1 0 1632 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1713453518
transform 1 0 1088 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1713453518
transform 1 0 2872 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1713453518
transform 1 0 2224 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1713453518
transform 1 0 1432 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1713453518
transform 1 0 1400 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1713453518
transform 1 0 984 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1713453518
transform 1 0 1784 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1713453518
transform 1 0 1712 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1713453518
transform 1 0 1016 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1713453518
transform 1 0 3056 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1713453518
transform 1 0 2632 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1713453518
transform 1 0 2760 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1713453518
transform 1 0 1000 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1713453518
transform 1 0 2472 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1713453518
transform 1 0 1768 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1713453518
transform 1 0 1080 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1713453518
transform 1 0 3112 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1713453518
transform 1 0 2736 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1713453518
transform 1 0 2808 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1713453518
transform 1 0 1024 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1713453518
transform 1 0 2392 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1713453518
transform 1 0 3088 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1713453518
transform 1 0 1392 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1713453518
transform 1 0 1056 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1713453518
transform 1 0 2320 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1713453518
transform 1 0 1832 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1713453518
transform 1 0 1088 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1713453518
transform 1 0 2872 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1713453518
transform 1 0 1528 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1713453518
transform 1 0 1064 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1713453518
transform 1 0 2344 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1713453518
transform 1 0 1832 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1713453518
transform 1 0 1152 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1713453518
transform 1 0 3176 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1713453518
transform 1 0 1632 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1713453518
transform 1 0 1000 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1713453518
transform 1 0 2312 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1713453518
transform 1 0 1800 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1713453518
transform 1 0 1080 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1713453518
transform 1 0 2880 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1713453518
transform 1 0 1520 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1713453518
transform 1 0 1024 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1713453518
transform 1 0 1880 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1713453518
transform 1 0 1776 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1713453518
transform 1 0 1064 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1713453518
transform 1 0 2696 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1713453518
transform 1 0 1248 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_163
timestamp 1713453518
transform 1 0 1216 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_164
timestamp 1713453518
transform 1 0 984 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_165
timestamp 1713453518
transform 1 0 1816 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_166
timestamp 1713453518
transform 1 0 1752 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_167
timestamp 1713453518
transform 1 0 1056 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_168
timestamp 1713453518
transform 1 0 2656 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_169
timestamp 1713453518
transform 1 0 2160 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_170
timestamp 1713453518
transform 1 0 1432 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_171
timestamp 1713453518
transform 1 0 1360 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_172
timestamp 1713453518
transform 1 0 1216 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_173
timestamp 1713453518
transform 1 0 1056 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_174
timestamp 1713453518
transform 1 0 2016 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_175
timestamp 1713453518
transform 1 0 1752 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_176
timestamp 1713453518
transform 1 0 1016 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_177
timestamp 1713453518
transform 1 0 3384 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_178
timestamp 1713453518
transform 1 0 2504 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_179
timestamp 1713453518
transform 1 0 2568 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_180
timestamp 1713453518
transform 1 0 1216 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_181
timestamp 1713453518
transform 1 0 960 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_182
timestamp 1713453518
transform 1 0 2232 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_183
timestamp 1713453518
transform 1 0 1728 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_184
timestamp 1713453518
transform 1 0 1032 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_185
timestamp 1713453518
transform 1 0 3304 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_186
timestamp 1713453518
transform 1 0 2512 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_187
timestamp 1713453518
transform 1 0 2448 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_188
timestamp 1713453518
transform 1 0 1232 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_189
timestamp 1713453518
transform 1 0 1064 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_190
timestamp 1713453518
transform 1 0 1768 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_191
timestamp 1713453518
transform 1 0 3184 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_192
timestamp 1713453518
transform 1 0 1432 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_193
timestamp 1713453518
transform 1 0 992 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_194
timestamp 1713453518
transform 1 0 2184 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_195
timestamp 1713453518
transform 1 0 1960 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_196
timestamp 1713453518
transform 1 0 1056 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_197
timestamp 1713453518
transform 1 0 2720 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_198
timestamp 1713453518
transform 1 0 1560 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_199
timestamp 1713453518
transform 1 0 1016 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_200
timestamp 1713453518
transform 1 0 2176 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_201
timestamp 1713453518
transform 1 0 1792 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_202
timestamp 1713453518
transform 1 0 1088 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_203
timestamp 1713453518
transform 1 0 2648 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_204
timestamp 1713453518
transform 1 0 1632 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_205
timestamp 1713453518
transform 1 0 1008 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_206
timestamp 1713453518
transform 1 0 2280 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_207
timestamp 1713453518
transform 1 0 1816 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_208
timestamp 1713453518
transform 1 0 1024 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_209
timestamp 1713453518
transform 1 0 2632 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_210
timestamp 1713453518
transform 1 0 1624 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_211
timestamp 1713453518
transform 1 0 960 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_212
timestamp 1713453518
transform 1 0 1800 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_213
timestamp 1713453518
transform 1 0 1976 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_214
timestamp 1713453518
transform 1 0 1712 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_215
timestamp 1713453518
transform 1 0 1264 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_216
timestamp 1713453518
transform 1 0 1496 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_217
timestamp 1713453518
transform 1 0 1408 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_218
timestamp 1713453518
transform 1 0 1024 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_219
timestamp 1713453518
transform 1 0 1840 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_220
timestamp 1713453518
transform 1 0 1912 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_221
timestamp 1713453518
transform 1 0 1872 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_222
timestamp 1713453518
transform 1 0 1056 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_223
timestamp 1713453518
transform 1 0 2040 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_224
timestamp 1713453518
transform 1 0 2008 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_225
timestamp 1713453518
transform 1 0 1384 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_226
timestamp 1713453518
transform 1 0 1808 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_227
timestamp 1713453518
transform 1 0 1760 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_228
timestamp 1713453518
transform 1 0 1056 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_229
timestamp 1713453518
transform 1 0 1904 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_230
timestamp 1713453518
transform 1 0 2104 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_231
timestamp 1713453518
transform 1 0 1704 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_232
timestamp 1713453518
transform 1 0 1000 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_233
timestamp 1713453518
transform 1 0 2136 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_234
timestamp 1713453518
transform 1 0 2056 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_235
timestamp 1713453518
transform 1 0 1416 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_236
timestamp 1713453518
transform 1 0 1920 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_237
timestamp 1713453518
transform 1 0 1688 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_238
timestamp 1713453518
transform 1 0 1008 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_239
timestamp 1713453518
transform 1 0 1832 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_240
timestamp 1713453518
transform 1 0 1944 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_241
timestamp 1713453518
transform 1 0 1800 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_242
timestamp 1713453518
transform 1 0 992 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_243
timestamp 1713453518
transform 1 0 2120 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_244
timestamp 1713453518
transform 1 0 2024 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_245
timestamp 1713453518
transform 1 0 1296 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_246
timestamp 1713453518
transform 1 0 1840 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_247
timestamp 1713453518
transform 1 0 1760 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_248
timestamp 1713453518
transform 1 0 848 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_249
timestamp 1713453518
transform 1 0 2056 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_250
timestamp 1713453518
transform 1 0 2208 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_251
timestamp 1713453518
transform 1 0 2208 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_252
timestamp 1713453518
transform 1 0 1520 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_253
timestamp 1713453518
transform 1 0 2024 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_254
timestamp 1713453518
transform 1 0 1712 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_255
timestamp 1713453518
transform 1 0 2752 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_256
timestamp 1713453518
transform 1 0 2792 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_257
timestamp 1713453518
transform 1 0 2896 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_258
timestamp 1713453518
transform 1 0 2824 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_259
timestamp 1713453518
transform 1 0 3320 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_260
timestamp 1713453518
transform 1 0 3216 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_261
timestamp 1713453518
transform 1 0 3384 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_262
timestamp 1713453518
transform 1 0 3152 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_263
timestamp 1713453518
transform 1 0 3360 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_264
timestamp 1713453518
transform 1 0 2352 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_265
timestamp 1713453518
transform 1 0 2120 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_266
timestamp 1713453518
transform 1 0 3112 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_267
timestamp 1713453518
transform 1 0 2976 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_268
timestamp 1713453518
transform 1 0 2736 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_269
timestamp 1713453518
transform 1 0 2664 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_270
timestamp 1713453518
transform 1 0 3104 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_271
timestamp 1713453518
transform 1 0 2000 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_272
timestamp 1713453518
transform 1 0 1944 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_273
timestamp 1713453518
transform 1 0 296 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_274
timestamp 1713453518
transform 1 0 472 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_275
timestamp 1713453518
transform 1 0 136 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_276
timestamp 1713453518
transform 1 0 560 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_277
timestamp 1713453518
transform 1 0 528 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_278
timestamp 1713453518
transform 1 0 248 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_279
timestamp 1713453518
transform 1 0 464 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_280
timestamp 1713453518
transform 1 0 560 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_281
timestamp 1713453518
transform 1 0 208 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_282
timestamp 1713453518
transform 1 0 640 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_283
timestamp 1713453518
transform 1 0 232 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_284
timestamp 1713453518
transform 1 0 608 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_285
timestamp 1713453518
transform 1 0 208 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_286
timestamp 1713453518
transform 1 0 552 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_287
timestamp 1713453518
transform 1 0 144 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_288
timestamp 1713453518
transform 1 0 648 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_289
timestamp 1713453518
transform 1 0 552 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_290
timestamp 1713453518
transform 1 0 600 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_291
timestamp 1713453518
transform 1 0 344 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_292
timestamp 1713453518
transform 1 0 576 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_293
timestamp 1713453518
transform 1 0 328 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_294
timestamp 1713453518
transform 1 0 712 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_295
timestamp 1713453518
transform 1 0 224 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_296
timestamp 1713453518
transform 1 0 616 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_297
timestamp 1713453518
transform 1 0 224 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_298
timestamp 1713453518
transform 1 0 664 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_299
timestamp 1713453518
transform 1 0 232 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_300
timestamp 1713453518
transform 1 0 568 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_301
timestamp 1713453518
transform 1 0 232 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_302
timestamp 1713453518
transform 1 0 664 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_303
timestamp 1713453518
transform 1 0 224 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_304
timestamp 1713453518
transform 1 0 720 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_305
timestamp 1713453518
transform 1 0 392 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_306
timestamp 1713453518
transform 1 0 688 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_307
timestamp 1713453518
transform 1 0 560 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_308
timestamp 1713453518
transform 1 0 608 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_309
timestamp 1713453518
transform 1 0 200 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_310
timestamp 1713453518
transform 1 0 576 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_311
timestamp 1713453518
transform 1 0 216 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_312
timestamp 1713453518
transform 1 0 632 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_313
timestamp 1713453518
transform 1 0 272 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_314
timestamp 1713453518
transform 1 0 736 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_315
timestamp 1713453518
transform 1 0 264 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_316
timestamp 1713453518
transform 1 0 712 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_317
timestamp 1713453518
transform 1 0 640 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_318
timestamp 1713453518
transform 1 0 568 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_319
timestamp 1713453518
transform 1 0 224 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_320
timestamp 1713453518
transform 1 0 688 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_321
timestamp 1713453518
transform 1 0 592 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_322
timestamp 1713453518
transform 1 0 776 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_323
timestamp 1713453518
transform 1 0 624 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_324
timestamp 1713453518
transform 1 0 800 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_325
timestamp 1713453518
transform 1 0 440 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_326
timestamp 1713453518
transform 1 0 832 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_327
timestamp 1713453518
transform 1 0 248 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_328
timestamp 1713453518
transform 1 0 528 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_329
timestamp 1713453518
transform 1 0 200 0 -1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_330
timestamp 1713453518
transform 1 0 616 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_331
timestamp 1713453518
transform 1 0 192 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_332
timestamp 1713453518
transform 1 0 576 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_333
timestamp 1713453518
transform 1 0 208 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_334
timestamp 1713453518
transform 1 0 560 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_335
timestamp 1713453518
transform 1 0 536 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_336
timestamp 1713453518
transform 1 0 448 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_337
timestamp 1713453518
transform 1 0 440 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_338
timestamp 1713453518
transform 1 0 480 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_339
timestamp 1713453518
transform 1 0 448 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_340
timestamp 1713453518
transform 1 0 504 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_341
timestamp 1713453518
transform 1 0 648 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_342
timestamp 1713453518
transform 1 0 640 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_343
timestamp 1713453518
transform 1 0 568 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_344
timestamp 1713453518
transform 1 0 1232 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_345
timestamp 1713453518
transform 1 0 1264 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_346
timestamp 1713453518
transform 1 0 736 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_347
timestamp 1713453518
transform 1 0 1464 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_348
timestamp 1713453518
transform 1 0 1384 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_349
timestamp 1713453518
transform 1 0 1288 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_350
timestamp 1713453518
transform 1 0 1680 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_351
timestamp 1713453518
transform 1 0 1512 0 -1 170
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1713453518
transform 1 0 1664 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1713453518
transform 1 0 2936 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1713453518
transform 1 0 2400 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1713453518
transform 1 0 1760 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1713453518
transform 1 0 2136 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1713453518
transform 1 0 1944 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1713453518
transform 1 0 2048 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1713453518
transform 1 0 1872 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1713453518
transform 1 0 1608 0 1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1713453518
transform 1 0 1608 0 -1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1713453518
transform 1 0 2080 0 -1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1713453518
transform 1 0 1416 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1713453518
transform 1 0 1296 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1713453518
transform 1 0 1344 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1713453518
transform 1 0 1168 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1713453518
transform 1 0 1400 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1713453518
transform 1 0 1160 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1713453518
transform 1 0 1616 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1713453518
transform 1 0 1432 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1713453518
transform 1 0 1600 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1713453518
transform 1 0 1656 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1713453518
transform 1 0 1304 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1713453518
transform 1 0 1592 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1713453518
transform 1 0 1456 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1713453518
transform 1 0 1560 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1713453518
transform 1 0 1488 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1713453518
transform 1 0 1576 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1713453518
transform 1 0 1400 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1713453518
transform 1 0 1544 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1713453518
transform 1 0 1384 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1713453518
transform 1 0 1368 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1713453518
transform 1 0 1192 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1713453518
transform 1 0 1288 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1713453518
transform 1 0 1144 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1713453518
transform 1 0 1656 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1713453518
transform 1 0 1352 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_36
timestamp 1713453518
transform 1 0 1496 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_37
timestamp 1713453518
transform 1 0 1432 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_38
timestamp 1713453518
transform 1 0 1496 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1713453518
transform 1 0 1440 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_40
timestamp 1713453518
transform 1 0 1616 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_41
timestamp 1713453518
transform 1 0 1488 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1713453518
transform 1 0 1760 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_43
timestamp 1713453518
transform 1 0 1464 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_44
timestamp 1713453518
transform 1 0 2256 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_45
timestamp 1713453518
transform 1 0 1328 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_46
timestamp 1713453518
transform 1 0 1432 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_47
timestamp 1713453518
transform 1 0 2320 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_48
timestamp 1713453518
transform 1 0 1352 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_49
timestamp 1713453518
transform 1 0 1440 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_50
timestamp 1713453518
transform 1 0 2376 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_51
timestamp 1713453518
transform 1 0 1320 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_52
timestamp 1713453518
transform 1 0 2312 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_53
timestamp 1713453518
transform 1 0 1800 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_54
timestamp 1713453518
transform 1 0 2424 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_55
timestamp 1713453518
transform 1 0 2248 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_56
timestamp 1713453518
transform 1 0 2928 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_57
timestamp 1713453518
transform 1 0 2848 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_58
timestamp 1713453518
transform 1 0 2752 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_59
timestamp 1713453518
transform 1 0 2216 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_60
timestamp 1713453518
transform 1 0 2152 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_61
timestamp 1713453518
transform 1 0 1936 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_62
timestamp 1713453518
transform 1 0 1864 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_63
timestamp 1713453518
transform 1 0 328 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_64
timestamp 1713453518
transform 1 0 432 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_65
timestamp 1713453518
transform 1 0 104 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_66
timestamp 1713453518
transform 1 0 208 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_67
timestamp 1713453518
transform 1 0 496 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_68
timestamp 1713453518
transform 1 0 784 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_69
timestamp 1713453518
transform 1 0 1504 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_70
timestamp 1713453518
transform 1 0 1392 0 1 170
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1713453518
transform 1 0 1376 0 1 370
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1713453518
transform 1 0 496 0 1 370
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1713453518
transform 1 0 2616 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1713453518
transform 1 0 2432 0 1 570
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1713453518
transform 1 0 2648 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1713453518
transform 1 0 3368 0 1 1370
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1713453518
transform 1 0 1512 0 1 3170
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1713453518
transform 1 0 1544 0 -1 3370
box -8 -3 40 105
use OR2X1  OR2X1_8
timestamp 1713453518
transform 1 0 1928 0 -1 3370
box -8 -3 40 105
use OR2X1  OR2X1_9
timestamp 1713453518
transform 1 0 1944 0 1 3170
box -8 -3 40 105
use OR2X1  OR2X1_10
timestamp 1713453518
transform 1 0 2848 0 1 2770
box -8 -3 40 105
use OR2X1  OR2X1_11
timestamp 1713453518
transform 1 0 2872 0 1 2970
box -8 -3 40 105
use OR2X1  OR2X1_12
timestamp 1713453518
transform 1 0 3192 0 -1 3170
box -8 -3 40 105
use OR2X1  OR2X1_13
timestamp 1713453518
transform 1 0 1656 0 1 2570
box -8 -3 40 105
use OR2X1  OR2X1_14
timestamp 1713453518
transform 1 0 1752 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_15
timestamp 1713453518
transform 1 0 2368 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_16
timestamp 1713453518
transform 1 0 1920 0 1 1770
box -8 -3 40 105
use OR2X1  OR2X1_17
timestamp 1713453518
transform 1 0 2224 0 -1 1770
box -8 -3 40 105
use OR2X1  OR2X1_18
timestamp 1713453518
transform 1 0 2048 0 1 1570
box -8 -3 40 105
use OR2X1  OR2X1_19
timestamp 1713453518
transform 1 0 1808 0 -1 1570
box -8 -3 40 105
use OR2X1  OR2X1_20
timestamp 1713453518
transform 1 0 2096 0 1 1370
box -8 -3 40 105
use OR2X1  OR2X1_21
timestamp 1713453518
transform 1 0 2168 0 -1 1370
box -8 -3 40 105
use OR2X1  OR2X1_22
timestamp 1713453518
transform 1 0 1768 0 1 970
box -8 -3 40 105
use OR2X1  OR2X1_23
timestamp 1713453518
transform 1 0 1248 0 -1 970
box -8 -3 40 105
use OR2X1  OR2X1_24
timestamp 1713453518
transform 1 0 1976 0 -1 370
box -8 -3 40 105
use OR2X1  OR2X1_25
timestamp 1713453518
transform 1 0 2312 0 1 170
box -8 -3 40 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1713453518
transform 1 0 3496 0 1 3417
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1713453518
transform 1 0 3496 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1713453518
transform 1 0 24 0 1 3417
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1713453518
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1713453518
transform 1 0 3472 0 1 3393
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1713453518
transform 1 0 3472 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1713453518
transform 1 0 48 0 1 3393
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1713453518
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1713453518
transform 1 0 3496 0 1 3270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1713453518
transform 1 0 3496 0 1 3070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1713453518
transform 1 0 3496 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1713453518
transform 1 0 3496 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1713453518
transform 1 0 3496 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1713453518
transform 1 0 3496 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1713453518
transform 1 0 3496 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1713453518
transform 1 0 3496 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1713453518
transform 1 0 3496 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1713453518
transform 1 0 3496 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1713453518
transform 1 0 3496 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1713453518
transform 1 0 3496 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1713453518
transform 1 0 3496 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1713453518
transform 1 0 3496 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1713453518
transform 1 0 3496 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1713453518
transform 1 0 3496 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1713453518
transform 1 0 3496 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1713453518
transform 1 0 24 0 1 3270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1713453518
transform 1 0 24 0 1 3070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1713453518
transform 1 0 24 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1713453518
transform 1 0 24 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1713453518
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1713453518
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1713453518
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1713453518
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1713453518
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1713453518
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1713453518
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1713453518
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1713453518
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1713453518
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1713453518
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1713453518
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1713453518
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1713453518
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1713453518
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1713453518
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1713453518
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1713453518
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1713453518
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1713453518
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1713453518
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1713453518
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1713453518
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1713453518
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1713453518
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1713453518
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1713453518
transform 1 0 48 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1713453518
transform 1 0 48 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1713453518
transform 1 0 48 0 1 3170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_50
timestamp 1713453518
transform 1 0 48 0 1 3370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_51
timestamp 1713453518
transform 1 0 3472 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_52
timestamp 1713453518
transform 1 0 3472 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_53
timestamp 1713453518
transform 1 0 3472 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_54
timestamp 1713453518
transform 1 0 3472 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_55
timestamp 1713453518
transform 1 0 3472 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_56
timestamp 1713453518
transform 1 0 3472 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_57
timestamp 1713453518
transform 1 0 3472 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_58
timestamp 1713453518
transform 1 0 3472 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_59
timestamp 1713453518
transform 1 0 3472 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_60
timestamp 1713453518
transform 1 0 3472 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_61
timestamp 1713453518
transform 1 0 3472 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_62
timestamp 1713453518
transform 1 0 3472 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_63
timestamp 1713453518
transform 1 0 3472 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_64
timestamp 1713453518
transform 1 0 3472 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_65
timestamp 1713453518
transform 1 0 3472 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_66
timestamp 1713453518
transform 1 0 3472 0 1 3170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_67
timestamp 1713453518
transform 1 0 3472 0 1 3370
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1713453518
transform 1 0 2800 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1713453518
transform 1 0 2944 0 -1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1713453518
transform 1 0 2880 0 -1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1713453518
transform 1 0 3352 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_3
timestamp 1713453518
transform 1 0 3392 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1713453518
transform 1 0 2304 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_5
timestamp 1713453518
transform 1 0 2448 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_6
timestamp 1713453518
transform 1 0 2592 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_7
timestamp 1713453518
transform 1 0 3192 0 1 170
box -8 -3 64 105
use XOR2X1  XOR2X1_8
timestamp 1713453518
transform 1 0 3168 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_9
timestamp 1713453518
transform 1 0 3264 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_10
timestamp 1713453518
transform 1 0 3280 0 -1 370
box -8 -3 64 105
<< labels >>
rlabel metal2 684 1 684 1 4 in_clka
rlabel metal3 2 945 2 945 4 in_clkb
rlabel metal2 1108 1 1108 1 4 in_restart
rlabel metal2 1788 1 1788 1 4 in_move[1]
rlabel metal2 1732 1 1732 1 4 in_move[0]
rlabel metal2 836 3438 836 3438 4 board_out[31]
rlabel metal2 852 3438 852 3438 4 board_out[30]
rlabel metal2 964 3438 964 3438 4 board_out[29]
rlabel metal3 2 2925 2 2925 4 board_out[28]
rlabel metal2 764 3438 764 3438 4 board_out[27]
rlabel metal2 812 3438 812 3438 4 board_out[26]
rlabel metal2 868 3438 868 3438 4 board_out[25]
rlabel metal3 2 2765 2 2765 4 board_out[24]
rlabel metal3 2 2615 2 2615 4 board_out[23]
rlabel metal3 2 2555 2 2555 4 board_out[22]
rlabel metal3 2 2495 2 2495 4 board_out[21]
rlabel metal3 2 2415 2 2415 4 board_out[20]
rlabel metal3 2 2345 2 2345 4 board_out[19]
rlabel metal3 2 2315 2 2315 4 board_out[18]
rlabel metal3 2 2155 2 2155 4 board_out[17]
rlabel metal3 2 2295 2 2295 4 board_out[16]
rlabel metal3 2 1995 2 1995 4 board_out[15]
rlabel metal3 2 1905 2 1905 4 board_out[14]
rlabel metal3 2 1845 2 1845 4 board_out[13]
rlabel metal3 2 1825 2 1825 4 board_out[12]
rlabel metal3 2 1635 2 1635 4 board_out[11]
rlabel metal3 2 1515 2 1515 4 board_out[10]
rlabel metal3 2 1485 2 1485 4 board_out[9]
rlabel metal3 2 1585 2 1585 4 board_out[8]
rlabel metal3 2 1095 2 1095 4 board_out[7]
rlabel metal3 2 1075 2 1075 4 board_out[6]
rlabel metal3 2 1045 2 1045 4 board_out[5]
rlabel metal3 2 1025 2 1025 4 board_out[4]
rlabel metal3 2 1005 2 1005 4 board_out[3]
rlabel metal3 2 985 2 985 4 board_out[2]
rlabel metal3 2 965 2 965 4 board_out[1]
rlabel metal3 2 925 2 925 4 board_out[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 22932.000 855.000 22932.000 1125.000 
<< end >>
