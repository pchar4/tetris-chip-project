magic
tech scmos
timestamp 1711653199
<< end >>
