magic
tech scmos
timestamp 1712698519
<< metal1 >>
rect -1370 4098 -1331 4120
rect -1063 4099 -1035 4117
rect -765 4101 -734 4125
rect -462 4097 -431 4116
rect -164 4096 -128 4116
rect 129 4094 174 4116
rect 734 4098 766 4115
rect 1034 4100 1069 4114
rect 1341 4094 1368 4117
rect 1633 4094 1671 4121
rect 1929 4094 1965 4115
rect 2233 4093 2272 4114
rect 2828 4094 2871 4113
rect 3131 4097 3180 4118
rect -1389 3381 -1385 3388
rect -1477 3377 -1385 3381
rect -1089 3381 -1085 3388
rect -1177 3377 -1085 3381
rect -789 3381 -785 3388
rect -877 3377 -785 3381
rect -489 3381 -485 3388
rect -577 3377 -485 3381
rect -189 3381 -185 3388
rect -277 3377 -185 3381
rect 111 3375 115 3388
rect 23 3371 115 3375
rect 435 3355 458 3407
rect 711 3375 715 3388
rect 623 3371 715 3375
rect 1011 3375 1015 3388
rect 923 3371 1015 3375
rect 1311 3375 1315 3388
rect 1223 3371 1315 3375
rect 1611 3375 1615 3388
rect 1911 3381 1915 3394
rect 1823 3377 1915 3381
rect 1523 3371 1615 3375
rect 2211 3375 2215 3388
rect 2811 3381 2815 3392
rect 2723 3377 2815 3381
rect 3111 3381 3115 3388
rect 3023 3377 3115 3381
rect 2123 3371 2215 3375
rect 435 3332 630 3355
rect -2224 3235 -2193 3269
rect -1492 3211 -1477 3215
rect -1481 3123 -1477 3211
rect -2227 2945 -2190 2969
rect -1488 2911 -1477 2915
rect -1481 2823 -1477 2911
rect -2220 2659 -2194 2671
rect 607 2660 630 3332
rect 3984 3230 4009 3265
rect 3992 2922 4014 2977
rect 3277 2911 3292 2915
rect 3277 2823 3281 2911
rect -2221 2647 -2193 2659
rect -2220 2629 -2194 2647
rect -881 2636 -816 2656
rect -1488 2611 -1477 2615
rect -1481 2523 -1477 2611
rect -2221 2325 -2188 2370
rect -1488 2311 -1477 2315
rect -1481 2223 -1477 2311
rect -1498 2040 -1434 2059
rect -1481 1789 -1477 1877
rect -1492 1785 -1477 1789
rect -2220 1731 -2192 1767
rect -1453 1765 -1434 2040
rect -881 1765 -861 2636
rect 3996 2629 4015 2657
rect 3277 2611 3289 2615
rect 3277 2523 3281 2611
rect 3989 2324 4012 2369
rect 3277 2311 3289 2315
rect 3277 2223 3281 2311
rect 3990 2023 4020 2076
rect 3277 2011 3289 2015
rect 3277 1923 3281 2011
rect -1453 1746 -861 1765
rect -2225 1424 -2196 1481
rect 3987 1423 4016 1473
rect -1492 1411 -1477 1415
rect -1481 1323 -1477 1411
rect 3277 1411 3289 1415
rect 3277 1323 3281 1411
rect -2218 1124 -2191 1183
rect 3988 1131 4012 1169
rect -1488 1111 -1477 1115
rect -1481 1023 -1477 1111
rect 3277 1111 3289 1115
rect 3277 1023 3281 1111
rect -2224 825 -2194 878
rect 3986 831 4011 869
rect -1496 811 -1495 815
rect -1488 811 -1477 815
rect -1481 723 -1477 811
rect 3277 811 3289 815
rect 3277 723 3281 811
rect -2220 534 -2190 577
rect 3989 533 4006 567
rect -1490 511 -1477 515
rect -1481 423 -1477 511
rect 3277 511 3289 515
rect 3277 423 3281 511
rect 3986 228 4011 272
rect -1481 -11 -1477 77
rect -1492 -15 -1477 -11
rect -2225 -77 -2186 -27
rect 3994 -370 4019 -326
rect 3988 -668 4012 -631
rect 3989 -965 4011 -934
<< m2contact >>
rect -1477 3381 -1471 3387
rect -1177 3381 -1171 3387
rect -877 3381 -871 3387
rect -577 3381 -571 3387
rect -277 3381 -271 3387
rect 23 3375 29 3381
rect 623 3375 629 3381
rect 923 3375 929 3381
rect 1223 3375 1229 3381
rect 1523 3375 1529 3381
rect 1823 3381 1829 3387
rect 2123 3375 2129 3381
rect 2723 3381 2729 3387
rect 3023 3381 3029 3387
rect -1487 3123 -1481 3129
rect -1487 2823 -1481 2829
rect 3281 2823 3287 2829
rect -1487 2523 -1481 2529
rect -1487 2223 -1481 2229
rect -1487 1871 -1481 1877
rect 3281 2523 3287 2529
rect 3281 2223 3287 2229
rect 3281 1923 3287 1929
rect -1487 1323 -1481 1329
rect 3281 1323 3287 1329
rect -1487 1023 -1481 1029
rect 3281 1023 3287 1029
rect -1487 723 -1481 729
rect 3281 723 3287 729
rect -1487 423 -1481 429
rect 3281 423 3287 429
rect -1487 71 -1481 77
<< metal2 >>
rect -1450 3335 -1447 3381
rect -1150 3341 -1147 3381
rect -850 3347 -847 3381
rect -550 3353 -547 3381
rect -250 3359 -247 3381
rect 50 3365 53 3381
rect 644 3371 647 3381
rect 612 3368 647 3371
rect 50 3362 609 3365
rect -250 3356 603 3359
rect -550 3350 597 3353
rect -850 3344 591 3347
rect -1150 3338 585 3341
rect -1450 3332 579 3335
rect -1481 3150 -1434 3153
rect -1482 2850 -1440 2853
rect -1481 2550 -1446 2553
rect -1481 2250 -1452 2253
rect -1481 1853 -1458 1856
rect -1461 1746 -1458 1853
rect -1455 1752 -1452 2250
rect -1449 1758 -1446 2550
rect -1443 1764 -1440 2850
rect -1437 1770 -1434 3150
rect -908 2744 55 2747
rect -908 1770 -905 2744
rect -1437 1767 -905 1770
rect -902 2738 23 2741
rect -902 1764 -899 2738
rect -1443 1761 -899 1764
rect -896 2732 -81 2735
rect -896 1758 -893 2732
rect -1449 1755 -893 1758
rect -890 2726 -113 2729
rect -890 1752 -887 2726
rect -1455 1749 -887 1752
rect -884 2720 -161 2723
rect -884 1746 -881 2720
rect -1461 1743 -881 1746
rect -878 2714 -225 2717
rect -878 1740 -875 2714
rect -1461 1737 -875 1740
rect -872 2708 -241 2711
rect -1461 1353 -1458 1737
rect -872 1734 -869 2708
rect -1482 1350 -1458 1353
rect -1455 1731 -869 1734
rect -866 2702 -257 2705
rect -1455 1053 -1452 1731
rect -866 1728 -863 2702
rect -1481 1050 -1452 1053
rect -1449 1725 -863 1728
rect -860 2696 -281 2699
rect -1449 753 -1446 1725
rect -860 1722 -857 2696
rect -1481 750 -1446 753
rect -1443 1719 -857 1722
rect -854 2690 -299 2693
rect -284 2690 -281 2696
rect -1443 453 -1440 1719
rect -854 1716 -851 2690
rect -260 2689 -257 2702
rect -244 2689 -241 2708
rect -228 2690 -225 2714
rect -164 2690 -161 2720
rect -116 2690 -113 2726
rect -84 2690 -81 2732
rect 20 2690 23 2738
rect 52 2690 55 2744
rect 576 2723 579 3332
rect 92 2720 579 2723
rect 92 2690 95 2720
rect 582 2717 585 3338
rect 172 2714 585 2717
rect 172 2690 175 2714
rect 588 2711 591 3344
rect 188 2708 591 2711
rect 188 2692 191 2708
rect 594 2705 597 3350
rect 204 2702 597 2705
rect 204 2692 207 2702
rect 600 2699 603 3356
rect 244 2696 603 2699
rect 244 2690 247 2696
rect 606 2693 609 3362
rect 327 2690 609 2693
rect 612 2690 615 3368
rect 944 3365 947 3381
rect 618 3362 947 3365
rect 618 2693 621 3362
rect 1250 3359 1253 3381
rect 624 3356 1253 3359
rect 624 2699 627 3356
rect 1550 3353 1553 3381
rect 630 3350 1553 3353
rect 630 2705 633 3350
rect 1850 3347 1853 3381
rect 636 3344 1853 3347
rect 636 2711 639 3344
rect 2144 3341 2147 3381
rect 642 3338 2147 3341
rect 642 2717 645 3338
rect 2744 3335 2747 3381
rect 648 3332 2747 3335
rect 648 2723 651 3332
rect 3044 3329 3047 3381
rect 654 3326 3047 3329
rect 3234 3363 3281 3366
rect 654 2729 657 3326
rect 1422 2744 2688 2747
rect 654 2726 1111 2729
rect 648 2720 1079 2723
rect 642 2714 1015 2717
rect 636 2708 999 2711
rect 630 2702 791 2705
rect 624 2696 775 2699
rect 772 2693 775 2696
rect 618 2690 692 2693
rect 788 2690 791 2702
rect 996 2693 999 2708
rect 1012 2693 1015 2714
rect 1076 2690 1079 2720
rect 1108 2690 1111 2726
rect 1422 2693 1425 2744
rect 1140 2690 1425 2693
rect 1428 2738 2682 2741
rect 1428 2689 1431 2738
rect 1468 2732 2676 2735
rect 1468 2690 1471 2732
rect 1524 2726 2670 2729
rect 1524 2693 1527 2726
rect 1572 2720 2664 2723
rect 1572 2693 1575 2720
rect 1588 2714 2658 2717
rect 1588 2693 1591 2714
rect 1620 2708 2652 2711
rect 1620 2693 1623 2708
rect 1636 2702 2646 2705
rect 1636 2693 1639 2702
rect 1724 2696 2640 2699
rect 1724 2693 1727 2696
rect 2015 2690 2634 2693
rect 2012 2686 2015 2689
rect 2631 1746 2634 2690
rect 2637 1752 2640 2696
rect 2643 1758 2646 2702
rect 2649 1764 2652 2708
rect 2655 1770 2658 2714
rect 2661 1776 2664 2720
rect 2667 1782 2670 2726
rect 2673 1788 2676 2732
rect 2679 1794 2682 2738
rect 2685 1800 2688 2744
rect 3234 1800 3237 3363
rect 3271 3195 3292 3199
rect 3271 3129 3275 3195
rect 3271 3125 3283 3129
rect 3271 3123 3282 3125
rect 2685 1797 3237 1800
rect 3240 2850 3281 2853
rect 3240 1794 3243 2850
rect 2679 1791 3243 1794
rect 3246 2550 3281 2553
rect 3246 1788 3249 2550
rect 2673 1785 3249 1788
rect 3252 2250 3281 2253
rect 3252 1782 3255 2250
rect 2667 1779 3255 1782
rect 3258 1950 3281 1953
rect 3258 1776 3261 1950
rect 2661 1773 3261 1776
rect 2655 1767 3261 1770
rect 2649 1761 3255 1764
rect 2643 1755 3249 1758
rect 2637 1749 3243 1752
rect 2631 1743 3237 1746
rect -1481 450 -1440 453
rect -1437 1713 -851 1716
rect 2631 1737 3231 1740
rect -1437 56 -1434 1713
rect 2631 1295 2634 1737
rect 2637 1731 3225 1734
rect 2637 1301 2640 1731
rect 2643 1725 3219 1728
rect 2643 1307 2646 1725
rect 2643 1304 2655 1307
rect 2637 1298 2645 1301
rect 2642 1295 2645 1298
rect 2652 1295 2655 1304
rect -1481 53 -1434 56
rect -1490 -405 -1471 -401
rect -1477 -471 -1471 -405
rect -1483 -477 -1471 -471
rect -1490 -705 -1471 -701
rect -1477 -771 -1471 -705
rect -1483 -777 -1471 -771
rect 3216 -834 3219 1725
rect 3222 -534 3225 1731
rect 3228 -234 3231 1737
rect 3234 366 3237 1743
rect 3240 453 3243 1749
rect 3246 753 3249 1755
rect 3252 1053 3255 1761
rect 3258 1353 3261 1767
rect 3258 1350 3281 1353
rect 3252 1050 3281 1053
rect 3246 750 3281 753
rect 3240 450 3281 453
rect 3234 363 3281 366
rect 3274 195 3288 199
rect 3274 129 3278 195
rect 3274 127 3281 129
rect 3274 123 3289 127
rect 3228 -237 3281 -234
rect 3271 -405 3292 -401
rect 3271 -471 3275 -405
rect 3271 -474 3289 -471
rect 3271 -477 3284 -474
rect 3222 -537 3281 -534
rect 3271 -705 3292 -701
rect 3271 -771 3275 -705
rect 3271 -777 3285 -771
rect 3216 -837 3281 -834
rect -1520 -979 -1501 -975
rect -1507 -1001 -1501 -979
rect -1509 -1005 -1503 -1001
rect -1490 -1005 -1471 -1001
rect -1507 -1035 -1501 -1005
rect -1513 -1051 -1501 -1046
rect -1477 -1071 -1471 -1005
rect -1483 -1077 -1471 -1071
rect 3271 -1005 3292 -1001
rect 3271 -1071 3275 -1005
rect 3271 -1073 3286 -1071
rect 3271 -1077 3287 -1073
rect -1490 -1305 -1471 -1301
rect -1477 -1371 -1471 -1305
rect 3272 -1305 3292 -1301
rect 3272 -1371 3276 -1305
rect -1483 -1377 -1471 -1371
rect -1477 -1381 -1471 -1377
rect -1177 -1377 -1101 -1371
rect -1177 -1381 -1171 -1377
rect -1105 -1392 -1101 -1377
rect -877 -1377 -801 -1371
rect -877 -1381 -871 -1377
rect -805 -1388 -801 -1377
rect -577 -1377 -501 -1371
rect -577 -1381 -571 -1377
rect -505 -1388 -501 -1377
rect 23 -1377 99 -1371
rect 23 -1381 29 -1377
rect 95 -1388 99 -1377
rect 323 -1377 399 -1371
rect 323 -1381 329 -1377
rect 395 -1388 399 -1377
rect 623 -1377 699 -1371
rect 623 -1381 629 -1377
rect 695 -1388 699 -1377
rect 923 -1377 999 -1371
rect 923 -1381 929 -1377
rect 995 -1388 999 -1377
rect 1223 -1377 1299 -1371
rect 1223 -1381 1229 -1377
rect 1295 -1388 1299 -1377
rect 1823 -1377 1899 -1371
rect 1823 -1381 1829 -1377
rect 1895 -1388 1899 -1377
rect 2123 -1377 2199 -1371
rect 2123 -1381 2129 -1377
rect 2195 -1388 2199 -1377
rect 2423 -1377 2499 -1371
rect 2423 -1381 2429 -1377
rect 2495 -1388 2499 -1377
rect 2723 -1377 2799 -1371
rect 2723 -1381 2729 -1377
rect 2795 -1388 2799 -1377
rect 3023 -1377 3099 -1371
rect 3272 -1373 3288 -1371
rect 3272 -1377 3286 -1373
rect 3023 -1381 3029 -1377
rect 3095 -1388 3099 -1377
<< m3contact >>
rect 2631 1290 2636 1295
rect 2642 1290 2647 1295
rect 2652 1290 2657 1295
<< metal3 >>
rect 2630 1295 2637 1296
rect 2630 1290 2631 1295
rect 2636 1290 2637 1295
rect 2630 1289 2637 1290
rect 2641 1295 2648 1296
rect 2641 1290 2642 1295
rect 2647 1290 2648 1295
rect 2641 1289 2648 1290
rect 2651 1295 2658 1296
rect 2651 1290 2652 1295
rect 2657 1290 2658 1295
rect 2651 1289 2658 1290
rect 2631 1275 2636 1289
rect 2642 170 2647 1289
rect 2637 165 2647 170
rect 2652 150 2657 1289
rect 2636 145 2657 150
use PadFC  16_0
timestamp 1681001061
transform 1 0 -2500 0 1 3400
box 327 -3 1003 673
use PadFC  16_1
timestamp 1681001061
transform 0 1 3300 -1 0 4400
box 327 -3 1003 673
use PadFC  16_2
timestamp 1681001061
transform 0 -1 -1500 1 0 -2400
box 327 -3 1003 673
use PadFC  16_3
timestamp 1681001061
transform -1 0 4300 0 -1 -1400
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1711830429
transform 1 0 -1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1711830429
transform 1 0 -1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1711830429
transform 1 0 -900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1711830429
transform 1 0 -600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1711830429
transform 1 0 -300 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_5
timestamp 1711830429
transform 1 0 0 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1711830429
transform 1 0 600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1711830429
transform 1 0 900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1711830429
transform 1 0 1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1711830429
transform 0 -1 -1500 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1711830429
transform 0 -1 -1500 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1711830429
transform 0 -1 -1500 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1711830429
transform 0 -1 -1500 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_13
timestamp 1711830429
transform 0 -1 -1500 -1 0 1900
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1711830429
transform 0 -1 -1500 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1711830429
transform 0 -1 -1500 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1711830429
transform 0 -1 -1500 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1711830429
transform 0 1 3300 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1711830429
transform 0 1 3300 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_19
timestamp 1711830429
transform 0 1 3300 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1711830429
transform 0 1 3300 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1711830429
transform 0 1 3300 1 0 1900
box -36 -19 303 1000
use PadBiDir  17_22
timestamp 1711830429
transform 0 1 3300 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1711830429
transform 0 1 3300 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1711830429
transform 0 1 3300 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1711830429
transform 0 -1 -1500 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_26
timestamp 1711830429
transform 1 0 -1500 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1711830429
transform 1 0 -1200 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1711830429
transform 1 0 -900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1711830429
transform 1 0 -600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_30
timestamp 1711830429
transform 1 0 0 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1711830429
transform 1 0 300 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1711830429
transform 1 0 600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1711830429
transform 1 0 900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1711830429
transform 0 1 3300 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1711830429
transform 1 0 1200 0 -1 -1400
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1711831643
transform 1 0 300 0 1 3400
box -3 -16 303 1000
use PadVdd  18_1
timestamp 1711831643
transform 1 0 -300 0 -1 -1400
box -3 -16 303 1000
use PadGnd  19_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 2200
box -3 -11 303 1000
use PadGnd  19_1
timestamp 1711831454
transform 0 1 3300 -1 0 1900
box -3 -11 303 1000
use PadBiDir  PadBiDir_0
timestamp 1711830429
transform 1 0 1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_1
timestamp 1711830429
transform 1 0 1800 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_2
timestamp 1711830429
transform 1 0 2100 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_3
timestamp 1711830429
transform 1 0 2700 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_4
timestamp 1711830429
transform 1 0 3000 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_5
timestamp 1711830429
transform 1 0 1800 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_6
timestamp 1711830429
transform 1 0 2100 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_7
timestamp 1711830429
transform 1 0 2400 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_8
timestamp 1711830429
transform 1 0 2700 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_9
timestamp 1711830429
transform 1 0 3000 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_10
timestamp 1711830429
transform 0 -1 -1500 -1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_11
timestamp 1711830429
transform 0 -1 -1500 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_12
timestamp 1711830429
transform 0 -1 -1500 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_13
timestamp 1711830429
transform 0 -1 -1500 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_14
timestamp 1711830429
transform 0 -1 -1500 1 0 1300
box -36 -19 303 1000
use PadBiDir  PadBiDir_15
timestamp 1711830429
transform 0 1 3300 1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_16
timestamp 1711830429
transform 0 1 3300 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_17
timestamp 1711830429
transform 0 1 3300 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_18
timestamp 1711830429
transform 0 1 3300 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_19
timestamp 1711830429
transform 0 1 3300 1 0 1300
box -36 -19 303 1000
use PadGnd  PadGnd_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 400
box -3 -11 303 1000
use PadGnd  PadGnd_1
timestamp 1711831454
transform 0 1 3300 -1 0 100
box -3 -11 303 1000
use PadVdd  PadVdd_0
timestamp 1711831643
transform 1 0 2400 0 1 3400
box -3 -16 303 1000
use PadVdd  PadVdd_1
timestamp 1711831643
transform 1 0 1500 0 -1 -1400
box -3 -16 303 1000
use top_module  top_module_0 ./foo
timestamp 1712693004
transform 1 0 -862 0 1 -647
box 14 13 3504 3340
<< labels >>
rlabel metal1 -2206 -51 -2206 -51 1 p_board_out[26]
rlabel metal1 -2205 555 -2205 555 1 p_board_out[25]
rlabel metal1 -2206 854 -2206 854 1 p_board_out[27]
rlabel metal1 -2205 1154 -2205 1154 1 p_board_out[24]
rlabel metal1 -2210 1453 -2210 1453 1 p_board_out[28]
rlabel metal1 -2207 1749 -2207 1749 1 p_board_out[29]
rlabel metal1 -2204 2350 -2204 2350 1 p_board_out[22]
rlabel metal1 -2207 2653 -2207 2653 1 p_board_out[23]
rlabel metal1 -2208 2956 -2208 2956 1 p_board_out[30]
rlabel metal1 -2208 3253 -2208 3253 1 p_board_out[21]
rlabel metal1 -1350 4109 -1350 4109 1 p_board_out[31]
rlabel metal1 -1049 4108 -1049 4108 1 p_board_out[20]
rlabel metal1 -744 4112 -744 4112 1 p_board_out[19]
rlabel metal1 -446 4107 -444 4107 1 p_board_out[18]
rlabel metal1 -145 4105 -145 4105 1 p_board_out[17]
rlabel metal1 152 4105 152 4105 1 p_board_out[16]
rlabel metal1 750 4106 750 4106 1 p_board_out[15]
rlabel metal1 1052 4107 1052 4107 1 p_board_out[14]
rlabel metal1 1353 4105 1353 4105 1 p_board_out[13]
rlabel metal1 1651 4108 1651 4108 1 p_board_out[12]
rlabel metal1 1950 4105 1950 4105 1 p_board_out[11]
rlabel metal1 2253 4103 2253 4103 1 p_board_out[8]
rlabel metal1 2852 4104 2852 4104 1 p_board_out[10]
rlabel metal1 3156 4108 3156 4108 1 p_board_out[9]
rlabel metal1 3996 3249 3996 3249 1 p_in_clkb
rlabel metal1 4002 2954 4002 2954 1 p_board_out[7]
rlabel metal1 4005 2645 4005 2645 1 p_board_out[3]
rlabel metal1 4001 2349 4001 2349 1 p_board_out[0]
rlabel metal1 4003 2051 4003 2051 1 p_board_out[6]
rlabel metal1 3998 1456 3998 1456 1 p_board_out[4]
rlabel metal1 3998 1146 3998 1146 1 p_board_out[1]
rlabel metal1 3995 849 3995 849 1 p_board_out[5]
rlabel metal1 3999 552 3999 552 1 p_board_out[2]
rlabel metal1 3998 251 3998 251 1 p_in_clka
rlabel metal1 4005 -347 4005 -347 1 p_in_restart
rlabel metal1 4000 -651 4000 -651 1 p_in_move[0]
rlabel metal1 4000 -948 4000 -948 1 p_in_move[1]
<< end >>
